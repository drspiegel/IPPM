
module s1196(GND, VDD, CK, G0, G1, G10, G11, G12, G13, G2, G3, G4, G45, G5, G530, G532, G535, G537, G539, G542, G546, G547, G548, G549, G550, G551, G552, G6, G7, G8, G9);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  input CK;
  wire \DFF_0.CK ;
  wire \DFF_0.D ;
  wire \DFF_0.Q ;
  wire \DFF_1.CK ;
  wire \DFF_1.D ;
  wire \DFF_1.Q ;
  wire \DFF_10.CK ;
  wire \DFF_10.D ;
  wire \DFF_10.Q ;
  wire \DFF_11.CK ;
  wire \DFF_11.D ;
  wire \DFF_11.Q ;
  wire \DFF_12.CK ;
  wire \DFF_12.D ;
  wire \DFF_12.Q ;
  wire \DFF_13.CK ;
  wire \DFF_13.D ;
  wire \DFF_13.Q ;
  wire \DFF_14.CK ;
  wire \DFF_14.D ;
  wire \DFF_14.Q ;
  wire \DFF_15.CK ;
  wire \DFF_15.D ;
  wire \DFF_15.Q ;
  wire \DFF_16.CK ;
  wire \DFF_16.D ;
  wire \DFF_16.Q ;
  wire \DFF_17.CK ;
  wire \DFF_17.D ;
  wire \DFF_17.Q ;
  wire \DFF_2.CK ;
  wire \DFF_2.D ;
  wire \DFF_2.Q ;
  wire \DFF_3.CK ;
  wire \DFF_3.D ;
  wire \DFF_3.Q ;
  wire \DFF_4.CK ;
  wire \DFF_4.D ;
  wire \DFF_4.Q ;
  wire \DFF_5.CK ;
  wire \DFF_5.D ;
  wire \DFF_5.Q ;
  wire \DFF_6.CK ;
  wire \DFF_6.D ;
  wire \DFF_6.Q ;
  wire \DFF_7.CK ;
  wire \DFF_7.D ;
  wire \DFF_7.Q ;
  wire \DFF_8.CK ;
  wire \DFF_8.D ;
  wire \DFF_8.Q ;
  wire \DFF_9.CK ;
  wire \DFF_9.D ;
  wire \DFF_9.Q ;
  input G0;
  input G1;
  input G10;
  wire G107;
  input G11;
  input G12;
  input G13;
  wire G153;
  wire G165;
  input G2;
  wire G228;
  wire G29;
  input G3;
  wire G30;
  wire G31;
  wire G32;
  wire G33;
  wire G334;
  wire G335;
  wire G34;
  wire G35;
  wire G36;
  wire G37;
  wire G38;
  wire G39;
  input G4;
  wire G40;
  wire G41;
  wire G42;
  wire G43;
  wire G44;
  output G45;
  wire G46;
  input G5;
  wire G502;
  wire G503;
  wire G504;
  wire G505;
  wire G506;
  wire G507;
  wire G508;
  wire G509;
  wire G510;
  wire G511;
  wire G512;
  wire G513;
  wire G514;
  wire G515;
  wire G516;
  wire G517;
  wire G518;
  wire G519;
  output G530;
  output G532;
  output G535;
  output G537;
  output G539;
  output G542;
  output G546;
  output G547;
  output G548;
  output G549;
  output G550;
  output G551;
  output G552;
  input G6;
  input G7;
  input G8;
  input G9;
  input GND;
  wire II218;
  wire II249;
  wire II374;
  input VDD;
  al_and2ft _268_ (
    .a(G6),
    .b(G9),
    .y(_237_)
  );
  al_and2ft _269_ (
    .a(G9),
    .b(G6),
    .y(_238_)
  );
  al_or2 _270_ (
    .a(_237_),
    .b(_238_),
    .y(\DFF_8.D )
  );
  al_oai21ftf _271_ (
    .a(G11),
    .b(G9),
    .c(G10),
    .y(\DFF_1.D )
  );
  al_nand3ftt _272_ (
    .a(G2),
    .b(G3),
    .c(G5),
    .y(_239_)
  );
  al_nand2ft _273_ (
    .a(G3),
    .b(G2),
    .y(_240_)
  );
  al_and2ft _274_ (
    .a(G5),
    .b(G2),
    .y(_241_)
  );
  al_nand3ftt _275_ (
    .a(_241_),
    .b(_239_),
    .c(_240_),
    .y(\DFF_10.D )
  );
  al_ao21ttf _276_ (
    .a(G11),
    .b(G9),
    .c(G10),
    .y(_242_)
  );
  al_ao21ftf _277_ (
    .a(G7),
    .b(G11),
    .c(_242_),
    .y(\DFF_2.D )
  );
  al_oai21ftf _278_ (
    .a(G6),
    .b(G4),
    .c(G5),
    .y(_243_)
  );
  al_nand3ftt _279_ (
    .a(G2),
    .b(G3),
    .c(_243_),
    .y(_244_)
  );
  al_and3 _280_ (
    .a(G3),
    .b(G4),
    .c(G6),
    .y(_245_)
  );
  al_or3fft _281_ (
    .a(G2),
    .b(G5),
    .c(_245_),
    .y(_246_)
  );
  al_nand3ftt _282_ (
    .a(G5),
    .b(G2),
    .c(G4),
    .y(_247_)
  );
  al_nand3 _283_ (
    .a(_247_),
    .b(_244_),
    .c(_246_),
    .y(\DFF_3.D )
  );
  al_inv _284_ (
    .a(G9),
    .y(_248_)
  );
  al_and2ft _285_ (
    .a(G10),
    .b(G7),
    .y(_249_)
  );
  al_nand3ftt _286_ (
    .a(G9),
    .b(G8),
    .c(_249_),
    .y(_250_)
  );
  al_and3fft _287_ (
    .a(G7),
    .b(G8),
    .c(G10),
    .y(_251_)
  );
  al_ao21ftf _288_ (
    .a(_248_),
    .b(_251_),
    .c(_250_),
    .y(_252_)
  );
  al_and3fft _289_ (
    .a(G8),
    .b(G9),
    .c(G7),
    .y(_253_)
  );
  al_and2ft _290_ (
    .a(G10),
    .b(_253_),
    .y(_254_)
  );
  al_mux2h _291_ (
    .a(_254_),
    .b(_252_),
    .s(G6),
    .y(\DFF_6.D )
  );
  al_nand2 _292_ (
    .a(G2),
    .b(G1),
    .y(_255_)
  );
  al_and3 _293_ (
    .a(G8),
    .b(G11),
    .c(G9),
    .y(_256_)
  );
  al_nand3 _294_ (
    .a(G7),
    .b(G10),
    .c(_256_),
    .y(_257_)
  );
  al_nand2 _295_ (
    .a(G3),
    .b(G0),
    .y(_258_)
  );
  al_and3 _296_ (
    .a(G4),
    .b(G6),
    .c(G5),
    .y(_259_)
  );
  al_or3ftt _297_ (
    .a(_259_),
    .b(_258_),
    .c(_257_),
    .y(_260_)
  );
  al_or2 _298_ (
    .a(G3),
    .b(G5),
    .y(_261_)
  );
  al_nand3ftt _299_ (
    .a(_261_),
    .b(_238_),
    .c(_251_),
    .y(_262_)
  );
  al_nand3 _300_ (
    .a(G3),
    .b(G8),
    .c(G5),
    .y(_263_)
  );
  al_or3fft _301_ (
    .a(\DFF_8.Q ),
    .b(_249_),
    .c(_263_),
    .y(_264_)
  );
  al_or3ftt _302_ (
    .a(G11),
    .b(G4),
    .c(G0),
    .y(_265_)
  );
  al_ao21 _303_ (
    .a(_264_),
    .b(_262_),
    .c(_265_),
    .y(_266_)
  );
  al_aoi21 _304_ (
    .a(_260_),
    .b(_266_),
    .c(_255_),
    .y(_267_)
  );
  al_nand2ft _305_ (
    .a(G5),
    .b(G4),
    .y(_000_)
  );
  al_ao21ttf _306_ (
    .a(G3),
    .b(G5),
    .c(G4),
    .y(_001_)
  );
  al_ao21ftf _307_ (
    .a(G1),
    .b(G5),
    .c(_001_),
    .y(_002_)
  );
  al_ao21 _308_ (
    .a(G2),
    .b(_002_),
    .c(_261_),
    .y(_003_)
  );
  al_and2ft _309_ (
    .a(G4),
    .b(G3),
    .y(_004_)
  );
  al_nand2ft _310_ (
    .a(G0),
    .b(_004_),
    .y(_005_)
  );
  al_ao21ttf _311_ (
    .a(_005_),
    .b(_003_),
    .c(_000_),
    .y(_006_)
  );
  al_inv _312_ (
    .a(G11),
    .y(_007_)
  );
  al_or3 _313_ (
    .a(G7),
    .b(G8),
    .c(G9),
    .y(_008_)
  );
  al_oa21 _314_ (
    .a(G6),
    .b(\DFF_1.Q ),
    .c(_008_),
    .y(_009_)
  );
  al_nand2 _315_ (
    .a(G8),
    .b(G10),
    .y(_010_)
  );
  al_nand3ftt _316_ (
    .a(G6),
    .b(G7),
    .c(\DFF_1.Q ),
    .y(_011_)
  );
  al_and3ftt _317_ (
    .a(\DFF_2.Q ),
    .b(G8),
    .c(_011_),
    .y(_012_)
  );
  al_ao21ftf _318_ (
    .a(_248_),
    .b(_010_),
    .c(_012_),
    .y(_013_)
  );
  al_aoi21 _319_ (
    .a(_009_),
    .b(_013_),
    .c(_007_),
    .y(_014_)
  );
  al_nand2 _320_ (
    .a(G8),
    .b(\DFF_2.Q ),
    .y(_015_)
  );
  al_oa21ttf _321_ (
    .a(G8),
    .b(G10),
    .c(G11),
    .y(_016_)
  );
  al_and3ftt _322_ (
    .a(G7),
    .b(G9),
    .c(_015_),
    .y(_017_)
  );
  al_aoi21ttf _323_ (
    .a(_016_),
    .b(_017_),
    .c(\DFF_17.Q ),
    .y(_018_)
  );
  al_nor2 _324_ (
    .a(G11),
    .b(G10),
    .y(_019_)
  );
  al_nand3ftt _325_ (
    .a(G9),
    .b(_011_),
    .c(_019_),
    .y(_020_)
  );
  al_aoi21ftf _326_ (
    .a(_020_),
    .b(_015_),
    .c(_018_),
    .y(_021_)
  );
  al_and3ftt _327_ (
    .a(_014_),
    .b(_006_),
    .c(_021_),
    .y(_022_)
  );
  al_nand2ft _328_ (
    .a(G13),
    .b(G12),
    .y(_023_)
  );
  al_and3fft _329_ (
    .a(_023_),
    .b(_022_),
    .c(_267_),
    .y(_024_)
  );
  al_inv _330_ (
    .a(G2),
    .y(_025_)
  );
  al_nand2ft _331_ (
    .a(G5),
    .b(G11),
    .y(_026_)
  );
  al_nor3fft _332_ (
    .a(\DFF_6.Q ),
    .b(_004_),
    .c(_026_),
    .y(_027_)
  );
  al_inv _333_ (
    .a(G5),
    .y(_028_)
  );
  al_inv _334_ (
    .a(_245_),
    .y(_029_)
  );
  al_nand3fft _335_ (
    .a(G7),
    .b(G8),
    .c(_019_),
    .y(_030_)
  );
  al_oai21ftt _336_ (
    .a(G9),
    .b(_030_),
    .c(_257_),
    .y(_031_)
  );
  al_nand3fft _337_ (
    .a(_028_),
    .b(_029_),
    .c(_031_),
    .y(_032_)
  );
  al_nand3fft _338_ (
    .a(_025_),
    .b(_027_),
    .c(_032_),
    .y(_033_)
  );
  al_nand2ft _339_ (
    .a(G6),
    .b(\DFF_7.Q ),
    .y(_034_)
  );
  al_nand3 _340_ (
    .a(G11),
    .b(_259_),
    .c(_252_),
    .y(_035_)
  );
  al_ao21 _341_ (
    .a(_034_),
    .b(_035_),
    .c(G3),
    .y(_036_)
  );
  al_and2ft _342_ (
    .a(G7),
    .b(G8),
    .y(_037_)
  );
  al_nand3ftt _343_ (
    .a(G10),
    .b(G9),
    .c(_037_),
    .y(_038_)
  );
  al_nand3ftt _344_ (
    .a(G5),
    .b(G11),
    .c(_245_),
    .y(_039_)
  );
  al_oai21ftf _345_ (
    .a(_038_),
    .b(_252_),
    .c(_039_),
    .y(_040_)
  );
  al_nand3 _346_ (
    .a(_025_),
    .b(_040_),
    .c(_036_),
    .y(_041_)
  );
  al_inv _347_ (
    .a(G12),
    .y(_042_)
  );
  al_and2 _348_ (
    .a(G7),
    .b(G10),
    .y(_043_)
  );
  al_and3ftt _349_ (
    .a(G10),
    .b(G7),
    .c(G9),
    .y(_044_)
  );
  al_aoi21 _350_ (
    .a(\DFF_1.Q ),
    .b(_037_),
    .c(_044_),
    .y(_045_)
  );
  al_ao21ftf _351_ (
    .a(_256_),
    .b(_043_),
    .c(_045_),
    .y(_046_)
  );
  al_aoi21 _352_ (
    .a(\DFF_3.Q ),
    .b(_046_),
    .c(G13),
    .y(_047_)
  );
  al_and2 _353_ (
    .a(_042_),
    .b(_047_),
    .y(_048_)
  );
  al_nand3 _354_ (
    .a(_033_),
    .b(_048_),
    .c(_041_),
    .y(_049_)
  );
  al_and2ft _355_ (
    .a(G1),
    .b(G3),
    .y(_050_)
  );
  al_nand3 _356_ (
    .a(G4),
    .b(G6),
    .c(_050_),
    .y(_051_)
  );
  al_and3ftt _357_ (
    .a(G4),
    .b(G3),
    .c(G1),
    .y(_052_)
  );
  al_nand2 _358_ (
    .a(G6),
    .b(_052_),
    .y(_053_)
  );
  al_nand3 _359_ (
    .a(G8),
    .b(_053_),
    .c(_051_),
    .y(_054_)
  );
  al_nor2 _360_ (
    .a(G4),
    .b(G6),
    .y(_055_)
  );
  al_ao21 _361_ (
    .a(_050_),
    .b(_055_),
    .c(G8),
    .y(_056_)
  );
  al_and3ftt _362_ (
    .a(G9),
    .b(G11),
    .c(_249_),
    .y(_057_)
  );
  al_nand3 _363_ (
    .a(_056_),
    .b(_057_),
    .c(_054_),
    .y(_058_)
  );
  al_and3ftt _364_ (
    .a(G8),
    .b(G11),
    .c(G9),
    .y(_059_)
  );
  al_and2 _365_ (
    .a(G10),
    .b(_059_),
    .y(_060_)
  );
  al_and2ft _366_ (
    .a(G10),
    .b(_256_),
    .y(_061_)
  );
  al_ao21ftt _367_ (
    .a(_051_),
    .b(_061_),
    .c(_060_),
    .y(_062_)
  );
  al_ao21 _368_ (
    .a(_053_),
    .b(_051_),
    .c(G7),
    .y(_063_)
  );
  al_ao21ftf _369_ (
    .a(_063_),
    .b(_062_),
    .c(_058_),
    .y(_064_)
  );
  al_or3fft _370_ (
    .a(G2),
    .b(G1),
    .c(_032_),
    .y(_065_)
  );
  al_ao21ttf _371_ (
    .a(_241_),
    .b(_064_),
    .c(_065_),
    .y(_066_)
  );
  al_nand3ftt _372_ (
    .a(G1),
    .b(G2),
    .c(_243_),
    .y(_067_)
  );
  al_inv _373_ (
    .a(G6),
    .y(_068_)
  );
  al_ao21ttf _374_ (
    .a(G2),
    .b(G5),
    .c(G4),
    .y(_069_)
  );
  al_aoi21 _375_ (
    .a(_240_),
    .b(_069_),
    .c(_068_),
    .y(_070_)
  );
  al_nand2 _376_ (
    .a(G2),
    .b(G4),
    .y(_071_)
  );
  al_nand2ft _377_ (
    .a(G4),
    .b(G5),
    .y(_072_)
  );
  al_aoi21 _378_ (
    .a(_072_),
    .b(_071_),
    .c(G6),
    .y(_073_)
  );
  al_or3ftt _379_ (
    .a(G4),
    .b(G3),
    .c(G5),
    .y(_074_)
  );
  al_nand3ftt _380_ (
    .a(G2),
    .b(G3),
    .c(G6),
    .y(_075_)
  );
  al_and2 _381_ (
    .a(G3),
    .b(G5),
    .y(_076_)
  );
  al_ao21ttf _382_ (
    .a(G4),
    .b(G6),
    .c(_076_),
    .y(_077_)
  );
  al_and3 _383_ (
    .a(_074_),
    .b(_075_),
    .c(_077_),
    .y(_078_)
  );
  al_nand3fft _384_ (
    .a(_070_),
    .b(_073_),
    .c(_078_),
    .y(_079_)
  );
  al_ao21ttf _385_ (
    .a(G1),
    .b(_079_),
    .c(_067_),
    .y(_080_)
  );
  al_nand2ft _386_ (
    .a(G12),
    .b(G13),
    .y(_081_)
  );
  al_aoi21 _387_ (
    .a(_046_),
    .b(_080_),
    .c(_081_),
    .y(_082_)
  );
  al_ao21ttf _388_ (
    .a(_066_),
    .b(_082_),
    .c(_049_),
    .y(_083_)
  );
  al_or2 _389_ (
    .a(_024_),
    .b(_083_),
    .y(\DFF_16.D )
  );
  al_ao21ttf _390_ (
    .a(G8),
    .b(G9),
    .c(\DFF_5.Q ),
    .y(_084_)
  );
  al_nand3ftt _391_ (
    .a(_023_),
    .b(G6),
    .c(_022_),
    .y(_085_)
  );
  al_nand2 _392_ (
    .a(G8),
    .b(\DFF_5.Q ),
    .y(_086_)
  );
  al_ao21ttf _393_ (
    .a(_086_),
    .b(_085_),
    .c(_044_),
    .y(_087_)
  );
  al_oai21ftf _394_ (
    .a(G7),
    .b(G8),
    .c(G10),
    .y(_088_)
  );
  al_oa21ftt _395_ (
    .a(G8),
    .b(G7),
    .c(G9),
    .y(_089_)
  );
  al_ao21ftt _396_ (
    .a(_089_),
    .b(_088_),
    .c(_060_),
    .y(_090_)
  );
  al_aoi21ftf _397_ (
    .a(_085_),
    .b(_090_),
    .c(_087_),
    .y(_091_)
  );
  al_ao21ftf _398_ (
    .a(_084_),
    .b(_043_),
    .c(_091_),
    .y(G542)
  );
  al_nand2ft _399_ (
    .a(G2),
    .b(G3),
    .y(_092_)
  );
  al_mux2l _400_ (
    .a(G3),
    .b(G5),
    .s(G4),
    .y(_093_)
  );
  al_nand3ftt _401_ (
    .a(G1),
    .b(G2),
    .c(_093_),
    .y(_094_)
  );
  al_aoi21ftf _402_ (
    .a(_092_),
    .b(_000_),
    .c(_094_),
    .y(\DFF_0.D )
  );
  al_nand3 _403_ (
    .a(G6),
    .b(_000_),
    .c(_072_),
    .y(_095_)
  );
  al_inv _404_ (
    .a(G1),
    .y(_096_)
  );
  al_nor2 _405_ (
    .a(G6),
    .b(G5),
    .y(_097_)
  );
  al_aoi21 _406_ (
    .a(_097_),
    .b(_071_),
    .c(_096_),
    .y(_098_)
  );
  al_ao21ttf _407_ (
    .a(_095_),
    .b(_098_),
    .c(_067_),
    .y(_099_)
  );
  al_nor3fft _408_ (
    .a(G6),
    .b(G1),
    .c(_092_),
    .y(_100_)
  );
  al_aoi21 _409_ (
    .a(G3),
    .b(_099_),
    .c(_100_),
    .y(\DFF_14.D )
  );
  al_and2 _410_ (
    .a(G6),
    .b(G9),
    .y(_101_)
  );
  al_nand3 _411_ (
    .a(G8),
    .b(G10),
    .c(_238_),
    .y(_102_)
  );
  al_aoi21ftf _412_ (
    .a(_043_),
    .b(_101_),
    .c(_102_),
    .y(_103_)
  );
  al_nand2ft _413_ (
    .a(G10),
    .b(G9),
    .y(_104_)
  );
  al_and2ft _414_ (
    .a(G6),
    .b(G7),
    .y(_105_)
  );
  al_aoi21 _415_ (
    .a(_104_),
    .b(_105_),
    .c(_253_),
    .y(_106_)
  );
  al_ao21 _416_ (
    .a(_106_),
    .b(_103_),
    .c(_007_),
    .y(\DFF_13.D )
  );
  al_aoi21 _417_ (
    .a(_030_),
    .b(_257_),
    .c(G5),
    .y(\DFF_7.D )
  );
  al_ao21ftf _418_ (
    .a(G10),
    .b(_256_),
    .c(_015_),
    .y(_107_)
  );
  al_and2 _419_ (
    .a(G7),
    .b(G9),
    .y(_108_)
  );
  al_nand3ftt _420_ (
    .a(G11),
    .b(G6),
    .c(_108_),
    .y(_109_)
  );
  al_ao21ttf _421_ (
    .a(_011_),
    .b(_109_),
    .c(G8),
    .y(_110_)
  );
  al_aoi21ftf _422_ (
    .a(_068_),
    .b(_107_),
    .c(_110_),
    .y(\DFF_11.D )
  );
  al_or3 _423_ (
    .a(G4),
    .b(G6),
    .c(G5),
    .y(_111_)
  );
  al_nand3ftt _424_ (
    .a(_111_),
    .b(_256_),
    .c(_043_),
    .y(_112_)
  );
  al_and2 _425_ (
    .a(G9),
    .b(_251_),
    .y(_113_)
  );
  al_nand3 _426_ (
    .a(G11),
    .b(_259_),
    .c(_113_),
    .y(_114_)
  );
  al_nand3ftt _427_ (
    .a(_008_),
    .b(_019_),
    .c(_097_),
    .y(_115_)
  );
  al_and3 _428_ (
    .a(_115_),
    .b(_112_),
    .c(_114_),
    .y(\DFF_15.D )
  );
  al_oai21ftf _429_ (
    .a(G4),
    .b(G5),
    .c(G3),
    .y(_116_)
  );
  al_ao21 _430_ (
    .a(G2),
    .b(_002_),
    .c(_116_),
    .y(_117_)
  );
  al_oa21 _431_ (
    .a(_092_),
    .b(_000_),
    .c(G0),
    .y(_118_)
  );
  al_ao21 _432_ (
    .a(_118_),
    .b(_117_),
    .c(G1),
    .y(_119_)
  );
  al_aoi21 _433_ (
    .a(G7),
    .b(G10),
    .c(G6),
    .y(_120_)
  );
  al_ao21ttf _434_ (
    .a(G7),
    .b(\DFF_1.Q ),
    .c(_120_),
    .y(_121_)
  );
  al_oai21ftt _435_ (
    .a(G3),
    .b(G4),
    .c(G0),
    .y(_122_)
  );
  al_ao21ftf _436_ (
    .a(G1),
    .b(G3),
    .c(_122_),
    .y(_123_)
  );
  al_or3fft _437_ (
    .a(G2),
    .b(_123_),
    .c(_002_),
    .y(_124_)
  );
  al_and3 _438_ (
    .a(_121_),
    .b(_124_),
    .c(_119_),
    .y(\DFF_17.D )
  );
  al_and3 _439_ (
    .a(_042_),
    .b(\DFF_3.Q ),
    .c(_046_),
    .y(_125_)
  );
  al_aoi21ftt _440_ (
    .a(_081_),
    .b(_046_),
    .c(_125_),
    .y(_126_)
  );
  al_oa21ftf _441_ (
    .a(G13),
    .b(_080_),
    .c(_126_),
    .y(\DFF_5.D )
  );
  al_and3ftt _442_ (
    .a(G4),
    .b(G1),
    .c(G0),
    .y(_127_)
  );
  al_nand3 _443_ (
    .a(G12),
    .b(_127_),
    .c(_022_),
    .y(_128_)
  );
  al_aoi21ftf _444_ (
    .a(_247_),
    .b(_125_),
    .c(_128_),
    .y(\DFF_4.D )
  );
  al_and2ft _445_ (
    .a(_023_),
    .b(_022_),
    .y(_129_)
  );
  al_nand3ftt _446_ (
    .a(_101_),
    .b(_043_),
    .c(_129_),
    .y(_130_)
  );
  al_inv _447_ (
    .a(\DFF_5.Q ),
    .y(_131_)
  );
  al_or3 _448_ (
    .a(_131_),
    .b(_010_),
    .c(_108_),
    .y(_132_)
  );
  al_and3 _449_ (
    .a(_132_),
    .b(_130_),
    .c(_087_),
    .y(\DFF_12.D )
  );
  al_inv _450_ (
    .a(\DFF_12.Q ),
    .y(G546)
  );
  al_ao21ttf _451_ (
    .a(_033_),
    .b(_041_),
    .c(_048_),
    .y(_133_)
  );
  al_or3 _452_ (
    .a(_267_),
    .b(_023_),
    .c(_022_),
    .y(_134_)
  );
  al_nand2 _453_ (
    .a(_046_),
    .b(_080_),
    .y(_135_)
  );
  al_inv _454_ (
    .a(_081_),
    .y(_136_)
  );
  al_or3fft _455_ (
    .a(_136_),
    .b(_135_),
    .c(_066_),
    .y(_137_)
  );
  al_nand3 _456_ (
    .a(_134_),
    .b(_133_),
    .c(_137_),
    .y(G539)
  );
  al_and3ftt _457_ (
    .a(\DFF_0.Q ),
    .b(G0),
    .c(_129_),
    .y(_138_)
  );
  al_and3ftt _458_ (
    .a(G0),
    .b(G4),
    .c(G1),
    .y(_139_)
  );
  al_and3 _459_ (
    .a(G3),
    .b(_139_),
    .c(_129_),
    .y(_140_)
  );
  al_and3 _460_ (
    .a(_046_),
    .b(_136_),
    .c(_080_),
    .y(_141_)
  );
  al_and3 _461_ (
    .a(G4),
    .b(G5),
    .c(G1),
    .y(_142_)
  );
  al_ao21 _462_ (
    .a(G4),
    .b(G1),
    .c(G5),
    .y(_143_)
  );
  al_nor3fft _463_ (
    .a(G2),
    .b(_143_),
    .c(_142_),
    .y(_144_)
  );
  al_nand2 _464_ (
    .a(_144_),
    .b(_141_),
    .y(_145_)
  );
  al_inv _465_ (
    .a(G13),
    .y(_146_)
  );
  al_nand3ftt _466_ (
    .a(\DFF_4.Q ),
    .b(G3),
    .c(_146_),
    .y(_147_)
  );
  al_and2 _467_ (
    .a(_146_),
    .b(_125_),
    .y(_148_)
  );
  al_nand3 _468_ (
    .a(_076_),
    .b(_071_),
    .c(_148_),
    .y(_149_)
  );
  al_and3 _469_ (
    .a(_147_),
    .b(_149_),
    .c(_145_),
    .y(_150_)
  );
  al_nand3fft _470_ (
    .a(_140_),
    .b(_138_),
    .c(_150_),
    .y(G550)
  );
  al_inv _471_ (
    .a(G3),
    .y(_151_)
  );
  al_and2 _472_ (
    .a(G2),
    .b(G0),
    .y(_152_)
  );
  al_mux2l _473_ (
    .a(G4),
    .b(G1),
    .s(_152_),
    .y(_153_)
  );
  al_and2 _474_ (
    .a(G4),
    .b(G1),
    .y(_154_)
  );
  al_mux2l _475_ (
    .a(G0),
    .b(_258_),
    .s(_154_),
    .y(_155_)
  );
  al_ao21ttf _476_ (
    .a(_151_),
    .b(_153_),
    .c(_155_),
    .y(_156_)
  );
  al_nand3 _477_ (
    .a(G5),
    .b(_156_),
    .c(_129_),
    .y(_157_)
  );
  al_nand3 _478_ (
    .a(G4),
    .b(\DFF_10.Q ),
    .c(_148_),
    .y(_158_)
  );
  al_nand3ftt _479_ (
    .a(G3),
    .b(G4),
    .c(G6),
    .y(_159_)
  );
  al_ao21ftf _480_ (
    .a(G4),
    .b(_075_),
    .c(_028_),
    .y(_160_)
  );
  al_ao21 _481_ (
    .a(_159_),
    .b(_160_),
    .c(_096_),
    .y(_161_)
  );
  al_and3ftt _482_ (
    .a(G1),
    .b(G2),
    .c(G4),
    .y(_162_)
  );
  al_aoi21ftt _483_ (
    .a(_092_),
    .b(_154_),
    .c(_162_),
    .y(_163_)
  );
  al_nand2 _484_ (
    .a(_163_),
    .b(_161_),
    .y(_164_)
  );
  al_or3fft _485_ (
    .a(_136_),
    .b(_164_),
    .c(_135_),
    .y(_165_)
  );
  al_nand3 _486_ (
    .a(_158_),
    .b(_165_),
    .c(_157_),
    .y(G551)
  );
  al_ao21ttf _487_ (
    .a(G4),
    .b(G1),
    .c(G2),
    .y(_166_)
  );
  al_or3fft _488_ (
    .a(_069_),
    .b(_166_),
    .c(_076_),
    .y(_167_)
  );
  al_and3 _489_ (
    .a(G6),
    .b(_167_),
    .c(_141_),
    .y(_168_)
  );
  al_and3fft _490_ (
    .a(\DFF_11.Q ),
    .b(_023_),
    .c(_022_),
    .y(_169_)
  );
  al_ao21 _491_ (
    .a(_000_),
    .b(_072_),
    .c(_068_),
    .y(_170_)
  );
  al_ao21 _492_ (
    .a(_159_),
    .b(_170_),
    .c(_025_),
    .y(_171_)
  );
  al_aoi21ftt _493_ (
    .a(G5),
    .b(G4),
    .c(_075_),
    .y(_172_)
  );
  al_ao21ftf _494_ (
    .a(_172_),
    .b(_171_),
    .c(_148_),
    .y(_173_)
  );
  al_or3ftt _495_ (
    .a(_173_),
    .b(_169_),
    .c(_168_),
    .y(G552)
  );
  al_and3 _496_ (
    .a(G7),
    .b(G10),
    .c(_237_),
    .y(_174_)
  );
  al_and3fft _497_ (
    .a(_059_),
    .b(_037_),
    .c(_104_),
    .y(_175_)
  );
  al_mux2l _498_ (
    .a(G9),
    .b(G11),
    .s(G10),
    .y(_176_)
  );
  al_ao21ftt _499_ (
    .a(_176_),
    .b(_037_),
    .c(_068_),
    .y(_177_)
  );
  al_oai21ttf _500_ (
    .a(_177_),
    .b(_175_),
    .c(_174_),
    .y(_178_)
  );
  al_aoi21ttf _501_ (
    .a(G8),
    .b(G10),
    .c(G7),
    .y(_179_)
  );
  al_ao21 _502_ (
    .a(G10),
    .b(_037_),
    .c(_179_),
    .y(_180_)
  );
  al_and3 _503_ (
    .a(G9),
    .b(\DFF_5.Q ),
    .c(_180_),
    .y(_181_)
  );
  al_ao21 _504_ (
    .a(_178_),
    .b(_129_),
    .c(_181_),
    .y(G547)
  );
  al_nand3 _505_ (
    .a(G11),
    .b(G9),
    .c(_179_),
    .y(_182_)
  );
  al_nor3fft _506_ (
    .a(G11),
    .b(_104_),
    .c(_089_),
    .y(_183_)
  );
  al_oai21 _507_ (
    .a(_043_),
    .b(_037_),
    .c(_183_),
    .y(_184_)
  );
  al_ao21 _508_ (
    .a(_182_),
    .b(_184_),
    .c(_131_),
    .y(_185_)
  );
  al_ao21ftf _509_ (
    .a(\DFF_13.Q ),
    .b(_129_),
    .c(_185_),
    .y(G548)
  );
  al_nand3 _510_ (
    .a(_258_),
    .b(_154_),
    .c(_129_),
    .y(_186_)
  );
  al_nor2ft _511_ (
    .a(G5),
    .b(_159_),
    .y(_187_)
  );
  al_ao21ftf _512_ (
    .a(G4),
    .b(G5),
    .c(_239_),
    .y(_188_)
  );
  al_ao21ftf _513_ (
    .a(G4),
    .b(G3),
    .c(_241_),
    .y(_189_)
  );
  al_nand3fft _514_ (
    .a(_188_),
    .b(_187_),
    .c(_189_),
    .y(_190_)
  );
  al_and3 _515_ (
    .a(G1),
    .b(_136_),
    .c(_046_),
    .y(_191_)
  );
  al_nand3 _516_ (
    .a(_190_),
    .b(_191_),
    .c(_080_),
    .y(_192_)
  );
  al_nand2 _517_ (
    .a(G3),
    .b(G4),
    .y(_193_)
  );
  al_and3 _518_ (
    .a(G2),
    .b(G5),
    .c(_193_),
    .y(_194_)
  );
  al_aoi21ttf _519_ (
    .a(_194_),
    .b(_148_),
    .c(_147_),
    .y(_195_)
  );
  al_nand3 _520_ (
    .a(_192_),
    .b(_195_),
    .c(_186_),
    .y(G549)
  );
  al_and3 _521_ (
    .a(G2),
    .b(G1),
    .c(_122_),
    .y(_196_)
  );
  al_ao21 _522_ (
    .a(_152_),
    .b(_002_),
    .c(_196_),
    .y(_197_)
  );
  al_and3ftt _523_ (
    .a(_023_),
    .b(_197_),
    .c(_022_),
    .y(_198_)
  );
  al_oai21ttf _524_ (
    .a(_036_),
    .b(_049_),
    .c(_198_),
    .y(G530)
  );
  al_nand3 _525_ (
    .a(_033_),
    .b(_047_),
    .c(_041_),
    .y(_199_)
  );
  al_ao21ftf _526_ (
    .a(_146_),
    .b(_066_),
    .c(_199_),
    .y(_200_)
  );
  al_ao21 _527_ (
    .a(G13),
    .b(_066_),
    .c(_245_),
    .y(_201_)
  );
  al_or3fft _528_ (
    .a(G5),
    .b(G9),
    .c(_030_),
    .y(_202_)
  );
  al_inv _529_ (
    .a(G4),
    .y(_203_)
  );
  al_oa21ftt _530_ (
    .a(_250_),
    .b(_113_),
    .c(_203_),
    .y(_204_)
  );
  al_oa21ftf _531_ (
    .a(_202_),
    .b(_204_),
    .c(_068_),
    .y(_205_)
  );
  al_ao21 _532_ (
    .a(_060_),
    .b(_201_),
    .c(_205_),
    .y(_206_)
  );
  al_and2ft _533_ (
    .a(G3),
    .b(_055_),
    .y(_207_)
  );
  al_ao21 _534_ (
    .a(_057_),
    .b(_187_),
    .c(_207_),
    .y(_208_)
  );
  al_or3 _535_ (
    .a(_146_),
    .b(\DFF_14.Q ),
    .c(_135_),
    .y(_209_)
  );
  al_oai21ftt _536_ (
    .a(_208_),
    .b(_199_),
    .c(_209_),
    .y(_210_)
  );
  al_ao21 _537_ (
    .a(_200_),
    .b(_206_),
    .c(_210_),
    .y(_211_)
  );
  al_nand3 _538_ (
    .a(G1),
    .b(_240_),
    .c(_193_),
    .y(_212_)
  );
  al_ao21ttf _539_ (
    .a(G3),
    .b(G1),
    .c(G2),
    .y(_213_)
  );
  al_ao21 _540_ (
    .a(_239_),
    .b(_213_),
    .c(_203_),
    .y(_214_)
  );
  al_nand3 _541_ (
    .a(_074_),
    .b(_212_),
    .c(_214_),
    .y(_215_)
  );
  al_and3 _542_ (
    .a(G0),
    .b(_215_),
    .c(_129_),
    .y(_216_)
  );
  al_ao21 _543_ (
    .a(_042_),
    .b(_211_),
    .c(_216_),
    .y(G532)
  );
  al_and2 _544_ (
    .a(G13),
    .b(_066_),
    .y(_217_)
  );
  al_oa21ttf _545_ (
    .a(G7),
    .b(G9),
    .c(G10),
    .y(_218_)
  );
  al_nand3ftt _546_ (
    .a(_000_),
    .b(_218_),
    .c(_217_),
    .y(_219_)
  );
  al_ao21ttf _547_ (
    .a(_204_),
    .b(_200_),
    .c(_219_),
    .y(_220_)
  );
  al_and2ft _548_ (
    .a(G12),
    .b(G6),
    .y(_221_)
  );
  al_and2 _549_ (
    .a(\DFF_8.Q ),
    .b(\DFF_9.Q ),
    .y(_222_)
  );
  al_nand3 _550_ (
    .a(_076_),
    .b(_222_),
    .c(_024_),
    .y(_223_)
  );
  al_nand3ftt _551_ (
    .a(_026_),
    .b(_245_),
    .c(_218_),
    .y(_224_)
  );
  al_ao21ftf _552_ (
    .a(\DFF_15.Q ),
    .b(_151_),
    .c(_224_),
    .y(_225_)
  );
  al_ao21ftf _553_ (
    .a(_049_),
    .b(_225_),
    .c(_223_),
    .y(_226_)
  );
  al_ao21 _554_ (
    .a(_221_),
    .b(_220_),
    .c(_226_),
    .y(G535)
  );
  al_oa21ftt _555_ (
    .a(_250_),
    .b(_113_),
    .c(_245_),
    .y(_227_)
  );
  al_oa21 _556_ (
    .a(_030_),
    .b(_111_),
    .c(_114_),
    .y(_228_)
  );
  al_or3 _557_ (
    .a(G6),
    .b(_000_),
    .c(_257_),
    .y(_229_)
  );
  al_and3ftt _558_ (
    .a(_227_),
    .b(_229_),
    .c(_228_),
    .y(_230_)
  );
  al_and3fft _559_ (
    .a(_230_),
    .b(_199_),
    .c(_042_),
    .y(_231_)
  );
  al_oa21ftt _560_ (
    .a(G6),
    .b(_250_),
    .c(_263_),
    .y(_232_)
  );
  al_ao21ttf _561_ (
    .a(_227_),
    .b(_217_),
    .c(_232_),
    .y(_233_)
  );
  al_ao21 _562_ (
    .a(\DFF_9.Q ),
    .b(_238_),
    .c(_043_),
    .y(_234_)
  );
  al_and3 _563_ (
    .a(_076_),
    .b(_234_),
    .c(_024_),
    .y(_235_)
  );
  al_ao21 _564_ (
    .a(_083_),
    .b(_233_),
    .c(_235_),
    .y(_236_)
  );
  al_ao21 _565_ (
    .a(G2),
    .b(_236_),
    .c(_231_),
    .y(G537)
  );
  al_and3fft _566_ (
    .a(G4),
    .b(G0),
    .c(_249_),
    .y(\DFF_9.D )
  );
  al_dffl _567_ (
    .clk(CK),
    .d(\DFF_0.D ),
    .q(\DFF_0.Q )
  );
  al_dffl _568_ (
    .clk(CK),
    .d(\DFF_1.D ),
    .q(\DFF_1.Q )
  );
  al_dffl _569_ (
    .clk(CK),
    .d(\DFF_2.D ),
    .q(\DFF_2.Q )
  );
  al_dffl _570_ (
    .clk(CK),
    .d(\DFF_3.D ),
    .q(\DFF_3.Q )
  );
  al_dffl _571_ (
    .clk(CK),
    .d(\DFF_4.D ),
    .q(\DFF_4.Q )
  );
  al_dffl _572_ (
    .clk(CK),
    .d(\DFF_5.D ),
    .q(\DFF_5.Q )
  );
  al_dffl _573_ (
    .clk(CK),
    .d(\DFF_6.D ),
    .q(\DFF_6.Q )
  );
  al_dffl _574_ (
    .clk(CK),
    .d(\DFF_7.D ),
    .q(\DFF_7.Q )
  );
  al_dffl _575_ (
    .clk(CK),
    .d(\DFF_8.D ),
    .q(\DFF_8.Q )
  );
  al_dffl _576_ (
    .clk(CK),
    .d(\DFF_9.D ),
    .q(\DFF_9.Q )
  );
  al_dffl _577_ (
    .clk(CK),
    .d(\DFF_10.D ),
    .q(\DFF_10.Q )
  );
  al_dffl _578_ (
    .clk(CK),
    .d(\DFF_11.D ),
    .q(\DFF_11.Q )
  );
  al_dffl _579_ (
    .clk(CK),
    .d(\DFF_12.D ),
    .q(\DFF_12.Q )
  );
  al_dffl _580_ (
    .clk(CK),
    .d(\DFF_13.D ),
    .q(\DFF_13.Q )
  );
  al_dffl _581_ (
    .clk(CK),
    .d(\DFF_14.D ),
    .q(\DFF_14.Q )
  );
  al_dffl _582_ (
    .clk(CK),
    .d(\DFF_15.D ),
    .q(\DFF_15.Q )
  );
  al_dffl _583_ (
    .clk(CK),
    .d(\DFF_16.D ),
    .q(\DFF_16.Q )
  );
  al_dffl _584_ (
    .clk(CK),
    .d(\DFF_17.D ),
    .q(\DFF_17.Q )
  );
  assign \DFF_0.CK  = CK;
  assign \DFF_1.CK  = CK;
  assign \DFF_10.CK  = CK;
  assign \DFF_11.CK  = CK;
  assign \DFF_12.CK  = CK;
  assign \DFF_13.CK  = CK;
  assign \DFF_14.CK  = CK;
  assign \DFF_15.CK  = CK;
  assign \DFF_16.CK  = CK;
  assign \DFF_17.CK  = CK;
  assign \DFF_2.CK  = CK;
  assign \DFF_3.CK  = CK;
  assign \DFF_4.CK  = CK;
  assign \DFF_5.CK  = CK;
  assign \DFF_6.CK  = CK;
  assign \DFF_7.CK  = CK;
  assign \DFF_8.CK  = CK;
  assign \DFF_9.CK  = CK;
  assign G107 = G0;
  assign G153 = G2;
  assign G165 = G6;
  assign G228 = G3;
  assign G29 = \DFF_0.Q ;
  assign G30 = \DFF_1.Q ;
  assign G31 = \DFF_2.Q ;
  assign G32 = \DFF_3.Q ;
  assign G33 = \DFF_4.Q ;
  assign G334 = G4;
  assign G335 = G1;
  assign G34 = \DFF_5.Q ;
  assign G35 = \DFF_6.Q ;
  assign G36 = \DFF_7.Q ;
  assign G37 = \DFF_8.Q ;
  assign G38 = \DFF_9.Q ;
  assign G39 = \DFF_10.Q ;
  assign G40 = \DFF_11.Q ;
  assign G41 = \DFF_12.Q ;
  assign G42 = \DFF_13.Q ;
  assign G43 = \DFF_14.Q ;
  assign G44 = \DFF_15.Q ;
  assign G45 = \DFF_16.Q ;
  assign G46 = \DFF_17.Q ;
  assign G502 = \DFF_0.D ;
  assign G503 = \DFF_1.D ;
  assign G504 = \DFF_2.D ;
  assign G505 = \DFF_3.D ;
  assign G506 = \DFF_4.D ;
  assign G507 = \DFF_5.D ;
  assign G508 = \DFF_6.D ;
  assign G509 = \DFF_7.D ;
  assign G510 = \DFF_8.D ;
  assign G511 = \DFF_9.D ;
  assign G512 = \DFF_10.D ;
  assign G513 = \DFF_11.D ;
  assign G514 = \DFF_12.D ;
  assign G515 = \DFF_13.D ;
  assign G516 = \DFF_14.D ;
  assign G517 = \DFF_15.D ;
  assign G518 = \DFF_16.D ;
  assign G519 = \DFF_17.D ;
  assign II218 = G5;
  assign II249 = G10;
  assign II374 = G0;
endmodule
