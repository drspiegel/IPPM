
module s9234(GND, VDD, CK, g102, g107, g1290, g1293, g22, g23, g2584, g301, g306, g310, g314, g319, g32, g3222, g36, g3600, g37, g38, g39, g40, g4098, g4099, g41, g4100, g4101, g4102, g4103, g4104, g4105, g4106, g4107, g4108, g4109, g4110, g4112, g4121, g42, g4307, g4321, g44, g4422, g45, g46, g47, g4809, g5137, g5468, g5469, g557, g558, g559, g560, g561, g562, g563, g564, g567, g5692, g6282, g6284, g6360, g6362, g6364, g6366, g6368, g6370, g6372, g6374, g639, g6728, g702, g705, g89, g94, g98);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  input CK;
  wire \DFF_0.CK ;
  wire \DFF_0.D ;
  wire \DFF_0.Q ;
  wire \DFF_1.CK ;
  wire \DFF_10.CK ;
  wire \DFF_10.D ;
  wire \DFF_10.Q ;
  wire \DFF_100.CK ;
  wire \DFF_101.CK ;
  wire \DFF_102.CK ;
  wire \DFF_102.D ;
  wire \DFF_102.Q ;
  wire \DFF_103.CK ;
  wire \DFF_103.D ;
  wire \DFF_103.Q ;
  wire \DFF_104.CK ;
  wire \DFF_105.CK ;
  wire \DFF_105.D ;
  wire \DFF_105.Q ;
  wire \DFF_106.CK ;
  wire \DFF_107.CK ;
  wire \DFF_108.CK ;
  wire \DFF_108.D ;
  wire \DFF_108.Q ;
  wire \DFF_109.CK ;
  wire \DFF_109.D ;
  wire \DFF_109.Q ;
  wire \DFF_11.CK ;
  wire \DFF_11.D ;
  wire \DFF_11.Q ;
  wire \DFF_110.CK ;
  wire \DFF_110.D ;
  wire \DFF_110.Q ;
  wire \DFF_111.CK ;
  wire \DFF_111.D ;
  wire \DFF_111.Q ;
  wire \DFF_112.CK ;
  wire \DFF_113.CK ;
  wire \DFF_113.D ;
  wire \DFF_113.Q ;
  wire \DFF_114.CK ;
  wire \DFF_114.D ;
  wire \DFF_114.Q ;
  wire \DFF_115.CK ;
  wire \DFF_116.CK ;
  wire \DFF_116.D ;
  wire \DFF_116.Q ;
  wire \DFF_117.CK ;
  wire \DFF_117.D ;
  wire \DFF_117.Q ;
  wire \DFF_118.CK ;
  wire \DFF_118.D ;
  wire \DFF_118.Q ;
  wire \DFF_119.CK ;
  wire \DFF_12.CK ;
  wire \DFF_120.CK ;
  wire \DFF_121.CK ;
  wire \DFF_121.D ;
  wire \DFF_121.Q ;
  wire \DFF_122.CK ;
  wire \DFF_122.D ;
  wire \DFF_122.Q ;
  wire \DFF_123.CK ;
  wire \DFF_123.D ;
  wire \DFF_123.Q ;
  wire \DFF_124.CK ;
  wire \DFF_124.D ;
  wire \DFF_124.Q ;
  wire \DFF_125.CK ;
  wire \DFF_125.D ;
  wire \DFF_125.Q ;
  wire \DFF_126.CK ;
  wire \DFF_126.D ;
  wire \DFF_126.Q ;
  wire \DFF_127.CK ;
  wire \DFF_127.D ;
  wire \DFF_127.Q ;
  wire \DFF_128.CK ;
  wire \DFF_128.D ;
  wire \DFF_128.Q ;
  wire \DFF_129.CK ;
  wire \DFF_129.D ;
  wire \DFF_129.Q ;
  wire \DFF_13.CK ;
  wire \DFF_13.D ;
  wire \DFF_13.Q ;
  wire \DFF_130.CK ;
  wire \DFF_131.CK ;
  wire \DFF_131.D ;
  wire \DFF_131.Q ;
  wire \DFF_132.CK ;
  wire \DFF_132.D ;
  wire \DFF_132.Q ;
  wire \DFF_133.CK ;
  wire \DFF_134.CK ;
  wire \DFF_134.D ;
  wire \DFF_134.Q ;
  wire \DFF_135.CK ;
  wire \DFF_135.D ;
  wire \DFF_135.Q ;
  wire \DFF_136.CK ;
  wire \DFF_137.CK ;
  wire \DFF_137.D ;
  wire \DFF_138.CK ;
  wire \DFF_138.D ;
  wire \DFF_138.Q ;
  wire \DFF_139.CK ;
  wire \DFF_139.D ;
  wire \DFF_139.Q ;
  wire \DFF_14.CK ;
  wire \DFF_14.D ;
  wire \DFF_14.Q ;
  wire \DFF_140.CK ;
  wire \DFF_140.D ;
  wire \DFF_140.Q ;
  wire \DFF_141.CK ;
  wire \DFF_141.D ;
  wire \DFF_141.Q ;
  wire \DFF_142.CK ;
  wire \DFF_142.D ;
  wire \DFF_142.Q ;
  wire \DFF_143.CK ;
  wire \DFF_143.D ;
  wire \DFF_143.Q ;
  wire \DFF_144.CK ;
  wire \DFF_144.D ;
  wire \DFF_144.Q ;
  wire \DFF_145.CK ;
  wire \DFF_146.CK ;
  wire \DFF_146.D ;
  wire \DFF_146.Q ;
  wire \DFF_147.CK ;
  wire \DFF_147.D ;
  wire \DFF_147.Q ;
  wire \DFF_148.CK ;
  wire \DFF_148.D ;
  wire \DFF_148.Q ;
  wire \DFF_149.CK ;
  wire \DFF_15.CK ;
  wire \DFF_15.D ;
  wire \DFF_15.Q ;
  wire \DFF_150.CK ;
  wire \DFF_151.CK ;
  wire \DFF_151.D ;
  wire \DFF_151.Q ;
  wire \DFF_152.CK ;
  wire \DFF_152.D ;
  wire \DFF_152.Q ;
  wire \DFF_153.CK ;
  wire \DFF_153.D ;
  wire \DFF_153.Q ;
  wire \DFF_154.CK ;
  wire \DFF_154.D ;
  wire \DFF_154.Q ;
  wire \DFF_155.CK ;
  wire \DFF_156.CK ;
  wire \DFF_156.D ;
  wire \DFF_156.Q ;
  wire \DFF_157.CK ;
  wire \DFF_157.D ;
  wire \DFF_157.Q ;
  wire \DFF_158.CK ;
  wire \DFF_158.D ;
  wire \DFF_158.Q ;
  wire \DFF_159.CK ;
  wire \DFF_16.CK ;
  wire \DFF_160.CK ;
  wire \DFF_161.CK ;
  wire \DFF_161.D ;
  wire \DFF_161.Q ;
  wire \DFF_162.CK ;
  wire \DFF_163.CK ;
  wire \DFF_163.D ;
  wire \DFF_163.Q ;
  wire \DFF_164.CK ;
  wire \DFF_164.D ;
  wire \DFF_164.Q ;
  wire \DFF_165.CK ;
  wire \DFF_166.CK ;
  wire \DFF_166.D ;
  wire \DFF_166.Q ;
  wire \DFF_167.CK ;
  wire \DFF_167.D ;
  wire \DFF_167.Q ;
  wire \DFF_168.CK ;
  wire \DFF_168.D ;
  wire \DFF_168.Q ;
  wire \DFF_169.CK ;
  wire \DFF_169.D ;
  wire \DFF_169.Q ;
  wire \DFF_17.CK ;
  wire \DFF_17.D ;
  wire \DFF_17.Q ;
  wire \DFF_170.CK ;
  wire \DFF_170.D ;
  wire \DFF_170.Q ;
  wire \DFF_171.CK ;
  wire \DFF_172.CK ;
  wire \DFF_172.D ;
  wire \DFF_172.Q ;
  wire \DFF_173.CK ;
  wire \DFF_173.D ;
  wire \DFF_173.Q ;
  wire \DFF_174.CK ;
  wire \DFF_175.CK ;
  wire \DFF_175.D ;
  wire \DFF_175.Q ;
  wire \DFF_176.CK ;
  wire \DFF_176.D ;
  wire \DFF_176.Q ;
  wire \DFF_177.CK ;
  wire \DFF_177.D ;
  wire \DFF_177.Q ;
  wire \DFF_178.CK ;
  wire \DFF_178.D ;
  wire \DFF_178.Q ;
  wire \DFF_179.CK ;
  wire \DFF_179.D ;
  wire \DFF_179.Q ;
  wire \DFF_18.CK ;
  wire \DFF_180.CK ;
  wire \DFF_180.D ;
  wire \DFF_180.Q ;
  wire \DFF_181.CK ;
  wire \DFF_182.CK ;
  wire \DFF_182.D ;
  wire \DFF_182.Q ;
  wire \DFF_183.CK ;
  wire \DFF_183.D ;
  wire \DFF_183.Q ;
  wire \DFF_184.CK ;
  wire \DFF_185.CK ;
  wire \DFF_186.CK ;
  wire \DFF_186.D ;
  wire \DFF_186.Q ;
  wire \DFF_187.CK ;
  wire \DFF_187.D ;
  wire \DFF_187.Q ;
  wire \DFF_188.CK ;
  wire \DFF_188.D ;
  wire \DFF_188.Q ;
  wire \DFF_189.CK ;
  wire \DFF_189.D ;
  wire \DFF_189.Q ;
  wire \DFF_19.CK ;
  wire \DFF_19.D ;
  wire \DFF_19.Q ;
  wire \DFF_190.CK ;
  wire \DFF_190.D ;
  wire \DFF_190.Q ;
  wire \DFF_191.CK ;
  wire \DFF_191.D ;
  wire \DFF_191.Q ;
  wire \DFF_192.CK ;
  wire \DFF_193.CK ;
  wire \DFF_194.CK ;
  wire \DFF_195.CK ;
  wire \DFF_195.D ;
  wire \DFF_195.Q ;
  wire \DFF_196.CK ;
  wire \DFF_196.D ;
  wire \DFF_196.Q ;
  wire \DFF_197.CK ;
  wire \DFF_197.D ;
  wire \DFF_197.Q ;
  wire \DFF_198.CK ;
  wire \DFF_199.CK ;
  wire \DFF_2.CK ;
  wire \DFF_20.CK ;
  wire \DFF_20.D ;
  wire \DFF_20.Q ;
  wire \DFF_200.CK ;
  wire \DFF_200.D ;
  wire \DFF_200.Q ;
  wire \DFF_201.CK ;
  wire \DFF_201.D ;
  wire \DFF_201.Q ;
  wire \DFF_202.CK ;
  wire \DFF_203.CK ;
  wire \DFF_204.CK ;
  wire \DFF_204.D ;
  wire \DFF_204.Q ;
  wire \DFF_205.CK ;
  wire \DFF_205.D ;
  wire \DFF_205.Q ;
  wire \DFF_206.CK ;
  wire \DFF_207.CK ;
  wire \DFF_207.D ;
  wire \DFF_207.Q ;
  wire \DFF_208.CK ;
  wire \DFF_208.D ;
  wire \DFF_208.Q ;
  wire \DFF_209.CK ;
  wire \DFF_209.D ;
  wire \DFF_209.Q ;
  wire \DFF_21.CK ;
  wire \DFF_21.D ;
  wire \DFF_21.Q ;
  wire \DFF_210.CK ;
  wire \DFF_22.CK ;
  wire \DFF_23.CK ;
  wire \DFF_23.D ;
  wire \DFF_23.Q ;
  wire \DFF_24.CK ;
  wire \DFF_24.D ;
  wire \DFF_24.Q ;
  wire \DFF_25.CK ;
  wire \DFF_25.D ;
  wire \DFF_25.Q ;
  wire \DFF_26.CK ;
  wire \DFF_26.D ;
  wire \DFF_26.Q ;
  wire \DFF_27.CK ;
  wire \DFF_27.D ;
  wire \DFF_27.Q ;
  wire \DFF_28.CK ;
  wire \DFF_28.D ;
  wire \DFF_28.Q ;
  wire \DFF_29.CK ;
  wire \DFF_3.CK ;
  wire \DFF_3.D ;
  wire \DFF_3.Q ;
  wire \DFF_30.CK ;
  wire \DFF_30.D ;
  wire \DFF_30.Q ;
  wire \DFF_31.CK ;
  wire \DFF_32.CK ;
  wire \DFF_33.CK ;
  wire \DFF_33.D ;
  wire \DFF_33.Q ;
  wire \DFF_34.CK ;
  wire \DFF_35.CK ;
  wire \DFF_35.D ;
  wire \DFF_35.Q ;
  wire \DFF_36.CK ;
  wire \DFF_36.D ;
  wire \DFF_36.Q ;
  wire \DFF_37.CK ;
  wire \DFF_37.D ;
  wire \DFF_37.Q ;
  wire \DFF_38.CK ;
  wire \DFF_38.D ;
  wire \DFF_38.Q ;
  wire \DFF_39.CK ;
  wire \DFF_4.CK ;
  wire \DFF_4.D ;
  wire \DFF_4.Q ;
  wire \DFF_40.CK ;
  wire \DFF_40.D ;
  wire \DFF_40.Q ;
  wire \DFF_41.CK ;
  wire \DFF_41.D ;
  wire \DFF_41.Q ;
  wire \DFF_42.CK ;
  wire \DFF_42.D ;
  wire \DFF_42.Q ;
  wire \DFF_43.CK ;
  wire \DFF_43.D ;
  wire \DFF_43.Q ;
  wire \DFF_44.CK ;
  wire \DFF_44.D ;
  wire \DFF_44.Q ;
  wire \DFF_45.CK ;
  wire \DFF_46.CK ;
  wire \DFF_46.D ;
  wire \DFF_46.Q ;
  wire \DFF_47.CK ;
  wire \DFF_47.D ;
  wire \DFF_47.Q ;
  wire \DFF_48.CK ;
  wire \DFF_48.D ;
  wire \DFF_48.Q ;
  wire \DFF_49.CK ;
  wire \DFF_5.CK ;
  wire \DFF_5.D ;
  wire \DFF_5.Q ;
  wire \DFF_50.CK ;
  wire \DFF_50.D ;
  wire \DFF_50.Q ;
  wire \DFF_51.CK ;
  wire \DFF_51.D ;
  wire \DFF_51.Q ;
  wire \DFF_52.CK ;
  wire \DFF_52.D ;
  wire \DFF_52.Q ;
  wire \DFF_53.CK ;
  wire \DFF_53.D ;
  wire \DFF_53.Q ;
  wire \DFF_54.CK ;
  wire \DFF_55.CK ;
  wire \DFF_55.D ;
  wire \DFF_55.Q ;
  wire \DFF_56.CK ;
  wire \DFF_56.D ;
  wire \DFF_56.Q ;
  wire \DFF_57.CK ;
  wire \DFF_57.D ;
  wire \DFF_57.Q ;
  wire \DFF_58.CK ;
  wire \DFF_58.D ;
  wire \DFF_58.Q ;
  wire \DFF_59.CK ;
  wire \DFF_59.D ;
  wire \DFF_59.Q ;
  wire \DFF_6.CK ;
  wire \DFF_6.D ;
  wire \DFF_6.Q ;
  wire \DFF_60.CK ;
  wire \DFF_60.D ;
  wire \DFF_60.Q ;
  wire \DFF_61.CK ;
  wire \DFF_61.D ;
  wire \DFF_61.Q ;
  wire \DFF_62.CK ;
  wire \DFF_63.CK ;
  wire \DFF_63.D ;
  wire \DFF_63.Q ;
  wire \DFF_64.CK ;
  wire \DFF_64.D ;
  wire \DFF_64.Q ;
  wire \DFF_65.CK ;
  wire \DFF_66.CK ;
  wire \DFF_66.D ;
  wire \DFF_66.Q ;
  wire \DFF_67.CK ;
  wire \DFF_68.CK ;
  wire \DFF_68.D ;
  wire \DFF_68.Q ;
  wire \DFF_69.CK ;
  wire \DFF_69.D ;
  wire \DFF_69.Q ;
  wire \DFF_7.CK ;
  wire \DFF_7.D ;
  wire \DFF_7.Q ;
  wire \DFF_70.CK ;
  wire \DFF_70.D ;
  wire \DFF_70.Q ;
  wire \DFF_71.CK ;
  wire \DFF_72.CK ;
  wire \DFF_72.D ;
  wire \DFF_72.Q ;
  wire \DFF_73.CK ;
  wire \DFF_73.D ;
  wire \DFF_73.Q ;
  wire \DFF_74.CK ;
  wire \DFF_74.D ;
  wire \DFF_74.Q ;
  wire \DFF_75.CK ;
  wire \DFF_75.D ;
  wire \DFF_75.Q ;
  wire \DFF_76.CK ;
  wire \DFF_76.D ;
  wire \DFF_76.Q ;
  wire \DFF_77.CK ;
  wire \DFF_77.D ;
  wire \DFF_77.Q ;
  wire \DFF_78.CK ;
  wire \DFF_78.D ;
  wire \DFF_78.Q ;
  wire \DFF_79.CK ;
  wire \DFF_79.D ;
  wire \DFF_79.Q ;
  wire \DFF_8.CK ;
  wire \DFF_80.CK ;
  wire \DFF_80.D ;
  wire \DFF_80.Q ;
  wire \DFF_81.CK ;
  wire \DFF_81.D ;
  wire \DFF_81.Q ;
  wire \DFF_82.CK ;
  wire \DFF_82.D ;
  wire \DFF_82.Q ;
  wire \DFF_83.CK ;
  wire \DFF_83.D ;
  wire \DFF_83.Q ;
  wire \DFF_84.CK ;
  wire \DFF_84.D ;
  wire \DFF_84.Q ;
  wire \DFF_85.CK ;
  wire \DFF_85.D ;
  wire \DFF_85.Q ;
  wire \DFF_86.CK ;
  wire \DFF_87.CK ;
  wire \DFF_87.D ;
  wire \DFF_87.Q ;
  wire \DFF_88.CK ;
  wire \DFF_88.D ;
  wire \DFF_88.Q ;
  wire \DFF_89.CK ;
  wire \DFF_89.D ;
  wire \DFF_89.Q ;
  wire \DFF_9.CK ;
  wire \DFF_9.D ;
  wire \DFF_9.Q ;
  wire \DFF_90.CK ;
  wire \DFF_90.D ;
  wire \DFF_90.Q ;
  wire \DFF_91.CK ;
  wire \DFF_92.CK ;
  wire \DFF_92.D ;
  wire \DFF_92.Q ;
  wire \DFF_93.CK ;
  wire \DFF_93.D ;
  wire \DFF_93.Q ;
  wire \DFF_94.CK ;
  wire \DFF_94.D ;
  wire \DFF_94.Q ;
  wire \DFF_95.CK ;
  wire \DFF_95.D ;
  wire \DFF_95.Q ;
  wire \DFF_96.CK ;
  wire \DFF_96.D ;
  wire \DFF_96.Q ;
  wire \DFF_97.CK ;
  wire \DFF_98.CK ;
  wire \DFF_98.D ;
  wire \DFF_98.Q ;
  wire \DFF_99.CK ;
  wire \DFF_99.D ;
  wire \DFF_99.Q ;
  input GND;
  wire I2029;
  wire I2033;
  wire I2165;
  wire I2172;
  wire I2290;
  wire I2293;
  wire I2296;
  wire I2306;
  wire I2312;
  wire I2321;
  wire I2364;
  wire I2370;
  wire I2373;
  wire I2379;
  wire I2388;
  wire I2445;
  wire I2449;
  wire I2453;
  wire I2460;
  wire I2464;
  wire I2473;
  wire I2476;
  wire I2479;
  wire I2521;
  wire I2537;
  wire I2552;
  wire I2584;
  wire I2596;
  wire I2608;
  wire I2614;
  wire I2627;
  wire I2630;
  wire I2635;
  wire I2638;
  wire I2643;
  wire I2716;
  wire I2731;
  wire I2735;
  wire I2753;
  wire I2756;
  wire I2773;
  wire I2776;
  wire I2802;
  wire I2805;
  wire I2821;
  wire I2825;
  wire I2839;
  wire I2867;
  wire I2877;
  wire I2880;
  wire I2883;
  wire I2887;
  wire I2890;
  wire I2907;
  wire I2910;
  wire I2916;
  wire I2929;
  wire I2940;
  wire I2943;
  wire I2946;
  wire I2952;
  wire I2955;
  wire I2961;
  wire I2982;
  wire I2992;
  wire I2995;
  wire I3004;
  wire I3007;
  wire I3016;
  wire I3019;
  wire I3022;
  wire I3025;
  wire I3037;
  wire I3040;
  wire I3047;
  wire I3050;
  wire I3062;
  wire I3065;
  wire I3068;
  wire I3074;
  wire I3077;
  wire I3083;
  wire I3086;
  wire I3093;
  wire I3096;
  wire I3102;
  wire I3105;
  wire I3112;
  wire I3137;
  wire I3140;
  wire I3144;
  wire I3152;
  wire I3198;
  wire I3202;
  wire I3206;
  wire I3215;
  wire I3251;
  wire I3255;
  wire I3268;
  wire I3278;
  wire I3284;
  wire I3288;
  wire I3291;
  wire I3294;
  wire I3298;
  wire I3301;
  wire I3304;
  wire I3307;
  wire I3313;
  wire I3316;
  wire I3325;
  wire I3434;
  wire I3452;
  wire I3462;
  wire I3471;
  wire I3474;
  wire I3478;
  wire I3481;
  wire I3485;
  wire I3488;
  wire I3493;
  wire I3496;
  wire I3499;
  wire I3502;
  wire I3505;
  wire I3509;
  wire I3513;
  wire I3516;
  wire I3519;
  wire I3522;
  wire I3525;
  wire I3534;
  wire I3537;
  wire I3543;
  wire I3550;
  wire I3553;
  wire I3556;
  wire I3563;
  wire I3569;
  wire I3572;
  wire I3575;
  wire I3578;
  wire I3581;
  wire I3587;
  wire I3590;
  wire I3593;
  wire I3596;
  wire I3599;
  wire I3602;
  wire I3608;
  wire I3614;
  wire I3617;
  wire I3620;
  wire I3623;
  wire I3632;
  wire I3635;
  wire I3638;
  wire I3641;
  wire I3650;
  wire I3653;
  wire I3656;
  wire I3659;
  wire I3665;
  wire I3672;
  wire I3675;
  wire I3681;
  wire I3711;
  wire I3714;
  wire I3726;
  wire I3729;
  wire I3733;
  wire I3736;
  wire I3746;
  wire I3755;
  wire I3758;
  wire I3767;
  wire I3770;
  wire I3779;
  wire I3782;
  wire I3785;
  wire I3797;
  wire I3800;
  wire I3808;
  wire I3811;
  wire I3823;
  wire I3826;
  wire I3836;
  wire I3840;
  wire I3843;
  wire I3855;
  wire I3861;
  wire I3868;
  wire I3871;
  wire I3883;
  wire I3890;
  wire I4019;
  wire I4031;
  wire I4170;
  wire I4189;
  wire I4192;
  wire I4217;
  wire I4220;
  wire I4226;
  wire I4240;
  wire I4243;
  wire I4249;
  wire I4252;
  wire I4258;
  wire I4261;
  wire I4267;
  wire I4270;
  wire I4276;
  wire I4282;
  wire I4285;
  wire I4294;
  wire I4297;
  wire I4303;
  wire I4306;
  wire I4309;
  wire I4312;
  wire I4318;
  wire I4321;
  wire I4324;
  wire I4327;
  wire I4331;
  wire I4337;
  wire I4340;
  wire I4343;
  wire I4347;
  wire I4354;
  wire I4358;
  wire I4362;
  wire I4371;
  wire I4398;
  wire I4410;
  wire I4414;
  wire I4424;
  wire I4468;
  wire I4903;
  wire I5337;
  wire I5415;
  wire I5418;
  wire I5542;
  wire I5929;
  input VDD;
  wire g1;
  wire g10;
  wire g1001;
  wire g1006;
  wire g1011;
  wire g1017;
  input g102;
  wire g1030;
  wire g1049;
  input g107;
  wire g1076;
  wire g1088;
  wire g1094;
  wire g11;
  wire g1101;
  wire g1106;
  wire g1107;
  wire g1108;
  wire g1109;
  wire g1110;
  wire g1111;
  wire g1113;
  wire g1114;
  wire g1116;
  wire g1119;
  wire g1122;
  wire g1123;
  wire g1142;
  wire g1143;
  wire g1156;
  wire g1160;
  wire g1161;
  wire g1173;
  wire g1176;
  wire g1177;
  wire g1189;
  wire g1190;
  wire g1193;
  wire g1203;
  wire g1209;
  wire g1219;
  wire g1220;
  wire g1222;
  wire g1232;
  wire g1233;
  wire g1236;
  wire g1246;
  wire g1249;
  wire g1256;
  wire g1257;
  wire g1263;
  wire g1267;
  wire g1270;
  wire g1273;
  wire g1274;
  wire g1275;
  wire g1276;
  wire g1279;
  wire g1282;
  wire g1283;
  wire g1284;
  wire g1285;
  wire g1286;
  wire g1287;
  wire g1288;
  wire g1289;
  output g1290;
  wire g1291;
  wire g1292;
  output g1293;
  wire g1294;
  wire g1318;
  wire g1320;
  wire g1321;
  wire g1322;
  wire g1323;
  wire g1324;
  wire g1325;
  wire g1327;
  wire g1328;
  wire g1329;
  wire g1330;
  wire g1331;
  wire g1332;
  wire g1333;
  wire g1334;
  wire g1335;
  wire g1337;
  wire g1338;
  wire g1339;
  wire g1340;
  wire g1341;
  wire g1344;
  wire g1345;
  wire g1348;
  wire g1352;
  wire g1355;
  wire g1363;
  wire g1366;
  wire g1372;
  wire g1375;
  wire g1378;
  wire g1381;
  wire g1384;
  wire g1391;
  wire g1395;
  wire g14;
  wire g1450;
  wire g1461;
  wire g1472;
  wire g1477;
  wire g1480;
  wire g1498;
  wire g15;
  wire g1503;
  wire g1504;
  wire g1513;
  wire g1519;
  wire g1528;
  wire g1533;
  wire g1539;
  wire g1542;
  wire g1549;
  wire g1556;
  wire g1559;
  wire g1586;
  wire g1587;
  wire g1593;
  wire g1594;
  wire g1608;
  wire g1623;
  wire g1631;
  wire g1636;
  wire g1640;
  wire g1641;
  wire g1643;
  wire g1644;
  wire g1645;
  wire g1646;
  wire g1647;
  wire g1648;
  wire g1649;
  wire g1653;
  wire g1654;
  wire g1655;
  wire g1659;
  wire g1660;
  wire g1664;
  wire g1665;
  wire g1670;
  wire g1671;
  wire g1673;
  wire g1674;
  wire g1678;
  wire g1679;
  wire g1681;
  wire g1684;
  wire g1685;
  wire g1688;
  wire g1692;
  wire g1696;
  wire g1699;
  wire g1703;
  wire g1711;
  wire g1721;
  wire g1724;
  wire g1726;
  wire g1732;
  wire g1733;
  wire g1734;
  wire g1735;
  wire g1739;
  wire g1747;
  wire g1748;
  wire g1759;
  wire g1760;
  wire g1761;
  wire g1762;
  wire g1771;
  wire g1772;
  wire g1773;
  wire g1774;
  wire g1775;
  wire g1781;
  wire g1782;
  wire g1783;
  wire g1787;
  wire g1788;
  wire g1789;
  wire g1790;
  wire g1791;
  wire g1792;
  wire g18;
  wire g1802;
  wire g1805;
  wire g1806;
  wire g1807;
  wire g1811;
  wire g1812;
  wire g1813;
  wire g1814;
  wire g1819;
  wire g1820;
  wire g1821;
  wire g1823;
  wire g1824;
  wire g1825;
  wire g1830;
  wire g1831;
  wire g1832;
  wire g1833;
  wire g1834;
  wire g1835;
  wire g1836;
  wire g1837;
  wire g1841;
  wire g1846;
  wire g1848;
  wire g1849;
  wire g1852;
  wire g1854;
  wire g1858;
  wire g1875;
  wire g1884;
  wire g1891;
  wire g1894;
  wire g1899;
  wire g19;
  wire g1902;
  wire g1911;
  wire g1914;
  wire g1925;
  wire g1928;
  wire g1931;
  wire g1937;
  wire g1947;
  wire g1950;
  wire g1960;
  wire g1969;
  wire g197;
  wire g1979;
  wire g1988;
  wire g1998;
  wire g2;
  wire g2004;
  wire g204;
  wire g2040;
  wire g2041;
  wire g2044;
  wire g205;
  wire g206;
  wire g207;
  wire g208;
  wire g2086;
  wire g2088;
  wire g209;
  wire g2090;
  wire g2096;
  wire g2097;
  wire g210;
  wire g2102;
  wire g2103;
  wire g2108;
  wire g2109;
  wire g211;
  wire g2117;
  wire g2118;
  wire g212;
  wire g2134;
  wire g2135;
  wire g2154;
  wire g2155;
  wire g2158;
  wire g2172;
  wire g2173;
  wire g2174;
  wire g2175;
  wire g2176;
  wire g2177;
  wire g2178;
  wire g2179;
  wire g218;
  wire g2194;
  wire g2195;
  wire g2196;
  wire g2197;
  input g22;
  wire g2212;
  wire g2213;
  wire g2214;
  wire g2215;
  wire g2230;
  wire g2231;
  wire g2232;
  wire g2233;
  wire g2234;
  wire g224;
  wire g2241;
  wire g2242;
  wire g2243;
  wire g2244;
  wire g2245;
  wire g2252;
  wire g2253;
  wire g2254;
  wire g2256;
  wire g2264;
  wire g2265;
  wire g2268;
  wire g2275;
  wire g2276;
  wire g2283;
  wire g2284;
  wire g2293;
  wire g2295;
  input g23;
  wire g230;
  wire g2308;
  wire g2312;
  wire g2315;
  wire g2316;
  wire g2317;
  wire g2320;
  wire g2324;
  wire g2327;
  wire g2333;
  wire g2343;
  wire g2347;
  wire g2357;
  wire g236;
  wire g2361;
  wire g2370;
  wire g2378;
  wire g2390;
  wire g2397;
  wire g24;
  wire g2405;
  wire g2408;
  wire g242;
  wire g2422;
  wire g2430;
  wire g2433;
  wire g2436;
  wire g2449;
  wire g2457;
  wire g2460;
  wire g2473;
  wire g248;
  wire g2481;
  wire g2484;
  wire g2497;
  wire g25;
  wire g2505;
  wire g2518;
  wire g2524;
  wire g254;
  wire g2544;
  wire g2550;
  wire g2554;
  wire g2574;
  wire g2575;
  wire g2576;
  wire g2580;
  wire g2581;
  output g2584;
  wire g2586;
  wire g2587;
  wire g2588;
  wire g2591;
  wire g2594;
  wire g2599;
  wire g260;
  wire g2604;
  wire g2609;
  wire g2612;
  wire g2618;
  wire g2619;
  wire g2622;
  wire g2631;
  wire g2634;
  wire g2644;
  wire g2647;
  wire g2650;
  wire g266;
  wire g2660;
  wire g2663;
  wire g2670;
  wire g2672;
  wire g2675;
  wire g2678;
  wire g2686;
  wire g2688;
  wire g269;
  wire g2691;
  wire g2701;
  wire g2705;
  wire g2706;
  wire g2709;
  wire g2712;
  wire g2722;
  wire g2726;
  wire g2727;
  wire g2734;
  wire g2738;
  wire g2739;
  wire g2740;
  wire g2743;
  wire g2744;
  wire g2748;
  wire g2752;
  wire g2753;
  wire g2754;
  wire g2755;
  wire g2756;
  wire g276;
  wire g2760;
  wire g2764;
  wire g2765;
  wire g2766;
  wire g2767;
  wire g2768;
  wire g277;
  wire g2772;
  wire g2776;
  wire g2777;
  wire g2778;
  wire g2779;
  wire g278;
  wire g2783;
  wire g2787;
  wire g2788;
  wire g2789;
  wire g279;
  wire g2790;
  wire g2792;
  wire g2796;
  wire g28;
  wire g280;
  wire g2800;
  wire g2801;
  wire g2802;
  wire g2803;
  wire g2805;
  wire g2806;
  wire g2809;
  wire g281;
  wire g2813;
  wire g2814;
  wire g2817;
  wire g2818;
  wire g2819;
  wire g282;
  wire g2820;
  wire g2822;
  wire g2826;
  wire g2827;
  wire g2828;
  wire g2829;
  wire g283;
  wire g2830;
  wire g2835;
  wire g2836;
  wire g2837;
  wire g2838;
  wire g2839;
  wire g284;
  wire g2840;
  wire g2841;
  wire g2845;
  wire g285;
  wire g2859;
  wire g286;
  wire g2861;
  wire g2864;
  wire g2866;
  wire g2867;
  wire g287;
  wire g2871;
  wire g2872;
  wire g2875;
  wire g2876;
  wire g288;
  wire g2883;
  wire g2884;
  wire g2885;
  wire g2886;
  wire g2888;
  wire g2889;
  wire g289;
  wire g2892;
  wire g2893;
  wire g29;
  wire g290;
  wire g2904;
  wire g2905;
  wire g291;
  wire g2912;
  wire g292;
  wire g293;
  wire g2945;
  wire g2967;
  wire g297;
  wire g2974;
  wire g2975;
  wire g2998;
  wire g3;
  wire g3001;
  input g301;
  wire g3016;
  wire g3022;
  wire g3031;
  wire g3040;
  wire g3043;
  wire g3052;
  wire g3054;
  input g306;
  wire g3063;
  wire g3064;
  wire g3073;
  wire g3082;
  wire g3093;
  input g310;
  wire g3104;
  wire g3118;
  wire g3128;
  wire g3136;
  input g314;
  wire g3150;
  wire g3158;
  wire g3162;
  wire g3173;
  wire g3177;
  wire g3183;
  wire g3187;
  input g319;
  wire g3192;
  wire g3196;
  input g32;
  wire g3200;
  wire g3204;
  wire g3209;
  wire g3212;
  wire g3216;
  wire g3219;
  output g3222;
  wire g3224;
  wire g3225;
  wire g3226;
  wire g3227;
  wire g3228;
  wire g3229;
  wire g3230;
  wire g3231;
  wire g3232;
  wire g3233;
  wire g3234;
  wire g3235;
  wire g3236;
  wire g3237;
  wire g3238;
  wire g3239;
  wire g3240;
  wire g3241;
  wire g3242;
  wire g3247;
  wire g3259;
  wire g3263;
  wire g3267;
  wire g3271;
  wire g3284;
  wire g3289;
  wire g3291;
  wire g3297;
  wire g3299;
  wire g33;
  wire g3306;
  wire g3308;
  wire g3320;
  wire g3322;
  wire g3331;
  wire g3332;
  wire g3342;
  wire g3343;
  wire g3354;
  wire g3355;
  wire g3363;
  wire g3364;
  wire g3370;
  wire g3440;
  wire g3451;
  wire g3452;
  wire g3453;
  wire g3454;
  wire g3455;
  wire g3456;
  wire g3457;
  wire g3458;
  wire g3459;
  wire g3460;
  wire g3462;
  wire g3463;
  wire g3477;
  wire g3478;
  wire g3482;
  wire g3483;
  wire g3486;
  wire g3488;
  wire g3491;
  wire g3527;
  wire g3534;
  wire g3537;
  wire g3541;
  wire g3545;
  wire g3546;
  wire g3557;
  wire g3559;
  wire g3564;
  wire g3567;
  wire g3571;
  wire g3589;
  wire g3593;
  wire g3599;
  input g36;
  output g3600;
  wire g3601;
  wire g3604;
  wire g3612;
  wire g3638;
  wire g3673;
  input g37;
  wire g3705;
  wire g3710;
  wire g3714;
  wire g3719;
  wire g3766;
  wire g3768;
  wire g3771;
  wire g3783;
  wire g3787;
  input g38;
  wire g3803;
  wire g3807;
  wire g3814;
  wire g3828;
  wire g3832;
  wire g3834;
  wire g3835;
  wire g3836;
  wire g3838;
  wire g3839;
  wire g3840;
  wire g3844;
  wire g3846;
  wire g3847;
  wire g3848;
  wire g3852;
  wire g3853;
  wire g3854;
  wire g3859;
  wire g3860;
  wire g3861;
  wire g3866;
  wire g3867;
  wire g3874;
  wire g3875;
  wire g3876;
  wire g3881;
  wire g3882;
  wire g3885;
  input g39;
  wire g3910;
  wire g3922;
  wire g3932;
  wire g3940;
  wire g3952;
  wire g3960;
  wire g3962;
  wire g3963;
  wire g3967;
  wire g3969;
  wire g3970;
  wire g3975;
  wire g3976;
  wire g3980;
  wire g3984;
  input g40;
  wire g4014;
  wire g4016;
  wire g402;
  wire g4034;
  wire g4036;
  wire g4040;
  wire g406;
  output g4098;
  output g4099;
  input g41;
  wire g410;
  output g4100;
  output g4101;
  output g4102;
  output g4103;
  output g4104;
  output g4105;
  output g4106;
  output g4107;
  output g4108;
  output g4109;
  output g4110;
  output g4112;
  output g4121;
  wire g4122;
  wire g4123;
  wire g4124;
  wire g4125;
  wire g4126;
  wire g4127;
  wire g4128;
  wire g4129;
  wire g4130;
  wire g4131;
  wire g4132;
  wire g4133;
  wire g4134;
  wire g4135;
  wire g4136;
  wire g4137;
  wire g4138;
  wire g4139;
  wire g414;
  wire g4140;
  wire g4141;
  wire g4142;
  wire g4143;
  wire g4144;
  wire g4145;
  wire g4146;
  wire g4147;
  wire g4148;
  wire g4149;
  wire g4150;
  wire g4152;
  wire g4153;
  wire g4157;
  wire g418;
  wire g4194;
  input g42;
  wire g4213;
  wire g4219;
  wire g422;
  wire g4228;
  wire g4249;
  wire g426;
  wire g4299;
  wire g43;
  wire g430;
  output g4307;
  wire g4308;
  wire g4320;
  output g4321;
  wire g4322;
  wire g434;
  wire g4343;
  wire g4350;
  wire g437;
  input g44;
  wire g441;
  output g4422;
  wire g4423;
  wire g4424;
  wire g4425;
  wire g4426;
  wire g4430;
  wire g4433;
  wire g4434;
  wire g4436;
  wire g4438;
  wire g4440;
  wire g4441;
  wire g4443;
  wire g4444;
  wire g4446;
  wire g4447;
  wire g445;
  wire g4450;
  wire g4451;
  wire g4454;
  wire g4455;
  wire g4458;
  wire g4460;
  wire g449;
  wire g4492;
  input g45;
  wire g4501;
  wire g4514;
  wire g4519;
  wire g453;
  wire g4562;
  wire g457;
  input g46;
  wire g4603;
  wire g4609;
  wire g461;
  wire g4644;
  wire g465;
  wire g4657;
  wire g4658;
  wire g4659;
  wire g4687;
  wire g4692;
  wire g4699;
  input g47;
  wire g4700;
  wire g4702;
  wire g4703;
  wire g4704;
  wire g4705;
  wire g4706;
  wire g4707;
  wire g471;
  wire g4711;
  wire g4712;
  wire g4714;
  wire g4715;
  wire g4718;
  wire g4719;
  wire g4721;
  wire g4758;
  wire g4761;
  wire g4765;
  wire g478;
  wire g4781;
  wire g4798;
  wire g48;
  output g4809;
  wire g4810;
  wire g4822;
  wire g4823;
  wire g4824;
  wire g4841;
  wire g4842;
  wire g4843;
  wire g4844;
  wire g4845;
  wire g4846;
  wire g4847;
  wire g4848;
  wire g4849;
  wire g485;
  wire g4850;
  wire g4851;
  wire g4852;
  wire g4853;
  wire g4854;
  wire g4855;
  wire g4856;
  wire g4857;
  wire g4858;
  wire g486;
  wire g4871;
  wire g4872;
  wire g489;
  wire g492;
  wire g496;
  wire g500;
  wire g5010;
  wire g5017;
  wire g5019;
  wire g504;
  wire g5051;
  wire g508;
  wire g5089;
  wire g5110;
  wire g512;
  wire g5135;
  wire g5136;
  output g5137;
  wire g5147;
  wire g5148;
  wire g5149;
  wire g5151;
  wire g516;
  wire g5167;
  wire g520;
  wire g5219;
  wire g5230;
  wire g5231;
  wire g524;
  wire g5273;
  wire g528;
  wire g5307;
  wire g5314;
  wire g5315;
  wire g5316;
  wire g532;
  wire g5328;
  wire g5329;
  wire g5330;
  wire g5355;
  wire g5358;
  wire g536;
  wire g5375;
  wire g5383;
  wire g5385;
  wire g5386;
  wire g5387;
  wire g541;
  wire g5432;
  wire g545;
  wire g5466;
  output g5468;
  output g5469;
  wire g548;
  wire g5489;
  wire g5490;
  wire g5491;
  wire g551;
  wire g5531;
  wire g5532;
  wire g5533;
  wire g5534;
  wire g5535;
  wire g554;
  wire g5540;
  input g557;
  wire g5579;
  input g558;
  wire g5580;
  wire g5581;
  wire g5582;
  wire g5584;
  wire g5587;
  input g559;
  wire g5590;
  wire g5593;
  input g560;
  input g561;
  input g562;
  wire g5622;
  wire g5624;
  wire g5625;
  wire g5626;
  wire g5627;
  wire g5628;
  wire g5629;
  input g563;
  wire g5630;
  input g564;
  wire g5645;
  input g567;
  output g5692;
  wire g5702;
  wire g5705;
  wire g5708;
  wire g571;
  wire g5711;
  wire g5714;
  wire g5717;
  wire g5720;
  wire g5723;
  wire g574;
  wire g5751;
  wire g5752;
  wire g5773;
  wire g5774;
  wire g578;
  wire g582;
  wire g586;
  wire g5875;
  wire g5876;
  wire g5877;
  wire g5878;
  wire g5879;
  wire g590;
  wire g5917;
  wire g5918;
  wire g5919;
  wire g5920;
  wire g5921;
  wire g5922;
  wire g5923;
  wire g5924;
  wire g594;
  wire g598;
  wire g6;
  wire g602;
  wire g6032;
  wire g606;
  wire g610;
  wire g6100;
  wire g6101;
  wire g6102;
  wire g6103;
  wire g6104;
  wire g6105;
  wire g6106;
  wire g6107;
  wire g6110;
  wire g613;
  wire g6137;
  wire g6142;
  wire g616;
  wire g6167;
  wire g6170;
  wire g6173;
  wire g6176;
  wire g6179;
  wire g6182;
  wire g6185;
  wire g6189;
  wire g619;
  wire g622;
  wire g625;
  wire g628;
  output g6282;
  wire g6283;
  output g6284;
  wire g6285;
  wire g6286;
  wire g6287;
  wire g6289;
  wire g6290;
  wire g6291;
  wire g6292;
  wire g6293;
  wire g6294;
  wire g6295;
  wire g6296;
  wire g6297;
  wire g6298;
  wire g6299;
  wire g6300;
  wire g6301;
  wire g6303;
  wire g6304;
  wire g6307;
  wire g6309;
  wire g631;
  wire g6310;
  wire g6312;
  wire g634;
  output g6360;
  wire g6361;
  output g6362;
  wire g6363;
  output g6364;
  wire g6365;
  output g6366;
  wire g6367;
  output g6368;
  wire g6369;
  output g6370;
  wire g6371;
  output g6372;
  wire g6373;
  output g6374;
  wire g6375;
  wire g638;
  input g639;
  wire g6407;
  wire g6410;
  wire g6411;
  wire g6412;
  wire g6413;
  wire g6414;
  wire g6415;
  wire g6416;
  wire g6417;
  wire g6418;
  wire g6419;
  wire g642;
  wire g6420;
  wire g6421;
  wire g6422;
  wire g6423;
  wire g6424;
  wire g6425;
  wire g6426;
  wire g6428;
  wire g6431;
  wire g6434;
  wire g6437;
  wire g6441;
  wire g646;
  wire g6479;
  wire g6480;
  wire g6481;
  wire g6482;
  wire g6483;
  wire g6485;
  wire g6497;
  wire g6498;
  wire g6499;
  wire g650;
  wire g6500;
  wire g6501;
  wire g6502;
  wire g6503;
  wire g6504;
  wire g6505;
  wire g6506;
  wire g6507;
  wire g6508;
  wire g6509;
  wire g6510;
  wire g6511;
  wire g6512;
  wire g6515;
  wire g6516;
  wire g6519;
  wire g6521;
  wire g6523;
  wire g6524;
  wire g6525;
  wire g6526;
  wire g6527;
  wire g6528;
  wire g6529;
  wire g6530;
  wire g6531;
  wire g6532;
  wire g654;
  wire g6574;
  wire g6575;
  wire g6576;
  wire g6577;
  wire g6578;
  wire g6579;
  wire g658;
  wire g6580;
  wire g6581;
  wire g6591;
  wire g6592;
  wire g6593;
  wire g6594;
  wire g6595;
  wire g6596;
  wire g6597;
  wire g6598;
  wire g6599;
  wire g6600;
  wire g6601;
  wire g6602;
  wire g662;
  wire g663;
  wire g664;
  wire g665;
  wire g6658;
  wire g666;
  wire g667;
  wire g668;
  wire g6684;
  wire g6685;
  wire g6686;
  wire g6687;
  wire g6688;
  wire g6689;
  wire g669;
  wire g6690;
  wire g6691;
  wire g6694;
  wire g6695;
  wire g6696;
  wire g6697;
  wire g6698;
  wire g6699;
  wire g6700;
  wire g6701;
  wire g6702;
  wire g6704;
  wire g6711;
  wire g672;
  wire g6720;
  wire g6721;
  wire g6722;
  wire g6723;
  wire g6724;
  wire g6725;
  wire g6726;
  wire g6727;
  output g6728;
  wire g6729;
  wire g6730;
  wire g6743;
  wire g6744;
  wire g6745;
  wire g675;
  wire g676;
  wire g677;
  wire g6774;
  wire g6778;
  wire g678;
  wire g6785;
  wire g6786;
  wire g6787;
  wire g6788;
  wire g6789;
  wire g679;
  wire g6790;
  wire g6791;
  wire g6792;
  wire g6793;
  wire g6794;
  wire g6796;
  wire g6797;
  wire g680;
  wire g6800;
  wire g6801;
  wire g6803;
  wire g6806;
  wire g6809;
  wire g681;
  wire g6812;
  wire g6817;
  wire g6818;
  wire g6819;
  wire g682;
  wire g6820;
  wire g6824;
  wire g6825;
  wire g6826;
  wire g6827;
  wire g683;
  wire g6832;
  wire g6833;
  wire g6834;
  wire g6835;
  wire g6836;
  wire g6837;
  wire g6838;
  wire g6839;
  wire g684;
  wire g6840;
  wire g6841;
  wire g6842;
  wire g6844;
  wire g6845;
  wire g6849;
  wire g685;
  wire g6850;
  wire g6853;
  wire g6854;
  wire g687;
  wire g688;
  wire g689;
  wire g690;
  wire g691;
  wire g692;
  wire g693;
  wire g694;
  wire g695;
  wire g696;
  wire g697;
  wire g698;
  wire g699;
  wire g7;
  input g702;
  input g705;
  wire g719;
  wire g729;
  wire g736;
  wire g743;
  wire g749;
  wire g754;
  wire g760;
  wire g766;
  wire g774;
  wire g784;
  wire g791;
  wire g798;
  wire g804;
  wire g809;
  wire g815;
  wire g821;
  input g89;
  wire g894;
  wire g898;
  wire g899;
  wire g900;
  wire g908;
  wire g909;
  wire g917;
  wire g922;
  wire g927;
  input g94;
  wire g952;
  wire g965;
  input g98;
  wire g980;
  wire g996;
  al_inv _0419_ (
    .a(\DFF_197.Q ),
    .y(\DFF_80.D )
  );
  al_inv _0420_ (
    .a(\DFF_208.Q ),
    .y(\DFF_153.D )
  );
  al_nand2ft _0421_ (
    .a(\DFF_69.Q ),
    .b(\DFF_21.Q ),
    .y(_0000_)
  );
  al_aoi21ftf _0422_ (
    .a(\DFF_153.Q ),
    .b(\DFF_135.Q ),
    .c(_0000_),
    .y(g4809)
  );
  al_nand2ft _0423_ (
    .a(\DFF_37.Q ),
    .b(\DFF_146.Q ),
    .y(_0001_)
  );
  al_and2ft _0424_ (
    .a(\DFF_146.Q ),
    .b(\DFF_37.Q ),
    .y(_0002_)
  );
  al_nand2ft _0425_ (
    .a(_0002_),
    .b(_0001_),
    .y(_0003_)
  );
  al_and3 _0426_ (
    .a(\DFF_178.Q ),
    .b(\DFF_52.Q ),
    .c(\DFF_168.Q ),
    .y(_0004_)
  );
  al_or3fft _0427_ (
    .a(\DFF_3.Q ),
    .b(_0004_),
    .c(_0001_),
    .y(_0005_)
  );
  al_or3 _0428_ (
    .a(\DFF_164.Q ),
    .b(\DFF_87.Q ),
    .c(\DFF_70.Q ),
    .y(_0006_)
  );
  al_aoi21 _0429_ (
    .a(_0005_),
    .b(_0003_),
    .c(_0006_),
    .y(_0007_)
  );
  al_and2 _0430_ (
    .a(\DFF_3.Q ),
    .b(_0004_),
    .y(_0008_)
  );
  al_and3 _0431_ (
    .a(\DFF_37.Q ),
    .b(\DFF_146.Q ),
    .c(_0008_),
    .y(_0009_)
  );
  al_nand2ft _0432_ (
    .a(\DFF_87.Q ),
    .b(\DFF_164.Q ),
    .y(_0010_)
  );
  al_mux2l _0433_ (
    .a(\DFF_188.Q ),
    .b(\DFF_200.Q ),
    .s(\DFF_178.Q ),
    .y(_0011_)
  );
  al_mux2l _0434_ (
    .a(\DFF_208.Q ),
    .b(\DFF_129.Q ),
    .s(\DFF_178.Q ),
    .y(_0012_)
  );
  al_mux2l _0435_ (
    .a(_0011_),
    .b(_0012_),
    .s(\DFF_168.Q ),
    .y(_0013_)
  );
  al_mux2l _0436_ (
    .a(\DFF_207.Q ),
    .b(\DFF_111.Q ),
    .s(\DFF_178.Q ),
    .y(_0014_)
  );
  al_mux2l _0437_ (
    .a(\DFF_26.Q ),
    .b(\DFF_51.Q ),
    .s(\DFF_178.Q ),
    .y(_0015_)
  );
  al_mux2l _0438_ (
    .a(_0014_),
    .b(_0015_),
    .s(\DFF_168.Q ),
    .y(_0016_)
  );
  al_mux2l _0439_ (
    .a(_0013_),
    .b(_0016_),
    .s(\DFF_52.Q ),
    .y(_0017_)
  );
  al_nand2 _0440_ (
    .a(\DFF_70.Q ),
    .b(_0017_),
    .y(_0018_)
  );
  al_inv _0441_ (
    .a(\DFF_70.Q ),
    .y(_0019_)
  );
  al_oa21ftf _0442_ (
    .a(_0019_),
    .b(_0017_),
    .c(_0003_),
    .y(_0020_)
  );
  al_nand3ftt _0443_ (
    .a(_0010_),
    .b(_0018_),
    .c(_0020_),
    .y(_0021_)
  );
  al_nand2 _0444_ (
    .a(\DFF_52.Q ),
    .b(_0013_),
    .y(_0022_)
  );
  al_nand2ft _0445_ (
    .a(\DFF_52.Q ),
    .b(_0016_),
    .y(_0023_)
  );
  al_nand3 _0446_ (
    .a(_0019_),
    .b(_0022_),
    .c(_0023_),
    .y(_0024_)
  );
  al_nand3ftt _0447_ (
    .a(_0003_),
    .b(_0024_),
    .c(_0018_),
    .y(_0025_)
  );
  al_ao21ftf _0448_ (
    .a(_0002_),
    .b(_0001_),
    .c(_0005_),
    .y(_0026_)
  );
  al_mux2h _0449_ (
    .a(_0005_),
    .b(_0026_),
    .s(_0019_),
    .y(_0027_)
  );
  al_and2 _0450_ (
    .a(\DFF_164.Q ),
    .b(\DFF_87.Q ),
    .y(_0028_)
  );
  al_ao21ttf _0451_ (
    .a(_0027_),
    .b(_0025_),
    .c(_0028_),
    .y(_0029_)
  );
  al_nand2ft _0452_ (
    .a(\DFF_164.Q ),
    .b(\DFF_87.Q ),
    .y(_0030_)
  );
  al_nand3 _0453_ (
    .a(_0021_),
    .b(_0030_),
    .c(_0029_),
    .y(_0031_)
  );
  al_nand2 _0454_ (
    .a(_0009_),
    .b(_0031_),
    .y(_0032_)
  );
  al_nand3ftt _0455_ (
    .a(_0007_),
    .b(\DFF_87.Q ),
    .c(_0032_),
    .y(_0033_)
  );
  al_inv _0456_ (
    .a(_0009_),
    .y(_0034_)
  );
  al_nand2 _0457_ (
    .a(_0021_),
    .b(_0029_),
    .y(_0035_)
  );
  al_and3ftt _0458_ (
    .a(_0010_),
    .b(_0009_),
    .c(_0025_),
    .y(_0036_)
  );
  al_aoi21 _0459_ (
    .a(_0034_),
    .b(_0035_),
    .c(_0036_),
    .y(_0037_)
  );
  al_aoi21 _0460_ (
    .a(\DFF_164.Q ),
    .b(_0027_),
    .c(_0028_),
    .y(_0038_)
  );
  al_ao21 _0461_ (
    .a(_0034_),
    .b(_0035_),
    .c(_0038_),
    .y(_0039_)
  );
  al_nand3ftt _0462_ (
    .a(_0007_),
    .b(_0032_),
    .c(_0039_),
    .y(_0040_)
  );
  al_ao21ttf _0463_ (
    .a(_0037_),
    .b(_0033_),
    .c(_0040_),
    .y(\DFF_161.D )
  );
  al_inv _0464_ (
    .a(g47),
    .y(\DFF_191.D )
  );
  al_and2ft _0465_ (
    .a(\DFF_209.Q ),
    .b(\DFF_117.Q ),
    .y(_0041_)
  );
  al_and2ft _0466_ (
    .a(\DFF_117.Q ),
    .b(\DFF_209.Q ),
    .y(_0042_)
  );
  al_or2 _0467_ (
    .a(_0041_),
    .b(_0042_),
    .y(_0043_)
  );
  al_or2 _0468_ (
    .a(\DFF_123.Q ),
    .b(\DFF_128.Q ),
    .y(_0044_)
  );
  al_nand2 _0469_ (
    .a(\DFF_123.Q ),
    .b(\DFF_128.Q ),
    .y(_0045_)
  );
  al_ao21 _0470_ (
    .a(_0044_),
    .b(_0045_),
    .c(_0043_),
    .y(_0046_)
  );
  al_nand3 _0471_ (
    .a(_0044_),
    .b(_0045_),
    .c(_0043_),
    .y(_0047_)
  );
  al_nand2ft _0472_ (
    .a(\DFF_98.Q ),
    .b(\DFF_127.Q ),
    .y(_0048_)
  );
  al_nand2ft _0473_ (
    .a(\DFF_127.Q ),
    .b(\DFF_98.Q ),
    .y(_0049_)
  );
  al_and3 _0474_ (
    .a(\DFF_10.Q ),
    .b(_0048_),
    .c(_0049_),
    .y(_0050_)
  );
  al_ao21 _0475_ (
    .a(_0048_),
    .b(_0049_),
    .c(\DFF_10.Q ),
    .y(_0051_)
  );
  al_and2ft _0476_ (
    .a(_0050_),
    .b(_0051_),
    .y(_0052_)
  );
  al_nand3 _0477_ (
    .a(_0047_),
    .b(_0046_),
    .c(_0052_),
    .y(_0053_)
  );
  al_ao21 _0478_ (
    .a(_0047_),
    .b(_0046_),
    .c(_0052_),
    .y(_0054_)
  );
  al_nor2 _0479_ (
    .a(\DFF_23.Q ),
    .b(\DFF_6.Q ),
    .y(_0055_)
  );
  al_nand2 _0480_ (
    .a(\DFF_23.Q ),
    .b(\DFF_6.Q ),
    .y(_0056_)
  );
  al_and2ft _0481_ (
    .a(_0055_),
    .b(_0056_),
    .y(_0057_)
  );
  al_nand3 _0482_ (
    .a(_0057_),
    .b(_0054_),
    .c(_0053_),
    .y(_0058_)
  );
  al_ao21 _0483_ (
    .a(_0054_),
    .b(_0053_),
    .c(_0057_),
    .y(_0059_)
  );
  al_and2ft _0484_ (
    .a(g37),
    .b(g38),
    .y(_0060_)
  );
  al_nand2ft _0485_ (
    .a(g38),
    .b(g37),
    .y(_0061_)
  );
  al_nand2ft _0486_ (
    .a(_0060_),
    .b(_0061_),
    .y(_0062_)
  );
  al_nand2ft _0487_ (
    .a(g39),
    .b(g40),
    .y(_0063_)
  );
  al_nand2ft _0488_ (
    .a(g40),
    .b(g39),
    .y(_0064_)
  );
  al_ao21 _0489_ (
    .a(_0063_),
    .b(_0064_),
    .c(_0062_),
    .y(_0065_)
  );
  al_and3 _0490_ (
    .a(_0063_),
    .b(_0064_),
    .c(_0062_),
    .y(_0066_)
  );
  al_and2ft _0491_ (
    .a(g32),
    .b(g36),
    .y(_0067_)
  );
  al_nand2ft _0492_ (
    .a(g36),
    .b(g32),
    .y(_0068_)
  );
  al_nand2ft _0493_ (
    .a(_0067_),
    .b(_0068_),
    .y(_0069_)
  );
  al_oai21ftf _0494_ (
    .a(_0065_),
    .b(_0066_),
    .c(_0069_),
    .y(_0070_)
  );
  al_nor3fft _0495_ (
    .a(_0069_),
    .b(_0065_),
    .c(_0066_),
    .y(_0071_)
  );
  al_and2ft _0496_ (
    .a(_0071_),
    .b(_0070_),
    .y(_0072_)
  );
  al_or3fft _0497_ (
    .a(_0058_),
    .b(_0059_),
    .c(_0072_),
    .y(_0073_)
  );
  al_aoi21ttf _0498_ (
    .a(_0058_),
    .b(_0059_),
    .c(_0072_),
    .y(_0074_)
  );
  al_nand2ft _0499_ (
    .a(_0074_),
    .b(_0073_),
    .y(\DFF_14.D )
  );
  al_inv _0500_ (
    .a(\DFF_188.Q ),
    .y(\DFF_69.D )
  );
  al_inv _0501_ (
    .a(\DFF_125.Q ),
    .y(_0075_)
  );
  al_nand2ft _0502_ (
    .a(\DFF_142.Q ),
    .b(\DFF_61.Q ),
    .y(_0076_)
  );
  al_and2ft _0503_ (
    .a(\DFF_61.Q ),
    .b(\DFF_142.Q ),
    .y(_0077_)
  );
  al_nand2ft _0504_ (
    .a(_0077_),
    .b(_0076_),
    .y(_0078_)
  );
  al_and3 _0505_ (
    .a(\DFF_43.Q ),
    .b(\DFF_201.Q ),
    .c(\DFF_17.Q ),
    .y(_0079_)
  );
  al_or3fft _0506_ (
    .a(\DFF_134.Q ),
    .b(_0079_),
    .c(_0076_),
    .y(_0080_)
  );
  al_or3 _0507_ (
    .a(\DFF_125.Q ),
    .b(\DFF_50.Q ),
    .c(\DFF_148.Q ),
    .y(_0081_)
  );
  al_aoi21 _0508_ (
    .a(_0080_),
    .b(_0078_),
    .c(_0081_),
    .y(_0082_)
  );
  al_and3 _0509_ (
    .a(\DFF_142.Q ),
    .b(\DFF_134.Q ),
    .c(_0079_),
    .y(_0083_)
  );
  al_and2 _0510_ (
    .a(\DFF_61.Q ),
    .b(_0083_),
    .y(_0084_)
  );
  al_inv _0511_ (
    .a(_0078_),
    .y(_0085_)
  );
  al_inv _0512_ (
    .a(\DFF_148.Q ),
    .y(_0086_)
  );
  al_inv _0513_ (
    .a(\DFF_17.Q ),
    .y(_0087_)
  );
  al_mux2l _0514_ (
    .a(\DFF_207.Q ),
    .b(\DFF_26.Q ),
    .s(\DFF_43.Q ),
    .y(_0088_)
  );
  al_or2ft _0515_ (
    .a(\DFF_201.Q ),
    .b(_0088_),
    .y(_0089_)
  );
  al_mux2l _0516_ (
    .a(\DFF_111.Q ),
    .b(\DFF_51.Q ),
    .s(\DFF_43.Q ),
    .y(_0090_)
  );
  al_or2 _0517_ (
    .a(\DFF_201.Q ),
    .b(_0090_),
    .y(_0091_)
  );
  al_nand3 _0518_ (
    .a(_0087_),
    .b(_0091_),
    .c(_0089_),
    .y(_0092_)
  );
  al_mux2l _0519_ (
    .a(\DFF_188.Q ),
    .b(\DFF_208.Q ),
    .s(\DFF_43.Q ),
    .y(_0093_)
  );
  al_mux2l _0520_ (
    .a(\DFF_200.Q ),
    .b(\DFF_129.Q ),
    .s(\DFF_43.Q ),
    .y(_0094_)
  );
  al_mux2l _0521_ (
    .a(_0093_),
    .b(_0094_),
    .s(\DFF_201.Q ),
    .y(_0095_)
  );
  al_nand2 _0522_ (
    .a(\DFF_17.Q ),
    .b(_0095_),
    .y(_0096_)
  );
  al_nand3 _0523_ (
    .a(_0086_),
    .b(_0092_),
    .c(_0096_),
    .y(_0097_)
  );
  al_or2 _0524_ (
    .a(_0087_),
    .b(_0095_),
    .y(_0098_)
  );
  al_ao21 _0525_ (
    .a(_0091_),
    .b(_0089_),
    .c(\DFF_17.Q ),
    .y(_0099_)
  );
  al_nand3 _0526_ (
    .a(\DFF_148.Q ),
    .b(_0098_),
    .c(_0099_),
    .y(_0100_)
  );
  al_nand3 _0527_ (
    .a(_0085_),
    .b(_0097_),
    .c(_0100_),
    .y(_0101_)
  );
  al_or3fft _0528_ (
    .a(_0075_),
    .b(\DFF_50.Q ),
    .c(_0101_),
    .y(_0102_)
  );
  al_nand3 _0529_ (
    .a(\DFF_148.Q ),
    .b(_0092_),
    .c(_0096_),
    .y(_0103_)
  );
  al_nand3 _0530_ (
    .a(_0086_),
    .b(_0098_),
    .c(_0099_),
    .y(_0104_)
  );
  al_nand3 _0531_ (
    .a(_0085_),
    .b(_0103_),
    .c(_0104_),
    .y(_0105_)
  );
  al_nand3 _0532_ (
    .a(_0086_),
    .b(_0080_),
    .c(_0078_),
    .y(_0106_)
  );
  al_ao21 _0533_ (
    .a(_0080_),
    .b(_0078_),
    .c(_0086_),
    .y(_0107_)
  );
  al_nand3 _0534_ (
    .a(_0078_),
    .b(_0106_),
    .c(_0107_),
    .y(_0108_)
  );
  al_and2 _0535_ (
    .a(\DFF_125.Q ),
    .b(\DFF_50.Q ),
    .y(_0109_)
  );
  al_nand3 _0536_ (
    .a(_0108_),
    .b(_0109_),
    .c(_0105_),
    .y(_0110_)
  );
  al_nand2ft _0537_ (
    .a(\DFF_50.Q ),
    .b(\DFF_125.Q ),
    .y(_0111_)
  );
  al_nand3 _0538_ (
    .a(_0111_),
    .b(_0110_),
    .c(_0102_),
    .y(_0112_)
  );
  al_nand2 _0539_ (
    .a(_0084_),
    .b(_0112_),
    .y(_0113_)
  );
  al_nand3fft _0540_ (
    .a(_0075_),
    .b(_0082_),
    .c(_0113_),
    .y(_0114_)
  );
  al_ao21 _0541_ (
    .a(_0110_),
    .b(_0102_),
    .c(_0084_),
    .y(_0115_)
  );
  al_and2ft _0542_ (
    .a(\DFF_125.Q ),
    .b(\DFF_50.Q ),
    .y(_0116_)
  );
  al_nand3 _0543_ (
    .a(_0084_),
    .b(_0116_),
    .c(_0101_),
    .y(_0117_)
  );
  al_and2 _0544_ (
    .a(_0117_),
    .b(_0115_),
    .y(_0118_)
  );
  al_oa21ftt _0545_ (
    .a(_0076_),
    .b(_0077_),
    .c(_0075_),
    .y(_0119_)
  );
  al_ao21ttf _0546_ (
    .a(_0106_),
    .b(_0107_),
    .c(_0119_),
    .y(_0120_)
  );
  al_nand3 _0547_ (
    .a(\DFF_50.Q ),
    .b(_0120_),
    .c(_0115_),
    .y(_0121_)
  );
  al_nand3ftt _0548_ (
    .a(_0082_),
    .b(_0113_),
    .c(_0121_),
    .y(_0122_)
  );
  al_ao21ttf _0549_ (
    .a(_0118_),
    .b(_0114_),
    .c(_0122_),
    .y(\DFF_190.D )
  );
  al_inv _0550_ (
    .a(g41),
    .y(_0123_)
  );
  al_inv _0551_ (
    .a(g22),
    .y(_0124_)
  );
  al_nand3 _0552_ (
    .a(_0123_),
    .b(_0058_),
    .c(_0059_),
    .y(_0125_)
  );
  al_and2 _0553_ (
    .a(\DFF_14.Q ),
    .b(_0125_),
    .y(_0126_)
  );
  al_nand3 _0554_ (
    .a(\DFF_147.Q ),
    .b(_0124_),
    .c(_0126_),
    .y(g6282)
  );
  al_and2ft _0555_ (
    .a(\DFF_187.Q ),
    .b(\DFF_90.Q ),
    .y(_0127_)
  );
  al_nand2ft _0556_ (
    .a(\DFF_90.Q ),
    .b(\DFF_187.Q ),
    .y(_0128_)
  );
  al_and2ft _0557_ (
    .a(\DFF_79.Q ),
    .b(\DFF_167.Q ),
    .y(_0129_)
  );
  al_nand2ft _0558_ (
    .a(\DFF_167.Q ),
    .b(\DFF_79.Q ),
    .y(_0130_)
  );
  al_nand2ft _0559_ (
    .a(_0129_),
    .b(_0130_),
    .y(_0131_)
  );
  al_and3ftt _0560_ (
    .a(_0127_),
    .b(_0128_),
    .c(_0131_),
    .y(_0132_)
  );
  al_ao21ftt _0561_ (
    .a(_0127_),
    .b(_0128_),
    .c(_0131_),
    .y(_0133_)
  );
  al_nand2ft _0562_ (
    .a(_0132_),
    .b(_0133_),
    .y(_0134_)
  );
  al_and2ft _0563_ (
    .a(\DFF_27.Q ),
    .b(\DFF_186.Q ),
    .y(_0135_)
  );
  al_nand2ft _0564_ (
    .a(\DFF_186.Q ),
    .b(\DFF_27.Q ),
    .y(_0136_)
  );
  al_and2ft _0565_ (
    .a(\DFF_44.Q ),
    .b(\DFF_63.Q ),
    .y(_0137_)
  );
  al_nand2ft _0566_ (
    .a(\DFF_63.Q ),
    .b(\DFF_44.Q ),
    .y(_0138_)
  );
  al_nand2ft _0567_ (
    .a(_0137_),
    .b(_0138_),
    .y(_0139_)
  );
  al_and3ftt _0568_ (
    .a(_0135_),
    .b(_0136_),
    .c(_0139_),
    .y(_0140_)
  );
  al_ao21ftt _0569_ (
    .a(_0135_),
    .b(_0136_),
    .c(_0139_),
    .y(_0141_)
  );
  al_aoi21ftf _0570_ (
    .a(_0140_),
    .b(_0141_),
    .c(_0134_),
    .y(_0142_)
  );
  al_or3ftt _0571_ (
    .a(_0141_),
    .b(_0140_),
    .c(_0134_),
    .y(_0143_)
  );
  al_nand2ft _0572_ (
    .a(_0142_),
    .b(_0143_),
    .y(\DFF_23.D )
  );
  al_or3 _0573_ (
    .a(_0123_),
    .b(\DFF_23.D ),
    .c(g6282),
    .y(g6284)
  );
  al_and2ft _0574_ (
    .a(g102),
    .b(g89),
    .y(g2584)
  );
  al_aoi21 _0575_ (
    .a(_0009_),
    .b(_0031_),
    .c(_0007_),
    .y(_0144_)
  );
  al_ao21ttf _0576_ (
    .a(\DFF_87.Q ),
    .b(_0144_),
    .c(_0037_),
    .y(_0145_)
  );
  al_mux2h _0577_ (
    .a(\DFF_51.Q ),
    .b(_0145_),
    .s(\DFF_179.Q ),
    .y(\DFF_87.D )
  );
  al_nand3 _0578_ (
    .a(\DFF_37.Q ),
    .b(\DFF_3.Q ),
    .c(_0004_),
    .y(_0146_)
  );
  al_oa21ftt _0579_ (
    .a(\DFF_146.Q ),
    .b(_0146_),
    .c(_0006_),
    .y(_0147_)
  );
  al_ao21 _0580_ (
    .a(\DFF_178.Q ),
    .b(\DFF_168.Q ),
    .c(\DFF_52.Q ),
    .y(_0148_)
  );
  al_and3ftt _0581_ (
    .a(_0004_),
    .b(_0148_),
    .c(_0147_),
    .y(_0149_)
  );
  al_mux2h _0582_ (
    .a(\DFF_200.Q ),
    .b(_0149_),
    .s(\DFF_179.Q ),
    .y(\DFF_52.D )
  );
  al_and3 _0583_ (
    .a(\DFF_140.Q ),
    .b(\DFF_126.Q ),
    .c(\DFF_144.Q ),
    .y(_0150_)
  );
  al_and3 _0584_ (
    .a(\DFF_154.Q ),
    .b(\DFF_36.Q ),
    .c(_0150_),
    .y(_0151_)
  );
  al_and3 _0585_ (
    .a(\DFF_15.Q ),
    .b(\DFF_40.Q ),
    .c(_0151_),
    .y(_0152_)
  );
  al_and3 _0586_ (
    .a(\DFF_64.Q ),
    .b(\DFF_121.Q ),
    .c(_0152_),
    .y(_0153_)
  );
  al_nand2 _0587_ (
    .a(\DFF_158.Q ),
    .b(_0153_),
    .y(_0154_)
  );
  al_inv _0588_ (
    .a(g639),
    .y(_0155_)
  );
  al_and2 _0589_ (
    .a(\DFF_158.Q ),
    .b(\DFF_189.Q ),
    .y(_0156_)
  );
  al_nand3 _0590_ (
    .a(\DFF_88.Q ),
    .b(_0156_),
    .c(_0153_),
    .y(_0157_)
  );
  al_or3fft _0591_ (
    .a(\DFF_24.Q ),
    .b(\DFF_83.Q ),
    .c(_0157_),
    .y(_0158_)
  );
  al_oa21ftf _0592_ (
    .a(\DFF_151.Q ),
    .b(_0158_),
    .c(_0155_),
    .y(_0159_)
  );
  al_or2 _0593_ (
    .a(\DFF_158.Q ),
    .b(_0153_),
    .y(_0160_)
  );
  al_and3 _0594_ (
    .a(_0154_),
    .b(_0160_),
    .c(_0159_),
    .y(\DFF_158.D )
  );
  al_or3 _0595_ (
    .a(_0123_),
    .b(\DFF_63.Q ),
    .c(g6282),
    .y(g6372)
  );
  al_and2ft _0596_ (
    .a(\DFF_82.Q ),
    .b(\DFF_129.Q ),
    .y(_0161_)
  );
  al_nand2 _0597_ (
    .a(\DFF_134.Q ),
    .b(_0079_),
    .y(_0162_)
  );
  al_nor2 _0598_ (
    .a(\DFF_134.Q ),
    .b(_0079_),
    .y(_0163_)
  );
  al_nand3ftt _0599_ (
    .a(_0081_),
    .b(_0080_),
    .c(_0078_),
    .y(_0164_)
  );
  al_aoi21ttf _0600_ (
    .a(\DFF_61.Q ),
    .b(_0083_),
    .c(_0164_),
    .y(_0165_)
  );
  al_ao21ftf _0601_ (
    .a(_0163_),
    .b(_0162_),
    .c(_0165_),
    .y(_0166_)
  );
  al_inv _0602_ (
    .a(\DFF_82.Q ),
    .y(_0167_)
  );
  al_nor2 _0603_ (
    .a(_0167_),
    .b(_0082_),
    .y(_0168_)
  );
  al_ao21 _0604_ (
    .a(_0168_),
    .b(_0166_),
    .c(_0161_),
    .y(\DFF_134.D )
  );
  al_mux2h _0605_ (
    .a(\DFF_111.Q ),
    .b(_0040_),
    .s(\DFF_179.Q ),
    .y(\DFF_164.D )
  );
  al_mux2h _0606_ (
    .a(\DFF_111.Q ),
    .b(_0122_),
    .s(\DFF_82.Q ),
    .y(\DFF_50.D )
  );
  al_or3 _0607_ (
    .a(_0123_),
    .b(\DFF_90.Q ),
    .c(g6282),
    .y(g6362)
  );
  al_nand2 _0608_ (
    .a(\DFF_43.Q ),
    .b(\DFF_201.Q ),
    .y(_0169_)
  );
  al_aoi21ttf _0609_ (
    .a(\DFF_61.Q ),
    .b(_0083_),
    .c(_0081_),
    .y(_0170_)
  );
  al_or2 _0610_ (
    .a(\DFF_43.Q ),
    .b(\DFF_201.Q ),
    .y(_0171_)
  );
  al_and3 _0611_ (
    .a(_0169_),
    .b(_0171_),
    .c(_0170_),
    .y(_0172_)
  );
  al_mux2h _0612_ (
    .a(\DFF_208.Q ),
    .b(_0172_),
    .s(\DFF_82.Q ),
    .y(\DFF_201.D )
  );
  al_oa21 _0613_ (
    .a(g567),
    .b(\DFF_19.Q ),
    .c(\DFF_139.Q ),
    .y(_0173_)
  );
  al_aoi21ttf _0614_ (
    .a(g567),
    .b(\DFF_19.Q ),
    .c(_0173_),
    .y(\DFF_19.D )
  );
  al_aoi21 _0615_ (
    .a(\DFF_3.Q ),
    .b(_0004_),
    .c(\DFF_37.Q ),
    .y(_0174_)
  );
  al_ao21ftf _0616_ (
    .a(_0174_),
    .b(_0146_),
    .c(_0147_),
    .y(_0175_)
  );
  al_mux2h _0617_ (
    .a(\DFF_207.Q ),
    .b(_0175_),
    .s(\DFF_179.Q ),
    .y(\DFF_37.D )
  );
  al_or3ftt _0618_ (
    .a(_0146_),
    .b(\DFF_146.Q ),
    .c(_0007_),
    .y(_0176_)
  );
  al_oa21ttf _0619_ (
    .a(_0006_),
    .b(_0026_),
    .c(_0009_),
    .y(_0177_)
  );
  al_nand3 _0620_ (
    .a(\DFF_179.Q ),
    .b(_0177_),
    .c(_0176_),
    .y(_0178_)
  );
  al_ao21ftf _0621_ (
    .a(\DFF_179.Q ),
    .b(\DFF_26.Q ),
    .c(_0178_),
    .y(\DFF_146.D )
  );
  al_or3 _0622_ (
    .a(_0123_),
    .b(\DFF_44.Q ),
    .c(g6282),
    .y(g6364)
  );
  al_and3 _0623_ (
    .a(g567),
    .b(\DFF_19.Q ),
    .c(\DFF_58.Q ),
    .y(_0179_)
  );
  al_ao21 _0624_ (
    .a(g567),
    .b(\DFF_19.Q ),
    .c(\DFF_58.Q ),
    .y(_0180_)
  );
  al_nor3fft _0625_ (
    .a(\DFF_139.Q ),
    .b(_0180_),
    .c(_0179_),
    .y(\DFF_58.D )
  );
  al_nand2 _0626_ (
    .a(\DFF_178.Q ),
    .b(\DFF_168.Q ),
    .y(_0181_)
  );
  al_or2 _0627_ (
    .a(\DFF_178.Q ),
    .b(\DFF_168.Q ),
    .y(_0182_)
  );
  al_and3 _0628_ (
    .a(_0181_),
    .b(_0182_),
    .c(_0147_),
    .y(_0183_)
  );
  al_mux2h _0629_ (
    .a(\DFF_208.Q ),
    .b(_0183_),
    .s(\DFF_179.Q ),
    .y(\DFF_178.D )
  );
  al_or3 _0630_ (
    .a(_0123_),
    .b(\DFF_27.Q ),
    .c(g6282),
    .y(g6370)
  );
  al_aoi21ttf _0631_ (
    .a(\DFF_140.Q ),
    .b(\DFF_144.Q ),
    .c(g639),
    .y(_0184_)
  );
  al_oa21 _0632_ (
    .a(\DFF_140.Q ),
    .b(\DFF_144.Q ),
    .c(_0184_),
    .y(\DFF_144.D )
  );
  al_and2ft _0633_ (
    .a(\DFF_197.Q ),
    .b(g45),
    .y(\DFF_197.D )
  );
  al_or3 _0634_ (
    .a(_0123_),
    .b(\DFF_167.Q ),
    .c(g6282),
    .y(g6360)
  );
  al_aoi21ftf _0635_ (
    .a(\DFF_151.Q ),
    .b(_0158_),
    .c(_0159_),
    .y(\DFF_151.D )
  );
  al_aoi21 _0636_ (
    .a(\DFF_15.Q ),
    .b(_0151_),
    .c(_0155_),
    .y(_0185_)
  );
  al_oa21 _0637_ (
    .a(\DFF_15.Q ),
    .b(_0151_),
    .c(_0185_),
    .y(\DFF_15.D )
  );
  al_and3 _0638_ (
    .a(\DFF_28.Q ),
    .b(\DFF_141.Q ),
    .c(_0179_),
    .y(_0186_)
  );
  al_and2 _0639_ (
    .a(\DFF_30.Q ),
    .b(_0186_),
    .y(_0187_)
  );
  al_or2 _0640_ (
    .a(\DFF_30.Q ),
    .b(_0186_),
    .y(_0188_)
  );
  al_nor3fft _0641_ (
    .a(\DFF_139.Q ),
    .b(_0188_),
    .c(_0187_),
    .y(\DFF_30.D )
  );
  al_and3fft _0642_ (
    .a(\DFF_168.Q ),
    .b(_0009_),
    .c(_0006_),
    .y(_0189_)
  );
  al_mux2h _0643_ (
    .a(\DFF_188.Q ),
    .b(_0189_),
    .s(\DFF_179.Q ),
    .y(\DFF_168.D )
  );
  al_aoi21 _0644_ (
    .a(_0084_),
    .b(_0112_),
    .c(_0082_),
    .y(_0190_)
  );
  al_ao21ttf _0645_ (
    .a(\DFF_125.Q ),
    .b(_0190_),
    .c(_0118_),
    .y(_0191_)
  );
  al_mux2h _0646_ (
    .a(\DFF_51.Q ),
    .b(_0191_),
    .s(\DFF_82.Q ),
    .y(\DFF_125.D )
  );
  al_aoi21 _0647_ (
    .a(\DFF_154.Q ),
    .b(_0150_),
    .c(\DFF_36.Q ),
    .y(_0192_)
  );
  al_nor3ftt _0648_ (
    .a(g639),
    .b(_0151_),
    .c(_0192_),
    .y(\DFF_36.D )
  );
  al_ao21 _0649_ (
    .a(\DFF_134.Q ),
    .b(_0079_),
    .c(\DFF_142.Q ),
    .y(_0193_)
  );
  al_ao21ftf _0650_ (
    .a(_0083_),
    .b(_0193_),
    .c(_0170_),
    .y(_0194_)
  );
  al_mux2h _0651_ (
    .a(\DFF_207.Q ),
    .b(_0194_),
    .s(\DFF_82.Q ),
    .y(\DFF_142.D )
  );
  al_or3 _0652_ (
    .a(\DFF_61.Q ),
    .b(_0083_),
    .c(_0082_),
    .y(_0195_)
  );
  al_nand3 _0653_ (
    .a(\DFF_82.Q ),
    .b(_0165_),
    .c(_0195_),
    .y(_0196_)
  );
  al_ao21ftf _0654_ (
    .a(\DFF_82.Q ),
    .b(\DFF_26.Q ),
    .c(_0196_),
    .y(\DFF_61.D )
  );
  al_aoi21 _0655_ (
    .a(\DFF_141.Q ),
    .b(_0179_),
    .c(\DFF_28.Q ),
    .y(_0197_)
  );
  al_nor3ftt _0656_ (
    .a(\DFF_139.Q ),
    .b(_0186_),
    .c(_0197_),
    .y(\DFF_28.D )
  );
  al_aoi21ttf _0657_ (
    .a(\DFF_141.Q ),
    .b(_0179_),
    .c(\DFF_139.Q ),
    .y(_0198_)
  );
  al_oa21 _0658_ (
    .a(\DFF_141.Q ),
    .b(_0179_),
    .c(_0198_),
    .y(\DFF_141.D )
  );
  al_and2ft _0659_ (
    .a(\DFF_179.Q ),
    .b(\DFF_129.Q ),
    .y(_0199_)
  );
  al_or2 _0660_ (
    .a(\DFF_3.Q ),
    .b(_0004_),
    .y(_0200_)
  );
  al_ao21ftf _0661_ (
    .a(_0008_),
    .b(_0200_),
    .c(_0177_),
    .y(_0201_)
  );
  al_aoi21ftf _0662_ (
    .a(_0006_),
    .b(_0026_),
    .c(\DFF_179.Q ),
    .y(_0202_)
  );
  al_ao21 _0663_ (
    .a(_0202_),
    .b(_0201_),
    .c(_0199_),
    .y(\DFF_3.D )
  );
  al_and2ft _0664_ (
    .a(\DFF_169.Q ),
    .b(g45),
    .y(\DFF_169.D )
  );
  al_and2ft _0665_ (
    .a(\DFF_140.Q ),
    .b(g639),
    .y(\DFF_140.D )
  );
  al_ao21 _0666_ (
    .a(\DFF_43.Q ),
    .b(\DFF_201.Q ),
    .c(\DFF_17.Q ),
    .y(_0203_)
  );
  al_and3ftt _0667_ (
    .a(_0079_),
    .b(_0203_),
    .c(_0170_),
    .y(_0204_)
  );
  al_mux2h _0668_ (
    .a(\DFF_200.Q ),
    .b(_0204_),
    .s(\DFF_82.Q ),
    .y(\DFF_17.D )
  );
  al_and3 _0669_ (
    .a(\DFF_170.Q ),
    .b(\DFF_30.Q ),
    .c(_0186_),
    .y(_0205_)
  );
  al_aoi21 _0670_ (
    .a(\DFF_30.Q ),
    .b(_0186_),
    .c(\DFF_170.Q ),
    .y(_0206_)
  );
  al_nor3ftt _0671_ (
    .a(\DFF_139.Q ),
    .b(_0205_),
    .c(_0206_),
    .y(\DFF_170.D )
  );
  al_aoi21 _0672_ (
    .a(\DFF_154.Q ),
    .b(_0150_),
    .c(_0155_),
    .y(_0207_)
  );
  al_oa21 _0673_ (
    .a(\DFF_154.Q ),
    .b(_0150_),
    .c(_0207_),
    .y(\DFF_154.D )
  );
  al_or3 _0674_ (
    .a(_0123_),
    .b(\DFF_79.Q ),
    .c(g6282),
    .y(g6366)
  );
  al_or3 _0675_ (
    .a(_0123_),
    .b(\DFF_187.Q ),
    .c(g6282),
    .y(g6374)
  );
  al_ao21 _0676_ (
    .a(\DFF_93.Q ),
    .b(_0205_),
    .c(\DFF_89.Q ),
    .y(_0208_)
  );
  al_nand3 _0677_ (
    .a(\DFF_93.Q ),
    .b(\DFF_89.Q ),
    .c(_0205_),
    .y(_0209_)
  );
  al_and3 _0678_ (
    .a(\DFF_139.Q ),
    .b(_0209_),
    .c(_0208_),
    .y(\DFF_89.D )
  );
  al_or3 _0679_ (
    .a(_0123_),
    .b(\DFF_186.Q ),
    .c(g6282),
    .y(g6368)
  );
  al_ao21 _0680_ (
    .a(_0156_),
    .b(_0153_),
    .c(\DFF_88.Q ),
    .y(_0210_)
  );
  al_and3 _0681_ (
    .a(_0157_),
    .b(_0210_),
    .c(_0159_),
    .y(\DFF_88.D )
  );
  al_nand3fft _0682_ (
    .a(_0167_),
    .b(\DFF_43.Q ),
    .c(_0170_),
    .y(_0211_)
  );
  al_ao21ftf _0683_ (
    .a(\DFF_69.D ),
    .b(_0167_),
    .c(_0211_),
    .y(\DFF_43.D )
  );
  al_aoi21 _0684_ (
    .a(\DFF_121.Q ),
    .b(_0152_),
    .c(_0155_),
    .y(_0212_)
  );
  al_oa21 _0685_ (
    .a(\DFF_121.Q ),
    .b(_0152_),
    .c(_0212_),
    .y(\DFF_121.D )
  );
  al_aoi21 _0686_ (
    .a(\DFF_15.Q ),
    .b(_0151_),
    .c(\DFF_40.Q ),
    .y(_0213_)
  );
  al_nor3ftt _0687_ (
    .a(g639),
    .b(_0152_),
    .c(_0213_),
    .y(\DFF_40.D )
  );
  al_ao21 _0688_ (
    .a(\DFF_158.Q ),
    .b(_0153_),
    .c(\DFF_189.Q ),
    .y(_0214_)
  );
  al_aoi21ttf _0689_ (
    .a(_0153_),
    .b(_0156_),
    .c(_0214_),
    .y(_0215_)
  );
  al_and2 _0690_ (
    .a(_0215_),
    .b(_0159_),
    .y(\DFF_189.D )
  );
  al_aoi21ttf _0691_ (
    .a(\DFF_93.Q ),
    .b(_0205_),
    .c(\DFF_139.Q ),
    .y(_0216_)
  );
  al_oa21 _0692_ (
    .a(\DFF_93.Q ),
    .b(_0205_),
    .c(_0216_),
    .y(\DFF_93.D )
  );
  al_aoi21 _0693_ (
    .a(\DFF_121.Q ),
    .b(_0152_),
    .c(\DFF_64.Q ),
    .y(_0217_)
  );
  al_nor3ftt _0694_ (
    .a(g639),
    .b(_0153_),
    .c(_0217_),
    .y(\DFF_64.D )
  );
  al_nand2ft _0695_ (
    .a(\DFF_114.Q ),
    .b(\DFF_55.Q ),
    .y(_0218_)
  );
  al_nand2ft _0696_ (
    .a(\DFF_55.Q ),
    .b(\DFF_114.Q ),
    .y(_0219_)
  );
  al_nand2ft _0697_ (
    .a(\DFF_176.Q ),
    .b(\DFF_109.Q ),
    .y(_0220_)
  );
  al_and2ft _0698_ (
    .a(\DFF_109.Q ),
    .b(\DFF_176.Q ),
    .y(_0221_)
  );
  al_and2ft _0699_ (
    .a(_0221_),
    .b(_0220_),
    .y(_0222_)
  );
  al_nand2ft _0700_ (
    .a(\DFF_157.Q ),
    .b(\DFF_60.Q ),
    .y(_0223_)
  );
  al_nand2ft _0701_ (
    .a(\DFF_60.Q ),
    .b(\DFF_157.Q ),
    .y(_0224_)
  );
  al_and3 _0702_ (
    .a(_0223_),
    .b(_0224_),
    .c(_0222_),
    .y(_0225_)
  );
  al_nand3 _0703_ (
    .a(_0218_),
    .b(_0219_),
    .c(_0225_),
    .y(_0226_)
  );
  al_nand2ft _0704_ (
    .a(\DFF_102.Q ),
    .b(\DFF_156.Q ),
    .y(_0227_)
  );
  al_aoi21ftf _0705_ (
    .a(\DFF_204.Q ),
    .b(\DFF_166.Q ),
    .c(_0227_),
    .y(_0228_)
  );
  al_nand2ft _0706_ (
    .a(\DFF_76.Q ),
    .b(\DFF_177.Q ),
    .y(_0229_)
  );
  al_nand2ft _0707_ (
    .a(\DFF_182.Q ),
    .b(\DFF_116.Q ),
    .y(_0230_)
  );
  al_and3 _0708_ (
    .a(_0229_),
    .b(_0230_),
    .c(_0228_),
    .y(_0231_)
  );
  al_nand2ft _0709_ (
    .a(\DFF_177.Q ),
    .b(\DFF_76.Q ),
    .y(_0232_)
  );
  al_ao21ftf _0710_ (
    .a(\DFF_116.Q ),
    .b(\DFF_182.Q ),
    .c(_0232_),
    .y(_0233_)
  );
  al_nand2ft _0711_ (
    .a(\DFF_156.Q ),
    .b(\DFF_102.Q ),
    .y(_0234_)
  );
  al_ao21ftf _0712_ (
    .a(\DFF_166.Q ),
    .b(\DFF_204.Q ),
    .c(_0234_),
    .y(_0235_)
  );
  al_nor2 _0713_ (
    .a(\DFF_172.Q ),
    .b(\DFF_152.Q ),
    .y(_0236_)
  );
  al_nand2 _0714_ (
    .a(\DFF_172.Q ),
    .b(\DFF_152.Q ),
    .y(_0237_)
  );
  al_nand2ft _0715_ (
    .a(_0236_),
    .b(_0237_),
    .y(_0238_)
  );
  al_nand2ft _0716_ (
    .a(\DFF_183.Q ),
    .b(\DFF_205.Q ),
    .y(_0239_)
  );
  al_nand2ft _0717_ (
    .a(\DFF_205.Q ),
    .b(\DFF_183.Q ),
    .y(_0240_)
  );
  al_and3 _0718_ (
    .a(_0239_),
    .b(_0240_),
    .c(_0238_),
    .y(_0241_)
  );
  al_nand3fft _0719_ (
    .a(_0233_),
    .b(_0235_),
    .c(_0241_),
    .y(_0242_)
  );
  al_nor3ftt _0720_ (
    .a(_0231_),
    .b(_0242_),
    .c(_0226_),
    .y(_0243_)
  );
  al_nand3fft _0721_ (
    .a(\DFF_110.Q ),
    .b(\DFF_105.Q ),
    .c(_0243_),
    .y(_0244_)
  );
  al_mux2l _0722_ (
    .a(\DFF_5.Q ),
    .b(\DFF_78.Q ),
    .s(_0244_),
    .y(\DFF_5.D )
  );
  al_mux2h _0723_ (
    .a(\DFF_173.Q ),
    .b(_0145_),
    .s(_0243_),
    .y(\DFF_173.D )
  );
  al_and2 _0724_ (
    .a(g702),
    .b(\DFF_191.Q ),
    .y(_0245_)
  );
  al_and3 _0725_ (
    .a(_0123_),
    .b(_0245_),
    .c(_0126_),
    .y(_0246_)
  );
  al_inv _0726_ (
    .a(\DFF_51.Q ),
    .y(_0247_)
  );
  al_and3ftt _0727_ (
    .a(\DFF_124.Q ),
    .b(\DFF_9.Q ),
    .c(\DFF_92.Q ),
    .y(_0248_)
  );
  al_and2 _0728_ (
    .a(\DFF_47.Q ),
    .b(_0248_),
    .y(_0249_)
  );
  al_nand3fft _0729_ (
    .a(\DFF_111.Q ),
    .b(_0247_),
    .c(_0249_),
    .y(_0250_)
  );
  al_nand2ft _0730_ (
    .a(_0250_),
    .b(_0246_),
    .y(_0251_)
  );
  al_mux2l _0731_ (
    .a(\DFF_75.Q ),
    .b(\DFF_129.Q ),
    .s(_0251_),
    .y(\DFF_75.D )
  );
  al_and3ftt _0732_ (
    .a(\DFF_169.Q ),
    .b(g41),
    .c(_0245_),
    .y(_0252_)
  );
  al_and2 _0733_ (
    .a(\DFF_80.Q ),
    .b(_0252_),
    .y(_0253_)
  );
  al_and3 _0734_ (
    .a(\DFF_14.Q ),
    .b(_0253_),
    .c(_0125_),
    .y(_0254_)
  );
  al_nor2 _0735_ (
    .a(\DFF_9.Q ),
    .b(\DFF_92.Q ),
    .y(_0255_)
  );
  al_and2ft _0736_ (
    .a(\DFF_124.Q ),
    .b(_0255_),
    .y(_0256_)
  );
  al_and2 _0737_ (
    .a(_0256_),
    .b(_0254_),
    .y(_0257_)
  );
  al_nand2ft _0738_ (
    .a(\DFF_92.Q ),
    .b(\DFF_9.Q ),
    .y(_0258_)
  );
  al_ao21ftf _0739_ (
    .a(\DFF_47.Q ),
    .b(_0248_),
    .c(_0258_),
    .y(_0259_)
  );
  al_and2 _0740_ (
    .a(_0259_),
    .b(_0254_),
    .y(_0260_)
  );
  al_inv _0741_ (
    .a(\DFF_200.Q ),
    .y(_0261_)
  );
  al_ao21ftf _0742_ (
    .a(\DFF_80.Q ),
    .b(\DFF_80.D ),
    .c(_0252_),
    .y(_0262_)
  );
  al_nor2 _0743_ (
    .a(\DFF_208.Q ),
    .b(_0262_),
    .y(_0263_)
  );
  al_and3 _0744_ (
    .a(\DFF_9.Q ),
    .b(\DFF_92.Q ),
    .c(\DFF_124.Q ),
    .y(_0264_)
  );
  al_and2ft _0745_ (
    .a(\DFF_129.Q ),
    .b(_0264_),
    .y(_0265_)
  );
  al_and3 _0746_ (
    .a(_0261_),
    .b(_0265_),
    .c(_0263_),
    .y(_0266_)
  );
  al_nor2 _0747_ (
    .a(_0250_),
    .b(_0262_),
    .y(_0267_)
  );
  al_and3fft _0748_ (
    .a(\DFF_153.D ),
    .b(_0262_),
    .c(_0265_),
    .y(_0268_)
  );
  al_or3 _0749_ (
    .a(_0267_),
    .b(_0268_),
    .c(_0266_),
    .y(_0269_)
  );
  al_nand3ftt _0750_ (
    .a(\DFF_26.Q ),
    .b(\DFF_47.Q ),
    .c(_0248_),
    .y(_0270_)
  );
  al_and3fft _0751_ (
    .a(_0247_),
    .b(_0262_),
    .c(\DFF_111.Q ),
    .y(_0271_)
  );
  al_and3ftt _0752_ (
    .a(_0270_),
    .b(\DFF_207.Q ),
    .c(_0271_),
    .y(_0272_)
  );
  al_and3ftt _0753_ (
    .a(\DFF_207.Q ),
    .b(\DFF_111.Q ),
    .c(\DFF_51.Q ),
    .y(_0273_)
  );
  al_and3fft _0754_ (
    .a(_0270_),
    .b(_0262_),
    .c(_0273_),
    .y(_0274_)
  );
  al_and3ftt _0755_ (
    .a(\DFF_200.Q ),
    .b(\DFF_129.Q ),
    .c(_0264_),
    .y(_0275_)
  );
  al_or3fft _0756_ (
    .a(\DFF_153.D ),
    .b(_0275_),
    .c(_0262_),
    .y(_0276_)
  );
  al_and3 _0757_ (
    .a(\DFF_26.Q ),
    .b(_0249_),
    .c(_0271_),
    .y(_0277_)
  );
  al_and3fft _0758_ (
    .a(_0274_),
    .b(_0277_),
    .c(_0276_),
    .y(_0278_)
  );
  al_and3fft _0759_ (
    .a(_0272_),
    .b(_0269_),
    .c(_0278_),
    .y(_0279_)
  );
  al_nor3ftt _0760_ (
    .a(_0279_),
    .b(_0257_),
    .c(_0260_),
    .y(_0280_)
  );
  al_nand3 _0761_ (
    .a(\DFF_188.Q ),
    .b(\DFF_60.Q ),
    .c(_0274_),
    .y(_0281_)
  );
  al_nand3 _0762_ (
    .a(\DFF_200.Q ),
    .b(g559),
    .c(_0268_),
    .y(_0282_)
  );
  al_and3 _0763_ (
    .a(\DFF_69.D ),
    .b(\DFF_84.Q ),
    .c(_0277_),
    .y(_0283_)
  );
  al_and2 _0764_ (
    .a(\DFF_188.Q ),
    .b(_0277_),
    .y(_0284_)
  );
  al_aoi21 _0765_ (
    .a(\DFF_163.Q ),
    .b(_0284_),
    .c(_0283_),
    .y(_0285_)
  );
  al_and3 _0766_ (
    .a(_0281_),
    .b(_0282_),
    .c(_0285_),
    .y(_0286_)
  );
  al_ao21ttf _0767_ (
    .a(\DFF_26.Q ),
    .b(_0260_),
    .c(_0286_),
    .y(_0287_)
  );
  al_inv _0768_ (
    .a(\DFF_99.Q ),
    .y(_0288_)
  );
  al_nand3 _0769_ (
    .a(_0288_),
    .b(\DFF_146.D ),
    .c(_0257_),
    .y(_0289_)
  );
  al_nand3 _0770_ (
    .a(\DFF_99.Q ),
    .b(_0256_),
    .c(_0254_),
    .y(_0290_)
  );
  al_aoi21ftf _0771_ (
    .a(_0290_),
    .b(\DFF_61.D ),
    .c(_0289_),
    .y(_0291_)
  );
  al_nand3fft _0772_ (
    .a(_0280_),
    .b(_0287_),
    .c(_0291_),
    .y(\DFF_167.D )
  );
  al_and3ftt _0773_ (
    .a(\DFF_26.Q ),
    .b(_0273_),
    .c(_0249_),
    .y(_0292_)
  );
  al_nand3 _0774_ (
    .a(\DFF_188.Q ),
    .b(_0292_),
    .c(_0246_),
    .y(_0293_)
  );
  al_nand2ft _0775_ (
    .a(\DFF_55.Q ),
    .b(_0293_),
    .y(\DFF_55.D )
  );
  al_mux2l _0776_ (
    .a(\DFF_179.Q ),
    .b(\DFF_188.Q ),
    .s(_0251_),
    .y(\DFF_179.D )
  );
  al_mux2l _0777_ (
    .a(\DFF_53.Q ),
    .b(\DFF_81.Q ),
    .s(_0244_),
    .y(\DFF_53.D )
  );
  al_nand3 _0778_ (
    .a(\DFF_179.Q ),
    .b(_0037_),
    .c(_0033_),
    .y(_0294_)
  );
  al_or2 _0779_ (
    .a(\DFF_51.Q ),
    .b(\DFF_179.Q ),
    .y(_0295_)
  );
  al_and3 _0780_ (
    .a(_0288_),
    .b(_0256_),
    .c(_0254_),
    .y(_0296_)
  );
  al_nand3 _0781_ (
    .a(_0295_),
    .b(_0296_),
    .c(_0294_),
    .y(_0297_)
  );
  al_nand3 _0782_ (
    .a(\DFF_82.Q ),
    .b(_0118_),
    .c(_0114_),
    .y(_0298_)
  );
  al_or2 _0783_ (
    .a(\DFF_51.Q ),
    .b(\DFF_82.Q ),
    .y(_0299_)
  );
  al_and3 _0784_ (
    .a(\DFF_99.Q ),
    .b(_0256_),
    .c(_0254_),
    .y(_0300_)
  );
  al_nand3 _0785_ (
    .a(_0299_),
    .b(_0300_),
    .c(_0298_),
    .y(_0301_)
  );
  al_aoi21ttf _0786_ (
    .a(_0259_),
    .b(_0254_),
    .c(_0279_),
    .y(_0302_)
  );
  al_nand3 _0787_ (
    .a(\DFF_51.Q ),
    .b(_0259_),
    .c(_0254_),
    .y(_0303_)
  );
  al_nand3 _0788_ (
    .a(\DFF_188.Q ),
    .b(\DFF_55.Q ),
    .c(_0274_),
    .y(_0304_)
  );
  al_and2 _0789_ (
    .a(\DFF_200.Q ),
    .b(_0268_),
    .y(_0305_)
  );
  al_nand3 _0790_ (
    .a(\DFF_69.D ),
    .b(\DFF_196.Q ),
    .c(_0277_),
    .y(_0306_)
  );
  al_aoi21ttf _0791_ (
    .a(g557),
    .b(_0305_),
    .c(_0306_),
    .y(_0307_)
  );
  al_aoi21ttf _0792_ (
    .a(\DFF_78.Q ),
    .b(_0284_),
    .c(_0307_),
    .y(_0308_)
  );
  al_and3 _0793_ (
    .a(_0304_),
    .b(_0308_),
    .c(_0303_),
    .y(_0309_)
  );
  al_ao21ftf _0794_ (
    .a(_0257_),
    .b(_0302_),
    .c(_0309_),
    .y(_0310_)
  );
  al_nand3ftt _0795_ (
    .a(_0310_),
    .b(_0301_),
    .c(_0297_),
    .y(\DFF_79.D )
  );
  al_nand3ftt _0796_ (
    .a(\DFF_189.Q ),
    .b(\DFF_111.Q ),
    .c(\DFF_158.Q ),
    .y(_0311_)
  );
  al_mux2l _0797_ (
    .a(\DFF_26.Q ),
    .b(\DFF_51.Q ),
    .s(\DFF_189.Q ),
    .y(_0312_)
  );
  al_nand3 _0798_ (
    .a(\DFF_207.Q ),
    .b(\DFF_158.Q ),
    .c(\DFF_189.Q ),
    .y(_0313_)
  );
  al_aoi21ftf _0799_ (
    .a(\DFF_158.Q ),
    .b(_0312_),
    .c(_0313_),
    .y(_0314_)
  );
  al_ao21 _0800_ (
    .a(_0311_),
    .b(_0314_),
    .c(\DFF_88.Q ),
    .y(_0315_)
  );
  al_mux2l _0801_ (
    .a(\DFF_208.Q ),
    .b(\DFF_129.Q ),
    .s(\DFF_189.Q ),
    .y(_0316_)
  );
  al_and3ftt _0802_ (
    .a(\DFF_189.Q ),
    .b(\DFF_158.Q ),
    .c(\DFF_200.Q ),
    .y(_0317_)
  );
  al_aoi21 _0803_ (
    .a(\DFF_188.Q ),
    .b(_0156_),
    .c(_0317_),
    .y(_0318_)
  );
  al_ao21ftf _0804_ (
    .a(\DFF_158.Q ),
    .b(_0316_),
    .c(_0318_),
    .y(_0319_)
  );
  al_nand2ft _0805_ (
    .a(\DFF_24.Q ),
    .b(\DFF_151.Q ),
    .y(_0320_)
  );
  al_and2ft _0806_ (
    .a(\DFF_151.Q ),
    .b(\DFF_24.Q ),
    .y(_0321_)
  );
  al_nand2ft _0807_ (
    .a(_0321_),
    .b(_0320_),
    .y(_0322_)
  );
  al_aoi21 _0808_ (
    .a(\DFF_88.Q ),
    .b(_0319_),
    .c(_0322_),
    .y(_0323_)
  );
  al_and3 _0809_ (
    .a(\DFF_83.Q ),
    .b(\DFF_88.Q ),
    .c(_0156_),
    .y(_0324_)
  );
  al_and2ft _0810_ (
    .a(_0320_),
    .b(_0324_),
    .y(_0325_)
  );
  al_aoi21 _0811_ (
    .a(_0315_),
    .b(_0323_),
    .c(_0325_),
    .y(\DFF_48.D )
  );
  al_nand3 _0812_ (
    .a(\DFF_69.D ),
    .b(\DFF_81.Q ),
    .c(_0277_),
    .y(_0326_)
  );
  al_aoi21ttf _0813_ (
    .a(g562),
    .b(_0305_),
    .c(_0326_),
    .y(_0327_)
  );
  al_aoi21ttf _0814_ (
    .a(\DFF_77.Q ),
    .b(_0284_),
    .c(_0327_),
    .y(_0328_)
  );
  al_nand3 _0815_ (
    .a(\DFF_188.Q ),
    .b(\DFF_172.Q ),
    .c(_0274_),
    .y(_0329_)
  );
  al_inv _0816_ (
    .a(\DFF_110.Q ),
    .y(_0330_)
  );
  al_nand3fft _0817_ (
    .a(_0330_),
    .b(\DFF_188.Q ),
    .c(_0274_),
    .y(_0331_)
  );
  al_nand2 _0818_ (
    .a(\DFF_94.Q ),
    .b(_0267_),
    .y(_0332_)
  );
  al_nand2 _0819_ (
    .a(\DFF_25.Q ),
    .b(_0272_),
    .y(_0333_)
  );
  al_and3 _0820_ (
    .a(_0331_),
    .b(_0332_),
    .c(_0333_),
    .y(_0334_)
  );
  al_nand3 _0821_ (
    .a(_0329_),
    .b(_0334_),
    .c(_0328_),
    .y(_0335_)
  );
  al_ao21 _0822_ (
    .a(\DFF_200.Q ),
    .b(_0260_),
    .c(_0335_),
    .y(_0336_)
  );
  al_nand3 _0823_ (
    .a(_0288_),
    .b(\DFF_52.D ),
    .c(_0257_),
    .y(_0337_)
  );
  al_aoi21ftf _0824_ (
    .a(_0290_),
    .b(\DFF_17.D ),
    .c(_0337_),
    .y(_0338_)
  );
  al_nand3fft _0825_ (
    .a(_0280_),
    .b(_0336_),
    .c(_0338_),
    .y(\DFF_27.D )
  );
  al_nand3 _0826_ (
    .a(\DFF_69.D ),
    .b(_0292_),
    .c(_0246_),
    .y(_0339_)
  );
  al_inv _0827_ (
    .a(\DFF_11.Q ),
    .y(_0340_)
  );
  al_mux2l _0828_ (
    .a(_0005_),
    .b(_0080_),
    .s(_0340_),
    .y(_0341_)
  );
  al_aoi21ftf _0829_ (
    .a(_0341_),
    .b(_0243_),
    .c(\DFF_110.Q ),
    .y(_0342_)
  );
  al_mux2l _0830_ (
    .a(_0342_),
    .b(\DFF_200.Q ),
    .s(_0339_),
    .y(\DFF_110.D )
  );
  al_mux2l _0831_ (
    .a(\DFF_77.Q ),
    .b(\DFF_175.Q ),
    .s(_0244_),
    .y(\DFF_77.D )
  );
  al_mux2l _0832_ (
    .a(\DFF_196.Q ),
    .b(\DFF_42.Q ),
    .s(_0244_),
    .y(\DFF_196.D )
  );
  al_and2 _0833_ (
    .a(_0324_),
    .b(_0153_),
    .y(_0343_)
  );
  al_nand2ft _0834_ (
    .a(\DFF_83.Q ),
    .b(_0157_),
    .y(_0344_)
  );
  al_ao21ftf _0835_ (
    .a(_0343_),
    .b(_0344_),
    .c(_0159_),
    .y(\DFF_83.D )
  );
  al_nand3 _0836_ (
    .a(_0288_),
    .b(_0256_),
    .c(_0254_),
    .y(_0345_)
  );
  al_nand3 _0837_ (
    .a(\DFF_99.Q ),
    .b(\DFF_142.D ),
    .c(_0257_),
    .y(_0346_)
  );
  al_aoi21ftf _0838_ (
    .a(_0345_),
    .b(\DFF_37.D ),
    .c(_0346_),
    .y(_0347_)
  );
  al_and3 _0839_ (
    .a(\DFF_188.Q ),
    .b(\DFF_109.Q ),
    .c(_0274_),
    .y(_0348_)
  );
  al_and3 _0840_ (
    .a(\DFF_188.Q ),
    .b(\DFF_73.Q ),
    .c(_0277_),
    .y(_0349_)
  );
  al_nand3 _0841_ (
    .a(\DFF_69.D ),
    .b(\DFF_96.Q ),
    .c(_0277_),
    .y(_0350_)
  );
  al_aoi21ttf _0842_ (
    .a(g560),
    .b(_0305_),
    .c(_0350_),
    .y(_0351_)
  );
  al_nand3fft _0843_ (
    .a(_0348_),
    .b(_0349_),
    .c(_0351_),
    .y(_0352_)
  );
  al_aoi21 _0844_ (
    .a(\DFF_207.Q ),
    .b(_0260_),
    .c(_0352_),
    .y(_0353_)
  );
  al_nand3ftt _0845_ (
    .a(_0280_),
    .b(_0353_),
    .c(_0347_),
    .y(\DFF_187.D )
  );
  al_mux2h _0846_ (
    .a(\DFF_20.Q ),
    .b(_0191_),
    .s(_0243_),
    .y(\DFF_20.D )
  );
  al_mux2l _0847_ (
    .a(\DFF_96.Q ),
    .b(\DFF_53.Q ),
    .s(_0244_),
    .y(\DFF_96.D )
  );
  al_oai21ftf _0848_ (
    .a(_0124_),
    .b(_0125_),
    .c(\DFF_131.Q ),
    .y(\DFF_131.D )
  );
  al_and2 _0849_ (
    .a(\DFF_109.Q ),
    .b(_0293_),
    .y(\DFF_109.D )
  );
  al_mux2l _0850_ (
    .a(\DFF_84.Q ),
    .b(\DFF_96.Q ),
    .s(_0244_),
    .y(\DFF_84.D )
  );
  al_mux2l _0851_ (
    .a(\DFF_172.Q ),
    .b(\DFF_200.Q ),
    .s(_0293_),
    .y(\DFF_172.D )
  );
  al_mux2l _0852_ (
    .a(\DFF_163.Q ),
    .b(\DFF_73.Q ),
    .s(_0244_),
    .y(\DFF_163.D )
  );
  al_mux2l _0853_ (
    .a(\DFF_175.Q ),
    .b(\DFF_74.Q ),
    .s(_0244_),
    .y(\DFF_175.D )
  );
  al_mux2l _0854_ (
    .a(\DFF_57.Q ),
    .b(\DFF_163.Q ),
    .s(_0244_),
    .y(\DFF_57.D )
  );
  al_inv _0855_ (
    .a(\DFF_105.Q ),
    .y(_0354_)
  );
  al_mux2l _0856_ (
    .a(_0009_),
    .b(_0084_),
    .s(_0340_),
    .y(_0355_)
  );
  al_nand3 _0857_ (
    .a(_0330_),
    .b(_0355_),
    .c(_0243_),
    .y(_0356_)
  );
  al_nand2 _0858_ (
    .a(_0354_),
    .b(_0356_),
    .y(_0357_)
  );
  al_mux2l _0859_ (
    .a(_0357_),
    .b(\DFF_129.Q ),
    .s(_0339_),
    .y(\DFF_105.D )
  );
  al_mux2l _0860_ (
    .a(\DFF_73.Q ),
    .b(\DFF_195.Q ),
    .s(_0244_),
    .y(\DFF_73.D )
  );
  al_mux2l _0861_ (
    .a(\DFF_68.Q ),
    .b(\DFF_5.Q ),
    .s(_0244_),
    .y(\DFF_68.D )
  );
  al_mux2l _0862_ (
    .a(\DFF_78.Q ),
    .b(\DFF_57.Q ),
    .s(_0244_),
    .y(\DFF_78.D )
  );
  al_aoi21 _0863_ (
    .a(_0324_),
    .b(_0153_),
    .c(\DFF_24.Q ),
    .y(_0358_)
  );
  al_ao21ftf _0864_ (
    .a(_0358_),
    .b(_0158_),
    .c(_0159_),
    .y(\DFF_24.D )
  );
  al_mux2l _0865_ (
    .a(\DFF_102.Q ),
    .b(\DFF_208.Q ),
    .s(_0293_),
    .y(\DFF_102.D )
  );
  al_mux2h _0866_ (
    .a(\DFF_113.Q ),
    .b(_0040_),
    .s(_0243_),
    .y(\DFF_113.D )
  );
  al_mux2l _0867_ (
    .a(\DFF_11.Q ),
    .b(\DFF_208.Q ),
    .s(_0339_),
    .y(\DFF_11.D )
  );
  al_and2 _0868_ (
    .a(\DFF_60.Q ),
    .b(_0293_),
    .y(\DFF_60.D )
  );
  al_mux2l _0869_ (
    .a(\DFF_148.Q ),
    .b(\DFF_70.Q ),
    .s(\DFF_11.Q ),
    .y(_0359_)
  );
  al_mux2l _0870_ (
    .a(\DFF_74.Q ),
    .b(_0359_),
    .s(_0244_),
    .y(\DFF_74.D )
  );
  al_mux2l _0871_ (
    .a(\DFF_82.Q ),
    .b(\DFF_208.Q ),
    .s(_0251_),
    .y(\DFF_82.D )
  );
  al_and2 _0872_ (
    .a(\DFF_205.Q ),
    .b(_0339_),
    .y(\DFF_205.D )
  );
  al_and2 _0873_ (
    .a(\DFF_69.D ),
    .b(_0277_),
    .y(_0360_)
  );
  al_nand3 _0874_ (
    .a(\DFF_188.Q ),
    .b(\DFF_175.Q ),
    .c(_0277_),
    .y(_0361_)
  );
  al_aoi21ttf _0875_ (
    .a(g563),
    .b(_0305_),
    .c(_0361_),
    .y(_0362_)
  );
  al_aoi21ttf _0876_ (
    .a(\DFF_68.Q ),
    .b(_0360_),
    .c(_0362_),
    .y(_0363_)
  );
  al_nor3fft _0877_ (
    .a(\DFF_188.Q ),
    .b(_0292_),
    .c(_0262_),
    .y(_0364_)
  );
  al_nand3fft _0878_ (
    .a(_0340_),
    .b(\DFF_188.Q ),
    .c(_0274_),
    .y(_0365_)
  );
  al_aoi21ttf _0879_ (
    .a(\DFF_102.Q ),
    .b(_0364_),
    .c(_0365_),
    .y(_0366_)
  );
  al_or3 _0880_ (
    .a(_0167_),
    .b(_0250_),
    .c(_0262_),
    .y(_0367_)
  );
  al_and3 _0881_ (
    .a(\DFF_131.Q ),
    .b(_0275_),
    .c(_0263_),
    .y(_0368_)
  );
  al_ao21 _0882_ (
    .a(\DFF_135.Q ),
    .b(_0266_),
    .c(_0368_),
    .y(_0369_)
  );
  al_nand3fft _0883_ (
    .a(\DFF_153.Q ),
    .b(\DFF_200.Q ),
    .c(_0268_),
    .y(_0370_)
  );
  al_ao21ttf _0884_ (
    .a(\DFF_173.Q ),
    .b(_0272_),
    .c(_0370_),
    .y(_0371_)
  );
  al_nor3ftt _0885_ (
    .a(_0367_),
    .b(_0371_),
    .c(_0369_),
    .y(_0372_)
  );
  al_nand3 _0886_ (
    .a(_0366_),
    .b(_0372_),
    .c(_0363_),
    .y(_0373_)
  );
  al_ao21 _0887_ (
    .a(\DFF_208.Q ),
    .b(_0260_),
    .c(_0373_),
    .y(_0374_)
  );
  al_nand3 _0888_ (
    .a(\DFF_99.Q ),
    .b(\DFF_201.D ),
    .c(_0257_),
    .y(_0375_)
  );
  al_aoi21ftf _0889_ (
    .a(_0345_),
    .b(\DFF_178.D ),
    .c(_0375_),
    .y(_0376_)
  );
  al_nand3fft _0890_ (
    .a(_0280_),
    .b(_0374_),
    .c(_0376_),
    .y(\DFF_186.D )
  );
  al_mux2l _0891_ (
    .a(\DFF_42.Q ),
    .b(\DFF_84.Q ),
    .s(_0244_),
    .y(\DFF_42.D )
  );
  al_mux2l _0892_ (
    .a(\DFF_204.Q ),
    .b(\DFF_129.Q ),
    .s(_0293_),
    .y(\DFF_204.D )
  );
  al_nand3 _0893_ (
    .a(\DFF_99.Q ),
    .b(\DFF_43.D ),
    .c(_0257_),
    .y(_0377_)
  );
  al_aoi21ftf _0894_ (
    .a(_0345_),
    .b(\DFF_168.D ),
    .c(_0377_),
    .y(_0378_)
  );
  al_and3ftt _0895_ (
    .a(\DFF_69.Q ),
    .b(_0261_),
    .c(_0268_),
    .y(_0379_)
  );
  al_aoi21 _0896_ (
    .a(\DFF_113.Q ),
    .b(_0272_),
    .c(_0379_),
    .y(_0380_)
  );
  al_aoi21ttf _0897_ (
    .a(\DFF_5.Q ),
    .b(_0360_),
    .c(_0380_),
    .y(_0381_)
  );
  al_and3 _0898_ (
    .a(\DFF_59.Q ),
    .b(_0275_),
    .c(_0263_),
    .y(_0382_)
  );
  al_aoi21 _0899_ (
    .a(\DFF_21.Q ),
    .b(_0266_),
    .c(_0382_),
    .y(_0383_)
  );
  al_aoi21ttf _0900_ (
    .a(\DFF_179.Q ),
    .b(_0267_),
    .c(_0383_),
    .y(_0384_)
  );
  al_nand3 _0901_ (
    .a(\DFF_200.Q ),
    .b(g564),
    .c(_0268_),
    .y(_0385_)
  );
  al_nand3 _0902_ (
    .a(\DFF_188.Q ),
    .b(\DFF_74.Q ),
    .c(_0277_),
    .y(_0386_)
  );
  al_and3 _0903_ (
    .a(_0385_),
    .b(_0386_),
    .c(_0384_),
    .y(_0387_)
  );
  al_inv _0904_ (
    .a(\DFF_177.Q ),
    .y(_0388_)
  );
  al_nand3 _0905_ (
    .a(\DFF_69.D ),
    .b(\DFF_205.Q ),
    .c(_0274_),
    .y(_0389_)
  );
  al_aoi21ftf _0906_ (
    .a(_0388_),
    .b(_0364_),
    .c(_0389_),
    .y(_0390_)
  );
  al_and3 _0907_ (
    .a(_0381_),
    .b(_0390_),
    .c(_0387_),
    .y(_0391_)
  );
  al_aoi21ftf _0908_ (
    .a(\DFF_69.D ),
    .b(_0260_),
    .c(_0391_),
    .y(_0392_)
  );
  al_nand3ftt _0909_ (
    .a(_0280_),
    .b(_0392_),
    .c(_0378_),
    .y(\DFF_44.D )
  );
  al_mux2l _0910_ (
    .a(\DFF_94.Q ),
    .b(\DFF_200.Q ),
    .s(_0251_),
    .y(\DFF_94.D )
  );
  al_nand2ft _0911_ (
    .a(\DFF_135.Q ),
    .b(_0110_),
    .y(\DFF_135.D )
  );
  al_mux2l _0912_ (
    .a(\DFF_81.Q ),
    .b(\DFF_68.Q ),
    .s(_0244_),
    .y(\DFF_81.D )
  );
  al_nand2 _0913_ (
    .a(_0388_),
    .b(_0293_),
    .y(\DFF_177.D )
  );
  al_mux2l _0914_ (
    .a(\DFF_195.Q ),
    .b(\DFF_77.Q ),
    .s(_0244_),
    .y(\DFF_195.D )
  );
  al_nand2ft _0915_ (
    .a(\DFF_21.Q ),
    .b(_0029_),
    .y(\DFF_21.D )
  );
  al_oai21ftf _0916_ (
    .a(_0124_),
    .b(\DFF_14.D ),
    .c(\DFF_59.Q ),
    .y(\DFF_59.D )
  );
  al_mux2h _0917_ (
    .a(\DFF_25.Q ),
    .b(_0122_),
    .s(_0243_),
    .y(\DFF_25.D )
  );
  al_ao21 _0918_ (
    .a(\DFF_140.Q ),
    .b(\DFF_144.Q ),
    .c(\DFF_126.Q ),
    .y(_0393_)
  );
  al_oai21ftf _0919_ (
    .a(_0393_),
    .b(_0150_),
    .c(_0155_),
    .y(\DFF_126.D )
  );
  al_nand3 _0920_ (
    .a(\DFF_188.Q ),
    .b(\DFF_195.Q ),
    .c(_0277_),
    .y(_0394_)
  );
  al_aoi21ttf _0921_ (
    .a(\DFF_20.Q ),
    .b(_0272_),
    .c(_0394_),
    .y(_0395_)
  );
  al_aoi21ttf _0922_ (
    .a(\DFF_53.Q ),
    .b(_0360_),
    .c(_0395_),
    .y(_0396_)
  );
  al_nand3 _0923_ (
    .a(\DFF_188.Q ),
    .b(\DFF_204.Q ),
    .c(_0274_),
    .y(_0397_)
  );
  al_nand3fft _0924_ (
    .a(\DFF_188.Q ),
    .b(_0354_),
    .c(_0274_),
    .y(_0398_)
  );
  al_and3 _0925_ (
    .a(\DFF_200.Q ),
    .b(g561),
    .c(_0268_),
    .y(_0399_)
  );
  al_nor3ftt _0926_ (
    .a(\DFF_75.Q ),
    .b(_0250_),
    .c(_0262_),
    .y(_0400_)
  );
  al_and3fft _0927_ (
    .a(_0400_),
    .b(_0399_),
    .c(_0398_),
    .y(_0401_)
  );
  al_nand3 _0928_ (
    .a(_0397_),
    .b(_0401_),
    .c(_0396_),
    .y(_0402_)
  );
  al_ao21 _0929_ (
    .a(\DFF_129.Q ),
    .b(_0260_),
    .c(_0402_),
    .y(_0403_)
  );
  al_nand3 _0930_ (
    .a(\DFF_99.Q ),
    .b(\DFF_134.D ),
    .c(_0257_),
    .y(_0404_)
  );
  al_aoi21ftf _0931_ (
    .a(_0345_),
    .b(\DFF_3.D ),
    .c(_0404_),
    .y(_0405_)
  );
  al_nand3fft _0932_ (
    .a(_0280_),
    .b(_0403_),
    .c(_0405_),
    .y(\DFF_63.D )
  );
  al_nand2ft _0933_ (
    .a(\DFF_182.Q ),
    .b(_0293_),
    .y(\DFF_182.D )
  );
  al_nand2 _0934_ (
    .a(\DFF_139.Q ),
    .b(g567),
    .y(g4121)
  );
  al_nand3 _0935_ (
    .a(\DFF_179.Q ),
    .b(_0039_),
    .c(_0144_),
    .y(_0406_)
  );
  al_or2 _0936_ (
    .a(\DFF_111.Q ),
    .b(\DFF_179.Q ),
    .y(_0407_)
  );
  al_and3 _0937_ (
    .a(_0407_),
    .b(_0296_),
    .c(_0406_),
    .y(_0408_)
  );
  al_nand3 _0938_ (
    .a(\DFF_82.Q ),
    .b(_0121_),
    .c(_0190_),
    .y(_0409_)
  );
  al_or2 _0939_ (
    .a(\DFF_111.Q ),
    .b(\DFF_82.Q ),
    .y(_0410_)
  );
  al_and3 _0940_ (
    .a(_0410_),
    .b(_0300_),
    .c(_0409_),
    .y(_0411_)
  );
  al_nand3 _0941_ (
    .a(\DFF_188.Q ),
    .b(\DFF_182.Q ),
    .c(_0274_),
    .y(_0412_)
  );
  al_nand3 _0942_ (
    .a(\DFF_69.D ),
    .b(\DFF_42.Q ),
    .c(_0277_),
    .y(_0413_)
  );
  al_nand3 _0943_ (
    .a(\DFF_188.Q ),
    .b(\DFF_57.Q ),
    .c(_0277_),
    .y(_0414_)
  );
  al_aoi21ttf _0944_ (
    .a(g558),
    .b(_0305_),
    .c(_0414_),
    .y(_0415_)
  );
  al_and3 _0945_ (
    .a(_0412_),
    .b(_0413_),
    .c(_0415_),
    .y(_0416_)
  );
  al_and3 _0946_ (
    .a(\DFF_111.Q ),
    .b(_0259_),
    .c(_0254_),
    .y(_0417_)
  );
  al_and3fft _0947_ (
    .a(_0417_),
    .b(_0280_),
    .c(_0416_),
    .y(_0418_)
  );
  al_nand3fft _0948_ (
    .a(_0411_),
    .b(_0408_),
    .c(_0418_),
    .y(\DFF_90.D )
  );
  al_buf _0949_ (
    .a(\DFF_44.Q ),
    .y(\DFF_209.D )
  );
  al_buf _0950_ (
    .a(\DFF_79.Q ),
    .y(\DFF_123.D )
  );
  al_buf _0951_ (
    .a(\DFF_187.Q ),
    .y(\DFF_128.D )
  );
  al_buf _0952_ (
    .a(\DFF_167.Q ),
    .y(\DFF_6.D )
  );
  al_buf _0953_ (
    .a(\DFF_27.Q ),
    .y(\DFF_98.D )
  );
  al_buf _0954_ (
    .a(\DFF_90.Q ),
    .y(\DFF_10.D )
  );
  al_buf _0955_ (
    .a(\DFF_186.Q ),
    .y(\DFF_117.D )
  );
  al_buf _0956_ (
    .a(\DFF_63.Q ),
    .y(\DFF_127.D )
  );
  al_dffl _0957_ (
    .clk(CK),
    .d(\DFF_3.D ),
    .q(\DFF_3.Q )
  );
  al_dffl _0958_ (
    .clk(CK),
    .d(\DFF_5.D ),
    .q(\DFF_5.Q )
  );
  al_dffl _0959_ (
    .clk(CK),
    .d(\DFF_6.D ),
    .q(\DFF_6.Q )
  );
  al_dffl _0960_ (
    .clk(CK),
    .d(g39),
    .q(\DFF_9.Q )
  );
  al_dffl _0961_ (
    .clk(CK),
    .d(\DFF_10.D ),
    .q(\DFF_10.Q )
  );
  al_dffl _0962_ (
    .clk(CK),
    .d(\DFF_11.D ),
    .q(\DFF_11.Q )
  );
  al_dffl _0963_ (
    .clk(CK),
    .d(\DFF_14.D ),
    .q(\DFF_14.Q )
  );
  al_dffl _0964_ (
    .clk(CK),
    .d(\DFF_15.D ),
    .q(\DFF_15.Q )
  );
  al_dffl _0965_ (
    .clk(CK),
    .d(\DFF_17.D ),
    .q(\DFF_17.Q )
  );
  al_dffl _0966_ (
    .clk(CK),
    .d(\DFF_19.D ),
    .q(\DFF_19.Q )
  );
  al_dffl _0967_ (
    .clk(CK),
    .d(\DFF_20.D ),
    .q(\DFF_20.Q )
  );
  al_dffl _0968_ (
    .clk(CK),
    .d(\DFF_21.D ),
    .q(\DFF_21.Q )
  );
  al_dffl _0969_ (
    .clk(CK),
    .d(\DFF_23.D ),
    .q(\DFF_23.Q )
  );
  al_dffl _0970_ (
    .clk(CK),
    .d(\DFF_24.D ),
    .q(\DFF_24.Q )
  );
  al_dffl _0971_ (
    .clk(CK),
    .d(\DFF_25.D ),
    .q(\DFF_25.Q )
  );
  al_dffl _0972_ (
    .clk(CK),
    .d(\DFF_6.Q ),
    .q(\DFF_26.Q )
  );
  al_dffl _0973_ (
    .clk(CK),
    .d(\DFF_27.D ),
    .q(\DFF_27.Q )
  );
  al_dffl _0974_ (
    .clk(CK),
    .d(\DFF_28.D ),
    .q(\DFF_28.Q )
  );
  al_dffl _0975_ (
    .clk(CK),
    .d(\DFF_30.D ),
    .q(\DFF_30.Q )
  );
  al_dffl _0976_ (
    .clk(CK),
    .d(\DFF_36.D ),
    .q(\DFF_36.Q )
  );
  al_dffl _0977_ (
    .clk(CK),
    .d(\DFF_37.D ),
    .q(\DFF_37.Q )
  );
  al_dffl _0978_ (
    .clk(CK),
    .d(\DFF_40.D ),
    .q(\DFF_40.Q )
  );
  al_dffl _0979_ (
    .clk(CK),
    .d(\DFF_42.D ),
    .q(\DFF_42.Q )
  );
  al_dffl _0980_ (
    .clk(CK),
    .d(\DFF_43.D ),
    .q(\DFF_43.Q )
  );
  al_dffl _0981_ (
    .clk(CK),
    .d(\DFF_44.D ),
    .q(\DFF_44.Q )
  );
  al_dffl _0982_ (
    .clk(CK),
    .d(g32),
    .q(\DFF_47.Q )
  );
  al_dffl _0983_ (
    .clk(CK),
    .d(\DFF_48.D ),
    .q(\DFF_48.Q )
  );
  al_dffl _0984_ (
    .clk(CK),
    .d(\DFF_50.D ),
    .q(\DFF_50.Q )
  );
  al_dffl _0985_ (
    .clk(CK),
    .d(\DFF_123.Q ),
    .q(\DFF_51.Q )
  );
  al_dffl _0986_ (
    .clk(CK),
    .d(\DFF_52.D ),
    .q(\DFF_52.Q )
  );
  al_dffl _0987_ (
    .clk(CK),
    .d(\DFF_53.D ),
    .q(\DFF_53.Q )
  );
  al_dffl _0988_ (
    .clk(CK),
    .d(\DFF_55.D ),
    .q(\DFF_55.Q )
  );
  al_dffl _0989_ (
    .clk(CK),
    .d(\DFF_57.D ),
    .q(\DFF_57.Q )
  );
  al_dffl _0990_ (
    .clk(CK),
    .d(\DFF_58.D ),
    .q(\DFF_58.Q )
  );
  al_dffl _0991_ (
    .clk(CK),
    .d(\DFF_59.D ),
    .q(\DFF_59.Q )
  );
  al_dffl _0992_ (
    .clk(CK),
    .d(\DFF_60.D ),
    .q(\DFF_60.Q )
  );
  al_dffl _0993_ (
    .clk(CK),
    .d(\DFF_61.D ),
    .q(\DFF_61.Q )
  );
  al_dffl _0994_ (
    .clk(CK),
    .d(\DFF_63.D ),
    .q(\DFF_63.Q )
  );
  al_dffl _0995_ (
    .clk(CK),
    .d(\DFF_64.D ),
    .q(\DFF_64.Q )
  );
  al_dffl _0996_ (
    .clk(CK),
    .d(\DFF_68.D ),
    .q(\DFF_68.Q )
  );
  al_dffl _0997_ (
    .clk(CK),
    .d(\DFF_69.D ),
    .q(\DFF_69.Q )
  );
  al_dffl _0998_ (
    .clk(CK),
    .d(\DFF_148.Q ),
    .q(\DFF_70.Q )
  );
  al_dffl _0999_ (
    .clk(CK),
    .d(\DFF_73.D ),
    .q(\DFF_73.Q )
  );
  al_dffl _1000_ (
    .clk(CK),
    .d(\DFF_74.D ),
    .q(\DFF_74.Q )
  );
  al_dffl _1001_ (
    .clk(CK),
    .d(\DFF_75.D ),
    .q(\DFF_75.Q )
  );
  al_dffl _1002_ (
    .clk(CK),
    .d(g567),
    .q(\DFF_76.Q )
  );
  al_dffl _1003_ (
    .clk(CK),
    .d(\DFF_77.D ),
    .q(\DFF_77.Q )
  );
  al_dffl _1004_ (
    .clk(CK),
    .d(\DFF_78.D ),
    .q(\DFF_78.Q )
  );
  al_dffl _1005_ (
    .clk(CK),
    .d(\DFF_79.D ),
    .q(\DFF_79.Q )
  );
  al_dffl _1006_ (
    .clk(CK),
    .d(\DFF_80.D ),
    .q(\DFF_80.Q )
  );
  al_dffl _1007_ (
    .clk(CK),
    .d(\DFF_81.D ),
    .q(\DFF_81.Q )
  );
  al_dffl _1008_ (
    .clk(CK),
    .d(\DFF_82.D ),
    .q(\DFF_82.Q )
  );
  al_dffl _1009_ (
    .clk(CK),
    .d(\DFF_83.D ),
    .q(\DFF_83.Q )
  );
  al_dffl _1010_ (
    .clk(CK),
    .d(\DFF_84.D ),
    .q(\DFF_84.Q )
  );
  al_dffl _1011_ (
    .clk(CK),
    .d(\DFF_87.D ),
    .q(\DFF_87.Q )
  );
  al_dffl _1012_ (
    .clk(CK),
    .d(\DFF_88.D ),
    .q(\DFF_88.Q )
  );
  al_dffl _1013_ (
    .clk(CK),
    .d(\DFF_89.D ),
    .q(\DFF_89.Q )
  );
  al_dffl _1014_ (
    .clk(CK),
    .d(\DFF_90.D ),
    .q(\DFF_90.Q )
  );
  al_dffl _1015_ (
    .clk(CK),
    .d(g40),
    .q(\DFF_92.Q )
  );
  al_dffl _1016_ (
    .clk(CK),
    .d(\DFF_93.D ),
    .q(\DFF_93.Q )
  );
  al_dffl _1017_ (
    .clk(CK),
    .d(\DFF_94.D ),
    .q(\DFF_94.Q )
  );
  al_dffl _1018_ (
    .clk(CK),
    .d(\DFF_96.D ),
    .q(\DFF_96.Q )
  );
  al_dffl _1019_ (
    .clk(CK),
    .d(\DFF_98.D ),
    .q(\DFF_98.Q )
  );
  al_dffl _1020_ (
    .clk(CK),
    .d(g37),
    .q(\DFF_99.Q )
  );
  al_dffl _1021_ (
    .clk(CK),
    .d(\DFF_102.D ),
    .q(\DFF_102.Q )
  );
  al_dffl _1022_ (
    .clk(CK),
    .d(\DFF_105.D ),
    .q(\DFF_105.Q )
  );
  al_dffl _1023_ (
    .clk(CK),
    .d(\DFF_109.D ),
    .q(\DFF_109.Q )
  );
  al_dffl _1024_ (
    .clk(CK),
    .d(\DFF_110.D ),
    .q(\DFF_110.Q )
  );
  al_dffl _1025_ (
    .clk(CK),
    .d(\DFF_10.Q ),
    .q(\DFF_111.Q )
  );
  al_dffl _1026_ (
    .clk(CK),
    .d(\DFF_113.D ),
    .q(\DFF_113.Q )
  );
  al_dffl _1027_ (
    .clk(CK),
    .d(\DFF_93.Q ),
    .q(\DFF_114.Q )
  );
  al_dffl _1028_ (
    .clk(CK),
    .d(\DFF_170.Q ),
    .q(\DFF_116.Q )
  );
  al_dffl _1029_ (
    .clk(CK),
    .d(\DFF_117.D ),
    .q(\DFF_117.Q )
  );
  al_dffl _1030_ (
    .clk(CK),
    .d(\DFF_121.D ),
    .q(\DFF_121.Q )
  );
  al_dffl _1031_ (
    .clk(CK),
    .d(\DFF_123.D ),
    .q(\DFF_123.Q )
  );
  al_dffl _1032_ (
    .clk(CK),
    .d(g38),
    .q(\DFF_124.Q )
  );
  al_dffl _1033_ (
    .clk(CK),
    .d(\DFF_125.D ),
    .q(\DFF_125.Q )
  );
  al_dffl _1034_ (
    .clk(CK),
    .d(\DFF_126.D ),
    .q(\DFF_126.Q )
  );
  al_dffl _1035_ (
    .clk(CK),
    .d(\DFF_127.D ),
    .q(\DFF_127.Q )
  );
  al_dffl _1036_ (
    .clk(CK),
    .d(\DFF_128.D ),
    .q(\DFF_128.Q )
  );
  al_dffl _1037_ (
    .clk(CK),
    .d(\DFF_127.Q ),
    .q(\DFF_129.Q )
  );
  al_dffl _1038_ (
    .clk(CK),
    .d(\DFF_131.D ),
    .q(\DFF_131.Q )
  );
  al_dffl _1039_ (
    .clk(CK),
    .d(g45),
    .q(\DFF_132.Q )
  );
  al_dffl _1040_ (
    .clk(CK),
    .d(\DFF_134.D ),
    .q(\DFF_134.Q )
  );
  al_dffl _1041_ (
    .clk(CK),
    .d(\DFF_135.D ),
    .q(\DFF_135.Q )
  );
  al_dffl _1042_ (
    .clk(CK),
    .d(\DFF_132.Q ),
    .q(\DFF_139.Q )
  );
  al_dffl _1043_ (
    .clk(CK),
    .d(\DFF_140.D ),
    .q(\DFF_140.Q )
  );
  al_dffl _1044_ (
    .clk(CK),
    .d(\DFF_141.D ),
    .q(\DFF_141.Q )
  );
  al_dffl _1045_ (
    .clk(CK),
    .d(\DFF_142.D ),
    .q(\DFF_142.Q )
  );
  al_dffl _1046_ (
    .clk(CK),
    .d(g42),
    .q(\DFF_143.Q )
  );
  al_dffl _1047_ (
    .clk(CK),
    .d(\DFF_144.D ),
    .q(\DFF_144.Q )
  );
  al_dffl _1048_ (
    .clk(CK),
    .d(\DFF_146.D ),
    .q(\DFF_146.Q )
  );
  al_dffl _1049_ (
    .clk(CK),
    .d(g702),
    .q(\DFF_147.Q )
  );
  al_dffl _1050_ (
    .clk(CK),
    .d(\DFF_143.Q ),
    .q(\DFF_148.Q )
  );
  al_dffl _1051_ (
    .clk(CK),
    .d(\DFF_151.D ),
    .q(\DFF_151.Q )
  );
  al_dffl _1052_ (
    .clk(CK),
    .d(\DFF_58.Q ),
    .q(\DFF_152.Q )
  );
  al_dffl _1053_ (
    .clk(CK),
    .d(\DFF_153.D ),
    .q(\DFF_153.Q )
  );
  al_dffl _1054_ (
    .clk(CK),
    .d(\DFF_154.D ),
    .q(\DFF_154.Q )
  );
  al_dffl _1055_ (
    .clk(CK),
    .d(\DFF_19.Q ),
    .q(\DFF_156.Q )
  );
  al_dffl _1056_ (
    .clk(CK),
    .d(\DFF_30.Q ),
    .q(\DFF_157.Q )
  );
  al_dffl _1057_ (
    .clk(CK),
    .d(\DFF_158.D ),
    .q(\DFF_158.Q )
  );
  al_dffl _1058_ (
    .clk(CK),
    .d(\DFF_161.D ),
    .q(\DFF_161.Q )
  );
  al_dffl _1059_ (
    .clk(CK),
    .d(\DFF_163.D ),
    .q(\DFF_163.Q )
  );
  al_dffl _1060_ (
    .clk(CK),
    .d(\DFF_164.D ),
    .q(\DFF_164.Q )
  );
  al_dffl _1061_ (
    .clk(CK),
    .d(\DFF_141.Q ),
    .q(\DFF_166.Q )
  );
  al_dffl _1062_ (
    .clk(CK),
    .d(\DFF_167.D ),
    .q(\DFF_167.Q )
  );
  al_dffl _1063_ (
    .clk(CK),
    .d(\DFF_168.D ),
    .q(\DFF_168.Q )
  );
  al_dffl _1064_ (
    .clk(CK),
    .d(\DFF_169.D ),
    .q(\DFF_169.Q )
  );
  al_dffl _1065_ (
    .clk(CK),
    .d(\DFF_170.D ),
    .q(\DFF_170.Q )
  );
  al_dffl _1066_ (
    .clk(CK),
    .d(\DFF_172.D ),
    .q(\DFF_172.Q )
  );
  al_dffl _1067_ (
    .clk(CK),
    .d(\DFF_173.D ),
    .q(\DFF_173.Q )
  );
  al_dffl _1068_ (
    .clk(CK),
    .d(\DFF_175.D ),
    .q(\DFF_175.Q )
  );
  al_dffl _1069_ (
    .clk(CK),
    .d(\DFF_28.Q ),
    .q(\DFF_176.Q )
  );
  al_dffl _1070_ (
    .clk(CK),
    .d(\DFF_177.D ),
    .q(\DFF_177.Q )
  );
  al_dffl _1071_ (
    .clk(CK),
    .d(\DFF_178.D ),
    .q(\DFF_178.Q )
  );
  al_dffl _1072_ (
    .clk(CK),
    .d(\DFF_179.D ),
    .q(\DFF_179.Q )
  );
  al_dffl _1073_ (
    .clk(CK),
    .d(g46),
    .q(\DFF_180.Q )
  );
  al_dffl _1074_ (
    .clk(CK),
    .d(\DFF_182.D ),
    .q(\DFF_182.Q )
  );
  al_dffl _1075_ (
    .clk(CK),
    .d(\DFF_89.Q ),
    .q(\DFF_183.Q )
  );
  al_dffl _1076_ (
    .clk(CK),
    .d(\DFF_186.D ),
    .q(\DFF_186.Q )
  );
  al_dffl _1077_ (
    .clk(CK),
    .d(\DFF_187.D ),
    .q(\DFF_187.Q )
  );
  al_dffl _1078_ (
    .clk(CK),
    .d(\DFF_209.Q ),
    .q(\DFF_188.Q )
  );
  al_dffl _1079_ (
    .clk(CK),
    .d(\DFF_189.D ),
    .q(\DFF_189.Q )
  );
  al_dffl _1080_ (
    .clk(CK),
    .d(\DFF_190.D ),
    .q(\DFF_190.Q )
  );
  al_dffl _1081_ (
    .clk(CK),
    .d(\DFF_191.D ),
    .q(\DFF_191.Q )
  );
  al_dffl _1082_ (
    .clk(CK),
    .d(\DFF_195.D ),
    .q(\DFF_195.Q )
  );
  al_dffl _1083_ (
    .clk(CK),
    .d(\DFF_196.D ),
    .q(\DFF_196.Q )
  );
  al_dffl _1084_ (
    .clk(CK),
    .d(\DFF_197.D ),
    .q(\DFF_197.Q )
  );
  al_dffl _1085_ (
    .clk(CK),
    .d(\DFF_98.Q ),
    .q(\DFF_200.Q )
  );
  al_dffl _1086_ (
    .clk(CK),
    .d(\DFF_201.D ),
    .q(\DFF_201.Q )
  );
  al_dffl _1087_ (
    .clk(CK),
    .d(\DFF_204.D ),
    .q(\DFF_204.Q )
  );
  al_dffl _1088_ (
    .clk(CK),
    .d(\DFF_205.D ),
    .q(\DFF_205.Q )
  );
  al_dffl _1089_ (
    .clk(CK),
    .d(\DFF_128.Q ),
    .q(\DFF_207.Q )
  );
  al_dffl _1090_ (
    .clk(CK),
    .d(\DFF_117.Q ),
    .q(\DFF_208.Q )
  );
  al_dffl _1091_ (
    .clk(CK),
    .d(\DFF_209.D ),
    .q(\DFF_209.Q )
  );
  assign \DFF_0.CK  = CK;
  assign \DFF_0.D  = \DFF_117.Q ;
  assign \DFF_0.Q  = \DFF_208.Q ;
  assign \DFF_1.CK  = CK;
  assign \DFF_10.CK  = CK;
  assign \DFF_100.CK  = CK;
  assign \DFF_101.CK  = CK;
  assign \DFF_102.CK  = CK;
  assign \DFF_103.CK  = CK;
  assign \DFF_103.D  = g42;
  assign \DFF_103.Q  = \DFF_143.Q ;
  assign \DFF_104.CK  = CK;
  assign \DFF_105.CK  = CK;
  assign \DFF_106.CK  = CK;
  assign \DFF_107.CK  = CK;
  assign \DFF_108.CK  = CK;
  assign \DFF_108.D  = \DFF_10.Q ;
  assign \DFF_108.Q  = \DFF_111.Q ;
  assign \DFF_109.CK  = CK;
  assign \DFF_11.CK  = CK;
  assign \DFF_110.CK  = CK;
  assign \DFF_111.CK  = CK;
  assign \DFF_111.D  = \DFF_10.Q ;
  assign \DFF_112.CK  = CK;
  assign \DFF_113.CK  = CK;
  assign \DFF_114.CK  = CK;
  assign \DFF_114.D  = \DFF_93.Q ;
  assign \DFF_115.CK  = CK;
  assign \DFF_116.CK  = CK;
  assign \DFF_116.D  = \DFF_170.Q ;
  assign \DFF_117.CK  = CK;
  assign \DFF_118.CK  = CK;
  assign \DFF_118.D  = \DFF_141.Q ;
  assign \DFF_118.Q  = \DFF_166.Q ;
  assign \DFF_119.CK  = CK;
  assign \DFF_12.CK  = CK;
  assign \DFF_120.CK  = CK;
  assign \DFF_121.CK  = CK;
  assign \DFF_122.CK  = CK;
  assign \DFF_122.D  = \DFF_98.Q ;
  assign \DFF_122.Q  = \DFF_200.Q ;
  assign \DFF_123.CK  = CK;
  assign \DFF_124.CK  = CK;
  assign \DFF_124.D  = g38;
  assign \DFF_125.CK  = CK;
  assign \DFF_126.CK  = CK;
  assign \DFF_127.CK  = CK;
  assign \DFF_128.CK  = CK;
  assign \DFF_129.CK  = CK;
  assign \DFF_129.D  = \DFF_127.Q ;
  assign \DFF_13.CK  = CK;
  assign \DFF_13.D  = \DFF_93.Q ;
  assign \DFF_13.Q  = \DFF_114.Q ;
  assign \DFF_130.CK  = CK;
  assign \DFF_131.CK  = CK;
  assign \DFF_132.CK  = CK;
  assign \DFF_132.D  = g45;
  assign \DFF_133.CK  = CK;
  assign \DFF_134.CK  = CK;
  assign \DFF_135.CK  = CK;
  assign \DFF_136.CK  = CK;
  assign \DFF_137.CK  = CK;
  assign \DFF_137.D  = g36;
  assign \DFF_138.CK  = CK;
  assign \DFF_138.D  = \DFF_28.Q ;
  assign \DFF_138.Q  = \DFF_176.Q ;
  assign \DFF_139.CK  = CK;
  assign \DFF_139.D  = \DFF_132.Q ;
  assign \DFF_14.CK  = CK;
  assign \DFF_140.CK  = CK;
  assign \DFF_141.CK  = CK;
  assign \DFF_142.CK  = CK;
  assign \DFF_143.CK  = CK;
  assign \DFF_143.D  = g42;
  assign \DFF_144.CK  = CK;
  assign \DFF_145.CK  = CK;
  assign \DFF_146.CK  = CK;
  assign \DFF_147.CK  = CK;
  assign \DFF_147.D  = g702;
  assign \DFF_148.CK  = CK;
  assign \DFF_148.D  = \DFF_143.Q ;
  assign \DFF_149.CK  = CK;
  assign \DFF_15.CK  = CK;
  assign \DFF_150.CK  = CK;
  assign \DFF_151.CK  = CK;
  assign \DFF_152.CK  = CK;
  assign \DFF_152.D  = \DFF_58.Q ;
  assign \DFF_153.CK  = CK;
  assign \DFF_154.CK  = CK;
  assign \DFF_155.CK  = CK;
  assign \DFF_156.CK  = CK;
  assign \DFF_156.D  = \DFF_19.Q ;
  assign \DFF_157.CK  = CK;
  assign \DFF_157.D  = \DFF_30.Q ;
  assign \DFF_158.CK  = CK;
  assign \DFF_159.CK  = CK;
  assign \DFF_16.CK  = CK;
  assign \DFF_160.CK  = CK;
  assign \DFF_161.CK  = CK;
  assign \DFF_162.CK  = CK;
  assign \DFF_163.CK  = CK;
  assign \DFF_164.CK  = CK;
  assign \DFF_165.CK  = CK;
  assign \DFF_166.CK  = CK;
  assign \DFF_166.D  = \DFF_141.Q ;
  assign \DFF_167.CK  = CK;
  assign \DFF_168.CK  = CK;
  assign \DFF_169.CK  = CK;
  assign \DFF_17.CK  = CK;
  assign \DFF_170.CK  = CK;
  assign \DFF_171.CK  = CK;
  assign \DFF_172.CK  = CK;
  assign \DFF_173.CK  = CK;
  assign \DFF_174.CK  = CK;
  assign \DFF_175.CK  = CK;
  assign \DFF_176.CK  = CK;
  assign \DFF_176.D  = \DFF_28.Q ;
  assign \DFF_177.CK  = CK;
  assign \DFF_178.CK  = CK;
  assign \DFF_179.CK  = CK;
  assign \DFF_18.CK  = CK;
  assign \DFF_180.CK  = CK;
  assign \DFF_180.D  = g46;
  assign \DFF_181.CK  = CK;
  assign \DFF_182.CK  = CK;
  assign \DFF_183.CK  = CK;
  assign \DFF_183.D  = \DFF_89.Q ;
  assign \DFF_184.CK  = CK;
  assign \DFF_185.CK  = CK;
  assign \DFF_186.CK  = CK;
  assign \DFF_187.CK  = CK;
  assign \DFF_188.CK  = CK;
  assign \DFF_188.D  = \DFF_209.Q ;
  assign \DFF_189.CK  = CK;
  assign \DFF_19.CK  = CK;
  assign \DFF_190.CK  = CK;
  assign \DFF_191.CK  = CK;
  assign \DFF_192.CK  = CK;
  assign \DFF_193.CK  = CK;
  assign \DFF_194.CK  = CK;
  assign \DFF_195.CK  = CK;
  assign \DFF_196.CK  = CK;
  assign \DFF_197.CK  = CK;
  assign \DFF_198.CK  = CK;
  assign \DFF_199.CK  = CK;
  assign \DFF_2.CK  = CK;
  assign \DFF_20.CK  = CK;
  assign \DFF_200.CK  = CK;
  assign \DFF_200.D  = \DFF_98.Q ;
  assign \DFF_201.CK  = CK;
  assign \DFF_202.CK  = CK;
  assign \DFF_203.CK  = CK;
  assign \DFF_204.CK  = CK;
  assign \DFF_205.CK  = CK;
  assign \DFF_206.CK  = CK;
  assign \DFF_207.CK  = CK;
  assign \DFF_207.D  = \DFF_128.Q ;
  assign \DFF_208.CK  = CK;
  assign \DFF_208.D  = \DFF_117.Q ;
  assign \DFF_209.CK  = CK;
  assign \DFF_21.CK  = CK;
  assign \DFF_210.CK  = CK;
  assign \DFF_22.CK  = CK;
  assign \DFF_23.CK  = CK;
  assign \DFF_24.CK  = CK;
  assign \DFF_25.CK  = CK;
  assign \DFF_26.CK  = CK;
  assign \DFF_26.D  = \DFF_6.Q ;
  assign \DFF_27.CK  = CK;
  assign \DFF_28.CK  = CK;
  assign \DFF_29.CK  = CK;
  assign \DFF_3.CK  = CK;
  assign \DFF_30.CK  = CK;
  assign \DFF_31.CK  = CK;
  assign \DFF_32.CK  = CK;
  assign \DFF_33.CK  = CK;
  assign \DFF_33.D  = \DFF_30.Q ;
  assign \DFF_33.Q  = \DFF_157.Q ;
  assign \DFF_34.CK  = CK;
  assign \DFF_35.CK  = CK;
  assign \DFF_35.D  = \DFF_123.Q ;
  assign \DFF_35.Q  = \DFF_51.Q ;
  assign \DFF_36.CK  = CK;
  assign \DFF_37.CK  = CK;
  assign \DFF_38.CK  = CK;
  assign \DFF_38.D  = \DFF_170.Q ;
  assign \DFF_38.Q  = \DFF_116.Q ;
  assign \DFF_39.CK  = CK;
  assign \DFF_4.CK  = CK;
  assign \DFF_4.D  = \DFF_6.Q ;
  assign \DFF_4.Q  = \DFF_26.Q ;
  assign \DFF_40.CK  = CK;
  assign \DFF_41.CK  = CK;
  assign \DFF_41.D  = \DFF_128.Q ;
  assign \DFF_41.Q  = \DFF_207.Q ;
  assign \DFF_42.CK  = CK;
  assign \DFF_43.CK  = CK;
  assign \DFF_44.CK  = CK;
  assign \DFF_45.CK  = CK;
  assign \DFF_46.CK  = CK;
  assign \DFF_46.D  = \DFF_58.Q ;
  assign \DFF_46.Q  = \DFF_152.Q ;
  assign \DFF_47.CK  = CK;
  assign \DFF_47.D  = g32;
  assign \DFF_48.CK  = CK;
  assign \DFF_49.CK  = CK;
  assign \DFF_5.CK  = CK;
  assign \DFF_50.CK  = CK;
  assign \DFF_51.CK  = CK;
  assign \DFF_51.D  = \DFF_123.Q ;
  assign \DFF_52.CK  = CK;
  assign \DFF_53.CK  = CK;
  assign \DFF_54.CK  = CK;
  assign \DFF_55.CK  = CK;
  assign \DFF_56.CK  = CK;
  assign \DFF_56.D  = g567;
  assign \DFF_56.Q  = \DFF_76.Q ;
  assign \DFF_57.CK  = CK;
  assign \DFF_58.CK  = CK;
  assign \DFF_59.CK  = CK;
  assign \DFF_6.CK  = CK;
  assign \DFF_60.CK  = CK;
  assign \DFF_61.CK  = CK;
  assign \DFF_62.CK  = CK;
  assign \DFF_63.CK  = CK;
  assign \DFF_64.CK  = CK;
  assign \DFF_65.CK  = CK;
  assign \DFF_66.CK  = CK;
  assign \DFF_66.D  = \DFF_127.Q ;
  assign \DFF_66.Q  = \DFF_129.Q ;
  assign \DFF_67.CK  = CK;
  assign \DFF_68.CK  = CK;
  assign \DFF_69.CK  = CK;
  assign \DFF_7.CK  = CK;
  assign \DFF_7.D  = \DFF_89.Q ;
  assign \DFF_7.Q  = \DFF_183.Q ;
  assign \DFF_70.CK  = CK;
  assign \DFF_70.D  = \DFF_148.Q ;
  assign \DFF_71.CK  = CK;
  assign \DFF_72.CK  = CK;
  assign \DFF_72.D  = \DFF_19.Q ;
  assign \DFF_72.Q  = \DFF_156.Q ;
  assign \DFF_73.CK  = CK;
  assign \DFF_74.CK  = CK;
  assign \DFF_75.CK  = CK;
  assign \DFF_76.CK  = CK;
  assign \DFF_76.D  = g567;
  assign \DFF_77.CK  = CK;
  assign \DFF_78.CK  = CK;
  assign \DFF_79.CK  = CK;
  assign \DFF_8.CK  = CK;
  assign \DFF_80.CK  = CK;
  assign \DFF_81.CK  = CK;
  assign \DFF_82.CK  = CK;
  assign \DFF_83.CK  = CK;
  assign \DFF_84.CK  = CK;
  assign \DFF_85.CK  = CK;
  assign \DFF_85.D  = \DFF_143.Q ;
  assign \DFF_85.Q  = \DFF_148.Q ;
  assign \DFF_86.CK  = CK;
  assign \DFF_87.CK  = CK;
  assign \DFF_88.CK  = CK;
  assign \DFF_89.CK  = CK;
  assign \DFF_9.CK  = CK;
  assign \DFF_9.D  = g39;
  assign \DFF_90.CK  = CK;
  assign \DFF_91.CK  = CK;
  assign \DFF_92.CK  = CK;
  assign \DFF_92.D  = g40;
  assign \DFF_93.CK  = CK;
  assign \DFF_94.CK  = CK;
  assign \DFF_95.CK  = CK;
  assign \DFF_95.D  = \DFF_209.Q ;
  assign \DFF_95.Q  = \DFF_188.Q ;
  assign \DFF_96.CK  = CK;
  assign \DFF_97.CK  = CK;
  assign \DFF_98.CK  = CK;
  assign \DFF_99.CK  = CK;
  assign \DFF_99.D  = g37;
  assign I2029 = \DFF_69.D ;
  assign I2033 = \DFF_153.D ;
  assign I2165 = \DFF_69.D ;
  assign I2172 = \DFF_153.D ;
  assign I2290 = \DFF_169.Q ;
  assign I2293 = \DFF_169.Q ;
  assign I2296 = g23;
  assign I2306 = g22;
  assign I2312 = g41;
  assign I2321 = g47;
  assign I2364 = \DFF_153.D ;
  assign I2370 = \DFF_69.D ;
  assign I2373 = \DFF_153.D ;
  assign I2379 = \DFF_69.D ;
  assign I2388 = g639;
  assign I2445 = \DFF_169.Q ;
  assign I2449 = \DFF_169.Q ;
  assign I2453 = \DFF_69.D ;
  assign I2460 = \DFF_69.D ;
  assign I2464 = \DFF_140.Q ;
  assign I2473 = \DFF_169.Q ;
  assign I2476 = \DFF_169.Q ;
  assign I2479 = \DFF_197.Q ;
  assign I2521 = \DFF_147.Q ;
  assign I2537 = \DFF_169.Q ;
  assign I2552 = \DFF_169.Q ;
  assign I2584 = g567;
  assign I2596 = \DFF_139.Q ;
  assign I2608 = \DFF_153.D ;
  assign I2614 = \DFF_69.D ;
  assign I2627 = \DFF_179.Q ;
  assign I2630 = \DFF_153.D ;
  assign I2635 = \DFF_82.Q ;
  assign I2638 = \DFF_69.D ;
  assign I2643 = \DFF_153.D ;
  assign I2716 = g40;
  assign I2731 = g32;
  assign I2735 = g36;
  assign I2753 = g37;
  assign I2756 = g42;
  assign I2773 = g38;
  assign I2776 = g44;
  assign I2802 = g39;
  assign I2805 = g45;
  assign I2821 = g46;
  assign I2825 = \DFF_153.D ;
  assign I2839 = \DFF_69.D ;
  assign I2867 = \DFF_153.D ;
  assign I2877 = \DFF_69.D ;
  assign I2880 = \DFF_153.D ;
  assign I2883 = \DFF_153.D ;
  assign I2887 = \DFF_69.D ;
  assign I2890 = \DFF_69.D ;
  assign I2907 = \DFF_197.Q ;
  assign I2910 = \DFF_69.D ;
  assign I2916 = \DFF_153.D ;
  assign I2929 = \DFF_69.D ;
  assign I2940 = \DFF_153.D ;
  assign I2943 = g40;
  assign I2946 = \DFF_188.Q ;
  assign I2952 = \DFF_208.Q ;
  assign I2955 = g32;
  assign I2961 = g36;
  assign I2982 = \DFF_169.Q ;
  assign I2992 = g37;
  assign I2995 = g42;
  assign I3004 = \DFF_169.Q ;
  assign I3007 = \DFF_169.Q ;
  assign I3016 = g38;
  assign I3019 = g44;
  assign I3022 = \DFF_169.Q ;
  assign I3025 = \DFF_169.Q ;
  assign I3037 = g39;
  assign I3040 = g45;
  assign I3047 = \DFF_169.Q ;
  assign I3050 = \DFF_169.Q ;
  assign I3062 = g46;
  assign I3065 = \DFF_169.Q ;
  assign I3068 = \DFF_169.Q ;
  assign I3074 = \DFF_169.Q ;
  assign I3077 = \DFF_169.Q ;
  assign I3083 = \DFF_169.Q ;
  assign I3086 = \DFF_169.Q ;
  assign I3093 = \DFF_169.Q ;
  assign I3096 = \DFF_169.Q ;
  assign I3102 = \DFF_169.Q ;
  assign I3105 = \DFF_169.Q ;
  assign I3112 = \DFF_169.Q ;
  assign I3137 = g23;
  assign I3140 = g22;
  assign I3144 = g41;
  assign I3152 = g47;
  assign I3198 = \DFF_69.D ;
  assign I3202 = \DFF_153.D ;
  assign I3206 = \DFF_69.D ;
  assign I3215 = \DFF_153.D ;
  assign I3251 = \DFF_140.Q ;
  assign I3255 = \DFF_179.Q ;
  assign I3268 = \DFF_82.Q ;
  assign I3278 = \DFF_6.Q ;
  assign I3284 = \DFF_10.Q ;
  assign I3288 = \DFF_209.Q ;
  assign I3291 = \DFF_123.Q ;
  assign I3294 = \DFF_117.Q ;
  assign I3298 = \DFF_98.Q ;
  assign I3301 = \DFF_127.Q ;
  assign I3304 = \DFF_128.Q ;
  assign I3307 = \DFF_69.D ;
  assign I3313 = \DFF_153.D ;
  assign I3316 = \DFF_69.D ;
  assign I3325 = \DFF_153.D ;
  assign I3434 = g567;
  assign I3452 = \DFF_69.D ;
  assign I3462 = \DFF_69.D ;
  assign I3471 = \DFF_69.D ;
  assign I3474 = \DFF_69.D ;
  assign I3478 = \DFF_69.D ;
  assign I3481 = \DFF_69.D ;
  assign I3485 = \DFF_69.D ;
  assign I3488 = \DFF_169.Q ;
  assign I3493 = \DFF_69.D ;
  assign I3496 = \DFF_23.Q ;
  assign I3499 = \DFF_69.D ;
  assign I3502 = \DFF_169.Q ;
  assign I3505 = \DFF_169.Q ;
  assign I3509 = \DFF_69.D ;
  assign I3513 = \DFF_69.D ;
  assign I3516 = \DFF_169.Q ;
  assign I3519 = \DFF_169.Q ;
  assign I3522 = \DFF_153.D ;
  assign I3525 = \DFF_69.D ;
  assign I3534 = \DFF_169.Q ;
  assign I3537 = \DFF_169.Q ;
  assign I3543 = \DFF_69.D ;
  assign I3550 = \DFF_169.Q ;
  assign I3553 = \DFF_169.Q ;
  assign I3556 = \DFF_169.Q ;
  assign I3563 = \DFF_69.D ;
  assign I3569 = \DFF_69.D ;
  assign I3572 = \DFF_169.Q ;
  assign I3575 = \DFF_169.Q ;
  assign I3578 = \DFF_169.Q ;
  assign I3581 = \DFF_169.Q ;
  assign I3587 = \DFF_69.D ;
  assign I3590 = \DFF_153.D ;
  assign I3593 = \DFF_169.Q ;
  assign I3596 = \DFF_169.Q ;
  assign I3599 = \DFF_169.Q ;
  assign I3602 = \DFF_169.Q ;
  assign I3608 = \DFF_69.D ;
  assign I3614 = \DFF_169.Q ;
  assign I3617 = \DFF_169.Q ;
  assign I3620 = \DFF_169.Q ;
  assign I3623 = \DFF_169.Q ;
  assign I3632 = \DFF_169.Q ;
  assign I3635 = \DFF_169.Q ;
  assign I3638 = \DFF_169.Q ;
  assign I3641 = \DFF_169.Q ;
  assign I3650 = \DFF_179.Q ;
  assign I3653 = \DFF_169.Q ;
  assign I3656 = \DFF_169.Q ;
  assign I3659 = \DFF_169.Q ;
  assign I3665 = \DFF_69.D ;
  assign I3672 = \DFF_82.Q ;
  assign I3675 = \DFF_169.Q ;
  assign I3681 = \DFF_153.D ;
  assign I3711 = \DFF_188.Q ;
  assign I3714 = \DFF_208.Q ;
  assign I3726 = g23;
  assign I3729 = \DFF_69.D ;
  assign I3733 = g22;
  assign I3736 = \DFF_153.D ;
  assign I3746 = g41;
  assign I3755 = \DFF_179.Q ;
  assign I3758 = g47;
  assign I3767 = \DFF_179.Q ;
  assign I3770 = \DFF_82.Q ;
  assign I3779 = \DFF_179.Q ;
  assign I3782 = \DFF_82.Q ;
  assign I3785 = \DFF_23.Q ;
  assign I3797 = \DFF_179.Q ;
  assign I3800 = \DFF_82.Q ;
  assign I3808 = \DFF_179.Q ;
  assign I3811 = \DFF_82.Q ;
  assign I3823 = \DFF_179.Q ;
  assign I3826 = \DFF_82.Q ;
  assign I3836 = \DFF_69.D ;
  assign I3840 = \DFF_179.Q ;
  assign I3843 = \DFF_82.Q ;
  assign I3855 = \DFF_69.D ;
  assign I3861 = \DFF_153.D ;
  assign I3868 = \DFF_179.Q ;
  assign I3871 = \DFF_82.Q ;
  assign I3883 = \DFF_153.D ;
  assign I3890 = \DFF_82.Q ;
  assign I4019 = \DFF_69.D ;
  assign I4031 = \DFF_153.D ;
  assign I4170 = \DFF_6.Q ;
  assign I4189 = \DFF_10.Q ;
  assign I4192 = g40;
  assign I4217 = \DFF_209.Q ;
  assign I4220 = \DFF_123.Q ;
  assign I4226 = \DFF_179.Q ;
  assign I4240 = \DFF_117.Q ;
  assign I4243 = g32;
  assign I4249 = \DFF_179.Q ;
  assign I4252 = \DFF_82.Q ;
  assign I4258 = \DFF_98.Q ;
  assign I4261 = g36;
  assign I4267 = \DFF_179.Q ;
  assign I4270 = \DFF_82.Q ;
  assign I4276 = \DFF_127.Q ;
  assign I4282 = \DFF_179.Q ;
  assign I4285 = \DFF_82.Q ;
  assign I4294 = \DFF_179.Q ;
  assign I4297 = \DFF_82.Q ;
  assign I4303 = g37;
  assign I4306 = g42;
  assign I4309 = \DFF_179.Q ;
  assign I4312 = \DFF_82.Q ;
  assign I4318 = \DFF_128.Q ;
  assign I4321 = g38;
  assign I4324 = g44;
  assign I4327 = \DFF_179.Q ;
  assign I4331 = \DFF_82.Q ;
  assign I4337 = g39;
  assign I4340 = g45;
  assign I4343 = \DFF_179.Q ;
  assign I4347 = \DFF_82.Q ;
  assign I4354 = g46;
  assign I4358 = \DFF_179.Q ;
  assign I4362 = \DFF_82.Q ;
  assign I4371 = \DFF_82.Q ;
  assign I4398 = \DFF_69.D ;
  assign I4410 = \DFF_153.D ;
  assign I4414 = \DFF_69.D ;
  assign I4424 = \DFF_153.D ;
  assign I4468 = g564;
  assign I4903 = g564;
  assign I5337 = \DFF_191.D ;
  assign I5415 = g564;
  assign I5418 = \DFF_191.D ;
  assign I5542 = g47;
  assign I5929 = g47;
  assign g1 = \DFF_209.Q ;
  assign g10 = \DFF_127.Q ;
  assign g1001 = \DFF_207.Q ;
  assign g1006 = \DFF_26.Q ;
  assign g1011 = \DFF_111.Q ;
  assign g1017 = \DFF_51.Q ;
  assign g1030 = \DFF_47.Q ;
  assign g1049 = \DFF_80.D ;
  assign g1076 = \DFF_99.Q ;
  assign g1088 = \DFF_124.Q ;
  assign g1094 = \DFF_9.Q ;
  assign g11 = \DFF_27.Q ;
  assign g1101 = \DFF_92.Q ;
  assign g1106 = \DFF_6.Q ;
  assign g1107 = \DFF_10.Q ;
  assign g1108 = g705;
  assign g1109 = \DFF_209.Q ;
  assign g1110 = \DFF_123.Q ;
  assign g1111 = \DFF_117.Q ;
  assign g1113 = \DFF_98.Q ;
  assign g1114 = \DFF_127.Q ;
  assign g1116 = \DFF_128.Q ;
  assign g1119 = \DFF_11.Q ;
  assign g1122 = \DFF_179.Q ;
  assign g1123 = \DFF_188.Q ;
  assign g1142 = \DFF_82.Q ;
  assign g1143 = \DFF_208.Q ;
  assign g1156 = \DFF_167.Q ;
  assign g1160 = \DFF_94.Q ;
  assign g1161 = \DFF_200.Q ;
  assign g1173 = \DFF_90.Q ;
  assign g1176 = \DFF_75.Q ;
  assign g1177 = \DFF_129.Q ;
  assign g1189 = \DFF_44.Q ;
  assign g1190 = \DFF_79.Q ;
  assign g1193 = \DFF_207.Q ;
  assign g1203 = \DFF_186.Q ;
  assign g1209 = \DFF_26.Q ;
  assign g1219 = \DFF_27.Q ;
  assign g1220 = \DFF_48.Q ;
  assign g1222 = \DFF_111.Q ;
  assign g1232 = \DFF_63.Q ;
  assign g1233 = \DFF_11.Q ;
  assign g1236 = \DFF_51.Q ;
  assign g1246 = \DFF_11.Q ;
  assign g1249 = \DFF_187.Q ;
  assign g1256 = g564;
  assign g1257 = \DFF_189.Q ;
  assign g1263 = \DFF_88.Q ;
  assign g1267 = \DFF_83.Q ;
  assign g1270 = \DFF_158.Q ;
  assign g1273 = g567;
  assign g1274 = \DFF_93.Q ;
  assign g1275 = \DFF_89.Q ;
  assign g1276 = \DFF_24.Q ;
  assign g1279 = \DFF_151.Q ;
  assign g1282 = \DFF_19.Q ;
  assign g1283 = \DFF_141.Q ;
  assign g1284 = \DFF_28.Q ;
  assign g1285 = \DFF_58.Q ;
  assign g1286 = \DFF_30.Q ;
  assign g1287 = \DFF_170.Q ;
  assign g1288 = \DFF_143.Q ;
  assign g1289 = \DFF_132.Q ;
  assign g1290 = \DFF_180.Q ;
  assign g1291 = \DFF_148.Q ;
  assign g1292 = \DFF_143.Q ;
  assign g1293 = \DFF_191.Q ;
  assign g1294 = g702;
  assign g1318 = \DFF_51.Q ;
  assign g1320 = \DFF_111.Q ;
  assign g1321 = \DFF_51.Q ;
  assign g1322 = \DFF_191.D ;
  assign g1323 = \DFF_26.Q ;
  assign g1324 = \DFF_111.Q ;
  assign g1325 = \DFF_179.Q ;
  assign g1327 = \DFF_207.Q ;
  assign g1328 = \DFF_26.Q ;
  assign g1329 = \DFF_82.Q ;
  assign g1330 = \DFF_129.Q ;
  assign g1331 = \DFF_207.Q ;
  assign g1332 = \DFF_94.Q ;
  assign g1333 = \DFF_200.Q ;
  assign g1334 = \DFF_129.Q ;
  assign g1335 = \DFF_75.Q ;
  assign g1337 = \DFF_208.Q ;
  assign g1338 = \DFF_200.Q ;
  assign g1339 = \DFF_188.Q ;
  assign g1340 = \DFF_208.Q ;
  assign g1341 = \DFF_52.Q ;
  assign g1344 = \DFF_188.Q ;
  assign g1345 = \DFF_178.Q ;
  assign g1348 = \DFF_17.Q ;
  assign g1352 = \DFF_201.Q ;
  assign g1355 = \DFF_178.Q ;
  assign g1363 = \DFF_52.Q ;
  assign g1366 = \DFF_201.Q ;
  assign g1372 = \DFF_178.Q ;
  assign g1375 = \DFF_3.Q ;
  assign g1378 = \DFF_17.Q ;
  assign g1381 = \DFF_201.Q ;
  assign g1384 = \DFF_134.Q ;
  assign g1391 = \DFF_178.Q ;
  assign g1395 = \DFF_201.Q ;
  assign g14 = \DFF_128.Q ;
  assign g1450 = \DFF_188.Q ;
  assign g1461 = \DFF_188.Q ;
  assign g1472 = \DFF_69.D ;
  assign g1477 = \DFF_69.D ;
  assign g1480 = \DFF_139.Q ;
  assign g1498 = \DFF_80.D ;
  assign g15 = \DFF_63.Q ;
  assign g1503 = g639;
  assign g1504 = \DFF_168.Q ;
  assign g1513 = g639;
  assign g1519 = \DFF_43.Q ;
  assign g1528 = g639;
  assign g1533 = g639;
  assign g1539 = g639;
  assign g1542 = g639;
  assign g1549 = g639;
  assign g1556 = g639;
  assign g1559 = \DFF_153.D ;
  assign g1586 = \DFF_161.Q ;
  assign g1587 = \DFF_69.D ;
  assign g1593 = \DFF_190.Q ;
  assign g1594 = \DFF_153.D ;
  assign g1608 = \DFF_111.Q ;
  assign g1623 = \DFF_26.Q ;
  assign g1631 = \DFF_207.Q ;
  assign g1636 = \DFF_129.Q ;
  assign g1640 = \DFF_200.Q ;
  assign g1641 = \DFF_111.Q ;
  assign g1643 = \DFF_208.Q ;
  assign g1644 = \DFF_26.Q ;
  assign g1645 = \DFF_188.Q ;
  assign g1646 = \DFF_207.Q ;
  assign g1647 = \DFF_129.Q ;
  assign g1648 = \DFF_200.Q ;
  assign g1649 = \DFF_139.Q ;
  assign g1653 = \DFF_208.Q ;
  assign g1654 = g639;
  assign g1655 = \DFF_139.Q ;
  assign g1659 = \DFF_188.Q ;
  assign g1660 = \DFF_139.Q ;
  assign g1664 = \DFF_208.Q ;
  assign g1665 = \DFF_139.Q ;
  assign g1670 = \DFF_200.Q ;
  assign g1671 = \DFF_139.Q ;
  assign g1673 = \DFF_129.Q ;
  assign g1674 = \DFF_139.Q ;
  assign g1678 = \DFF_207.Q ;
  assign g1679 = \DFF_139.Q ;
  assign g1681 = \DFF_26.Q ;
  assign g1684 = \DFF_111.Q ;
  assign g1685 = \DFF_51.Q ;
  assign g1688 = \DFF_47.Q ;
  assign g1692 = \DFF_167.Q ;
  assign g1696 = \DFF_90.Q ;
  assign g1699 = \DFF_44.Q ;
  assign g1703 = \DFF_79.Q ;
  assign g1711 = \DFF_186.Q ;
  assign g1721 = \DFF_27.Q ;
  assign g1724 = \DFF_48.Q ;
  assign g1726 = \DFF_63.Q ;
  assign g1732 = \DFF_51.Q ;
  assign g1733 = \DFF_111.Q ;
  assign g1734 = \DFF_69.D ;
  assign g1735 = \DFF_187.Q ;
  assign g1739 = \DFF_26.Q ;
  assign g1747 = \DFF_207.Q ;
  assign g1748 = \DFF_51.Q ;
  assign g1759 = \DFF_129.Q ;
  assign g1760 = \DFF_111.Q ;
  assign g1761 = \DFF_51.Q ;
  assign g1762 = \DFF_51.Q ;
  assign g1771 = \DFF_200.Q ;
  assign g1772 = \DFF_26.Q ;
  assign g1773 = \DFF_111.Q ;
  assign g1774 = \DFF_111.Q ;
  assign g1775 = \DFF_69.D ;
  assign g1781 = \DFF_208.Q ;
  assign g1782 = \DFF_207.Q ;
  assign g1783 = \DFF_26.Q ;
  assign g1787 = \DFF_26.Q ;
  assign g1788 = \DFF_139.Q ;
  assign g1789 = \DFF_188.Q ;
  assign g1790 = \DFF_129.Q ;
  assign g1791 = \DFF_207.Q ;
  assign g1792 = \DFF_207.Q ;
  assign g18 = \DFF_6.Q ;
  assign g1802 = g2584;
  assign g1805 = \DFF_51.Q ;
  assign g1806 = \DFF_200.Q ;
  assign g1807 = \DFF_129.Q ;
  assign g1811 = \DFF_129.Q ;
  assign g1812 = \DFF_208.Q ;
  assign g1813 = \DFF_200.Q ;
  assign g1814 = \DFF_200.Q ;
  assign g1819 = \DFF_188.Q ;
  assign g1820 = \DFF_208.Q ;
  assign g1821 = \DFF_208.Q ;
  assign g1823 = \DFF_188.Q ;
  assign g1824 = \DFF_188.Q ;
  assign g1825 = \DFF_51.Q ;
  assign g1830 = g564;
  assign g1831 = \DFF_80.D ;
  assign g1832 = \DFF_188.Q ;
  assign g1833 = \DFF_207.Q ;
  assign g1834 = \DFF_208.Q ;
  assign g1835 = \DFF_26.Q ;
  assign g1836 = \DFF_111.Q ;
  assign g1837 = \DFF_51.Q ;
  assign g1841 = \DFF_188.Q ;
  assign g1846 = \DFF_208.Q ;
  assign g1848 = \DFF_69.D ;
  assign g1849 = \DFF_88.Q ;
  assign g1852 = \DFF_153.D ;
  assign g1854 = \DFF_189.Q ;
  assign g1858 = \DFF_189.Q ;
  assign g1875 = \DFF_168.Q ;
  assign g1884 = \DFF_88.Q ;
  assign g1891 = \DFF_168.Q ;
  assign g1894 = \DFF_43.Q ;
  assign g1899 = \DFF_189.Q ;
  assign g19 = \DFF_187.Q ;
  assign g1902 = \DFF_83.Q ;
  assign g1911 = \DFF_168.Q ;
  assign g1914 = \DFF_43.Q ;
  assign g1925 = \DFF_168.Q ;
  assign g1928 = \DFF_168.Q ;
  assign g1931 = \DFF_43.Q ;
  assign g1937 = \DFF_189.Q ;
  assign g1947 = \DFF_43.Q ;
  assign g1950 = \DFF_43.Q ;
  assign g1960 = \DFF_168.Q ;
  assign g1969 = \DFF_43.Q ;
  assign g197 = \DFF_179.Q ;
  assign g1979 = \DFF_168.Q ;
  assign g1988 = \DFF_43.Q ;
  assign g1998 = \DFF_168.Q ;
  assign g2 = \DFF_117.Q ;
  assign g2004 = \DFF_43.Q ;
  assign g204 = \DFF_168.Q ;
  assign g2040 = g705;
  assign g2041 = \DFF_191.D ;
  assign g2044 = \DFF_158.Q ;
  assign g205 = \DFF_178.Q ;
  assign g206 = \DFF_52.Q ;
  assign g207 = \DFF_3.Q ;
  assign g208 = \DFF_37.Q ;
  assign g2086 = \DFF_188.Q ;
  assign g2088 = \DFF_208.Q ;
  assign g209 = \DFF_146.Q ;
  assign g2090 = \DFF_188.Q ;
  assign g2096 = \DFF_200.Q ;
  assign g2097 = \DFF_208.Q ;
  assign g210 = \DFF_164.Q ;
  assign g2102 = \DFF_129.Q ;
  assign g2103 = \DFF_200.Q ;
  assign g2108 = \DFF_207.Q ;
  assign g2109 = \DFF_129.Q ;
  assign g211 = \DFF_87.Q ;
  assign g2117 = \DFF_26.Q ;
  assign g2118 = \DFF_207.Q ;
  assign g212 = \DFF_76.Q ;
  assign g2134 = \DFF_111.Q ;
  assign g2135 = \DFF_26.Q ;
  assign g2154 = \DFF_51.Q ;
  assign g2155 = \DFF_111.Q ;
  assign g2158 = \DFF_51.Q ;
  assign g2172 = \DFF_188.Q ;
  assign g2173 = \DFF_200.Q ;
  assign g2174 = \DFF_208.Q ;
  assign g2175 = \DFF_188.Q ;
  assign g2176 = \DFF_129.Q ;
  assign g2177 = \DFF_200.Q ;
  assign g2178 = \DFF_208.Q ;
  assign g2179 = g567;
  assign g218 = \DFF_156.Q ;
  assign g2194 = \DFF_207.Q ;
  assign g2195 = \DFF_129.Q ;
  assign g2196 = \DFF_200.Q ;
  assign g2197 = \DFF_19.Q ;
  assign g2212 = \DFF_26.Q ;
  assign g2213 = \DFF_207.Q ;
  assign g2214 = \DFF_129.Q ;
  assign g2215 = \DFF_58.Q ;
  assign g2230 = \DFF_111.Q ;
  assign g2231 = \DFF_26.Q ;
  assign g2232 = \DFF_207.Q ;
  assign g2233 = \DFF_200.Q ;
  assign g2234 = \DFF_141.Q ;
  assign g224 = \DFF_152.Q ;
  assign g2241 = \DFF_51.Q ;
  assign g2242 = \DFF_111.Q ;
  assign g2243 = \DFF_26.Q ;
  assign g2244 = \DFF_129.Q ;
  assign g2245 = \DFF_28.Q ;
  assign g2252 = \DFF_51.Q ;
  assign g2253 = \DFF_111.Q ;
  assign g2254 = \DFF_207.Q ;
  assign g2256 = \DFF_30.Q ;
  assign g2264 = \DFF_51.Q ;
  assign g2265 = \DFF_26.Q ;
  assign g2268 = \DFF_170.Q ;
  assign g2275 = \DFF_111.Q ;
  assign g2276 = \DFF_93.Q ;
  assign g2283 = \DFF_51.Q ;
  assign g2284 = \DFF_89.Q ;
  assign g2293 = \DFF_169.Q ;
  assign g2295 = \DFF_169.Q ;
  assign g230 = \DFF_166.Q ;
  assign g2308 = \DFF_188.Q ;
  assign g2312 = \DFF_188.Q ;
  assign g2315 = \DFF_48.Q ;
  assign g2316 = g2584;
  assign g2317 = \DFF_188.Q ;
  assign g2320 = \DFF_188.Q ;
  assign g2324 = \DFF_188.Q ;
  assign g2327 = \DFF_188.Q ;
  assign g2333 = \DFF_188.Q ;
  assign g2343 = \DFF_188.Q ;
  assign g2347 = \DFF_188.Q ;
  assign g2357 = \DFF_188.Q ;
  assign g236 = \DFF_176.Q ;
  assign g2361 = \DFF_188.Q ;
  assign g2370 = \DFF_208.Q ;
  assign g2378 = \DFF_188.Q ;
  assign g2390 = \DFF_190.Q ;
  assign g2397 = \DFF_200.Q ;
  assign g24 = \DFF_10.Q ;
  assign g2405 = \DFF_188.Q ;
  assign g2408 = \DFF_161.Q ;
  assign g242 = \DFF_157.Q ;
  assign g2422 = \DFF_129.Q ;
  assign g2430 = \DFF_188.Q ;
  assign g2433 = g4809;
  assign g2436 = \DFF_188.Q ;
  assign g2449 = \DFF_207.Q ;
  assign g2457 = \DFF_188.Q ;
  assign g2460 = \DFF_208.Q ;
  assign g2473 = \DFF_26.Q ;
  assign g248 = \DFF_116.Q ;
  assign g2481 = \DFF_188.Q ;
  assign g2484 = \DFF_200.Q ;
  assign g2497 = \DFF_111.Q ;
  assign g25 = \DFF_167.Q ;
  assign g2505 = \DFF_129.Q ;
  assign g2518 = \DFF_51.Q ;
  assign g2524 = \DFF_207.Q ;
  assign g254 = \DFF_114.Q ;
  assign g2544 = \DFF_47.Q ;
  assign g2550 = \DFF_188.Q ;
  assign g2554 = \DFF_26.Q ;
  assign g2574 = \DFF_208.Q ;
  assign g2575 = \DFF_111.Q ;
  assign g2576 = \DFF_200.Q ;
  assign g2580 = \DFF_51.Q ;
  assign g2581 = \DFF_129.Q ;
  assign g2586 = \DFF_69.D ;
  assign g2587 = \DFF_153.D ;
  assign g2588 = \DFF_51.Q ;
  assign g2591 = \DFF_111.Q ;
  assign g2594 = \DFF_51.Q ;
  assign g2599 = \DFF_188.Q ;
  assign g260 = \DFF_183.Q ;
  assign g2604 = \DFF_208.Q ;
  assign g2609 = \DFF_200.Q ;
  assign g2612 = \DFF_158.Q ;
  assign g2618 = \DFF_191.D ;
  assign g2619 = \DFF_129.Q ;
  assign g2622 = \DFF_158.Q ;
  assign g2631 = \DFF_207.Q ;
  assign g2634 = \DFF_158.Q ;
  assign g2644 = \DFF_26.Q ;
  assign g2647 = \DFF_158.Q ;
  assign g2650 = \DFF_158.Q ;
  assign g266 = \DFF_197.Q ;
  assign g2660 = \DFF_111.Q ;
  assign g2663 = \DFF_69.D ;
  assign g2670 = \DFF_144.D ;
  assign g2672 = \DFF_51.Q ;
  assign g2675 = \DFF_158.Q ;
  assign g2678 = \DFF_69.D ;
  assign g2686 = g567;
  assign g2688 = \DFF_188.Q ;
  assign g269 = \DFF_82.Q ;
  assign g2691 = \DFF_69.D ;
  assign g2701 = \DFF_188.Q ;
  assign g2705 = \DFF_19.Q ;
  assign g2706 = \DFF_208.Q ;
  assign g2709 = \DFF_158.Q ;
  assign g2712 = \DFF_69.D ;
  assign g2722 = \DFF_208.Q ;
  assign g2726 = \DFF_58.Q ;
  assign g2727 = \DFF_69.D ;
  assign g2734 = \DFF_200.Q ;
  assign g2738 = \DFF_69.D ;
  assign g2739 = \DFF_141.Q ;
  assign g2740 = \DFF_158.Q ;
  assign g2743 = \DFF_69.D ;
  assign g2744 = \DFF_169.Q ;
  assign g2748 = \DFF_129.Q ;
  assign g2752 = \DFF_69.D ;
  assign g2753 = \DFF_28.Q ;
  assign g2754 = \DFF_69.D ;
  assign g2755 = \DFF_169.Q ;
  assign g2756 = \DFF_169.Q ;
  assign g276 = \DFF_43.Q ;
  assign g2760 = \DFF_207.Q ;
  assign g2764 = \DFF_69.D ;
  assign g2765 = \DFF_30.Q ;
  assign g2766 = \DFF_69.D ;
  assign g2767 = \DFF_169.Q ;
  assign g2768 = \DFF_169.Q ;
  assign g277 = \DFF_201.Q ;
  assign g2772 = \DFF_26.Q ;
  assign g2776 = \DFF_69.D ;
  assign g2777 = \DFF_170.Q ;
  assign g2778 = \DFF_169.Q ;
  assign g2779 = \DFF_169.Q ;
  assign g278 = \DFF_17.Q ;
  assign g2783 = \DFF_111.Q ;
  assign g2787 = \DFF_69.D ;
  assign g2788 = \DFF_93.Q ;
  assign g2789 = \DFF_169.Q ;
  assign g279 = \DFF_134.Q ;
  assign g2790 = \DFF_169.Q ;
  assign g2792 = \DFF_169.Q ;
  assign g2796 = \DFF_51.Q ;
  assign g28 = \DFF_123.Q ;
  assign g280 = \DFF_142.Q ;
  assign g2800 = \DFF_69.D ;
  assign g2801 = \DFF_89.Q ;
  assign g2802 = \DFF_169.Q ;
  assign g2803 = \DFF_169.Q ;
  assign g2805 = \DFF_169.Q ;
  assign g2806 = \DFF_169.Q ;
  assign g2809 = \DFF_188.Q ;
  assign g281 = \DFF_61.Q ;
  assign g2813 = \DFF_69.D ;
  assign g2814 = \DFF_48.Q ;
  assign g2817 = \DFF_169.Q ;
  assign g2818 = \DFF_169.Q ;
  assign g2819 = \DFF_169.Q ;
  assign g282 = \DFF_50.Q ;
  assign g2820 = \DFF_169.Q ;
  assign g2822 = \DFF_208.Q ;
  assign g2826 = \DFF_69.D ;
  assign g2827 = \DFF_169.Q ;
  assign g2828 = \DFF_169.Q ;
  assign g2829 = \DFF_169.Q ;
  assign g283 = \DFF_125.Q ;
  assign g2830 = \DFF_169.Q ;
  assign g2835 = \DFF_169.Q ;
  assign g2836 = \DFF_169.Q ;
  assign g2837 = \DFF_169.Q ;
  assign g2838 = \DFF_169.Q ;
  assign g2839 = \DFF_169.Q ;
  assign g284 = \DFF_76.Q ;
  assign g2840 = \DFF_169.Q ;
  assign g2841 = \DFF_169.Q ;
  assign g2845 = \DFF_169.Q ;
  assign g285 = \DFF_156.Q ;
  assign g2859 = \DFF_19.D ;
  assign g286 = \DFF_152.Q ;
  assign g2861 = \DFF_140.D ;
  assign g2864 = \DFF_169.Q ;
  assign g2866 = \DFF_169.Q ;
  assign g2867 = \DFF_169.Q ;
  assign g287 = \DFF_166.Q ;
  assign g2871 = \DFF_169.Q ;
  assign g2872 = \DFF_169.Q ;
  assign g2875 = \DFF_169.Q ;
  assign g2876 = \DFF_169.Q ;
  assign g288 = \DFF_176.Q ;
  assign g2883 = \DFF_169.Q ;
  assign g2884 = \DFF_169.Q ;
  assign g2885 = \DFF_169.Q ;
  assign g2886 = \DFF_169.Q ;
  assign g2888 = \DFF_169.Q ;
  assign g2889 = \DFF_169.Q ;
  assign g289 = \DFF_157.Q ;
  assign g2892 = \DFF_169.Q ;
  assign g2893 = \DFF_169.Q ;
  assign g29 = \DFF_90.Q ;
  assign g290 = \DFF_116.Q ;
  assign g2904 = \DFF_169.Q ;
  assign g2905 = \DFF_169.Q ;
  assign g291 = \DFF_114.Q ;
  assign g2912 = \DFF_169.Q ;
  assign g292 = \DFF_183.Q ;
  assign g293 = \DFF_94.Q ;
  assign g2945 = g705;
  assign g2967 = \DFF_190.Q ;
  assign g297 = \DFF_75.Q ;
  assign g2974 = \DFF_161.Q ;
  assign g2975 = \DFF_170.Q ;
  assign g2998 = \DFF_200.Q ;
  assign g3 = \DFF_44.Q ;
  assign g3001 = \DFF_93.Q ;
  assign g3016 = \DFF_129.Q ;
  assign g3022 = \DFF_89.Q ;
  assign g3031 = \DFF_207.Q ;
  assign g3040 = g567;
  assign g3043 = \DFF_26.Q ;
  assign g3052 = \DFF_19.Q ;
  assign g3054 = \DFF_111.Q ;
  assign g3063 = \DFF_58.Q ;
  assign g3064 = \DFF_51.Q ;
  assign g3073 = \DFF_141.Q ;
  assign g3082 = \DFF_28.Q ;
  assign g3093 = \DFF_30.Q ;
  assign g3104 = \DFF_200.Q ;
  assign g3118 = \DFF_129.Q ;
  assign g3128 = \DFF_207.Q ;
  assign g3136 = \DFF_26.Q ;
  assign g3150 = \DFF_111.Q ;
  assign g3158 = \DFF_188.Q ;
  assign g3162 = \DFF_51.Q ;
  assign g3173 = \DFF_208.Q ;
  assign g3177 = \DFF_188.Q ;
  assign g3183 = \DFF_200.Q ;
  assign g3187 = \DFF_208.Q ;
  assign g3192 = \DFF_129.Q ;
  assign g3196 = \DFF_200.Q ;
  assign g3200 = \DFF_207.Q ;
  assign g3204 = \DFF_129.Q ;
  assign g3209 = \DFF_26.Q ;
  assign g3212 = \DFF_207.Q ;
  assign g3216 = \DFF_111.Q ;
  assign g3219 = \DFF_26.Q ;
  assign g3222 = g705;
  assign g3224 = g567;
  assign g3225 = \DFF_19.Q ;
  assign g3226 = \DFF_58.Q ;
  assign g3227 = \DFF_141.Q ;
  assign g3228 = \DFF_28.Q ;
  assign g3229 = \DFF_30.Q ;
  assign g3230 = \DFF_170.Q ;
  assign g3231 = \DFF_93.Q ;
  assign g3232 = \DFF_89.Q ;
  assign g3233 = g567;
  assign g3234 = \DFF_19.Q ;
  assign g3235 = \DFF_58.Q ;
  assign g3236 = \DFF_141.Q ;
  assign g3237 = \DFF_28.Q ;
  assign g3238 = \DFF_30.Q ;
  assign g3239 = \DFF_170.Q ;
  assign g3240 = \DFF_93.Q ;
  assign g3241 = \DFF_89.Q ;
  assign g3242 = \DFF_128.Q ;
  assign g3247 = \DFF_6.Q ;
  assign g3259 = \DFF_10.Q ;
  assign g3263 = \DFF_123.Q ;
  assign g3267 = g32;
  assign g3271 = g36;
  assign g3284 = \DFF_179.Q ;
  assign g3289 = \DFF_179.Q ;
  assign g3291 = \DFF_82.Q ;
  assign g3297 = \DFF_179.Q ;
  assign g3299 = \DFF_82.Q ;
  assign g33 = \DFF_79.Q ;
  assign g3306 = \DFF_179.Q ;
  assign g3308 = \DFF_82.Q ;
  assign g3320 = \DFF_179.Q ;
  assign g3322 = \DFF_82.Q ;
  assign g3331 = \DFF_179.Q ;
  assign g3332 = \DFF_82.Q ;
  assign g3342 = \DFF_179.Q ;
  assign g3343 = \DFF_82.Q ;
  assign g3354 = \DFF_179.Q ;
  assign g3355 = \DFF_82.Q ;
  assign g3363 = \DFF_179.Q ;
  assign g3364 = \DFF_82.Q ;
  assign g3370 = \DFF_82.Q ;
  assign g3440 = \DFF_144.D ;
  assign g3451 = \DFF_179.Q ;
  assign g3452 = \DFF_179.Q ;
  assign g3453 = \DFF_82.Q ;
  assign g3454 = \DFF_58.D ;
  assign g3455 = \DFF_179.Q ;
  assign g3456 = \DFF_82.Q ;
  assign g3457 = \DFF_179.Q ;
  assign g3458 = \DFF_82.Q ;
  assign g3459 = \DFF_179.Q ;
  assign g3460 = \DFF_82.Q ;
  assign g3462 = \DFF_179.Q ;
  assign g3463 = \DFF_82.Q ;
  assign g3477 = \DFF_179.Q ;
  assign g3478 = \DFF_82.Q ;
  assign g3482 = \DFF_179.Q ;
  assign g3483 = \DFF_82.Q ;
  assign g3486 = g4809;
  assign g3488 = \DFF_82.Q ;
  assign g3491 = g41;
  assign g3527 = \DFF_51.Q ;
  assign g3534 = \DFF_19.D ;
  assign g3537 = \DFF_140.D ;
  assign g3541 = \DFF_23.Q ;
  assign g3545 = g44;
  assign g3546 = g45;
  assign g3557 = g23;
  assign g3559 = g22;
  assign g3564 = g47;
  assign g3567 = g37;
  assign g3571 = g38;
  assign g3589 = g39;
  assign g3593 = g40;
  assign g3599 = g4121;
  assign g3600 = \DFF_48.Q ;
  assign g3601 = \DFF_48.Q ;
  assign g3604 = \DFF_190.Q ;
  assign g3612 = \DFF_161.Q ;
  assign g3638 = g46;
  assign g3673 = g42;
  assign g3705 = \DFF_209.Q ;
  assign g3710 = \DFF_117.Q ;
  assign g3714 = \DFF_98.Q ;
  assign g3719 = \DFF_127.Q ;
  assign g3766 = g42;
  assign g3768 = \DFF_154.D ;
  assign g3771 = g42;
  assign g3783 = g45;
  assign g3787 = g46;
  assign g3803 = \DFF_161.Q ;
  assign g3807 = \DFF_190.Q ;
  assign g3814 = \DFF_169.D ;
  assign g3828 = \DFF_126.D ;
  assign g3832 = \DFF_123.Q ;
  assign g3834 = g32;
  assign g3835 = \DFF_128.Q ;
  assign g3836 = \DFF_51.Q ;
  assign g3838 = \DFF_209.Q ;
  assign g3839 = g36;
  assign g3840 = \DFF_6.Q ;
  assign g3844 = \DFF_141.D ;
  assign g3846 = \DFF_117.Q ;
  assign g3847 = g37;
  assign g3848 = \DFF_10.Q ;
  assign g3852 = \DFF_98.Q ;
  assign g3853 = g38;
  assign g3854 = \DFF_123.Q ;
  assign g3859 = \DFF_127.Q ;
  assign g3860 = g39;
  assign g3861 = g40;
  assign g3866 = \DFF_128.Q ;
  assign g3867 = \DFF_209.Q ;
  assign g3874 = \DFF_144.D ;
  assign g3875 = \DFF_6.Q ;
  assign g3876 = \DFF_117.Q ;
  assign g3881 = \DFF_10.Q ;
  assign g3882 = \DFF_98.Q ;
  assign g3885 = \DFF_127.Q ;
  assign g3910 = \DFF_197.D ;
  assign g3922 = \DFF_58.D ;
  assign g3932 = g40;
  assign g3940 = g32;
  assign g3952 = g36;
  assign g3960 = \DFF_19.D ;
  assign g3962 = g37;
  assign g3963 = g42;
  assign g3967 = \DFF_140.D ;
  assign g3969 = g38;
  assign g3970 = g44;
  assign g3975 = g39;
  assign g3976 = g45;
  assign g3980 = g46;
  assign g3984 = \DFF_191.D ;
  assign g4014 = g23;
  assign g4016 = g22;
  assign g402 = \DFF_74.Q ;
  assign g4034 = g41;
  assign g4036 = g47;
  assign g4040 = g4121;
  assign g406 = \DFF_175.Q ;
  assign g4098 = g23;
  assign g4099 = g32;
  assign g410 = \DFF_77.Q ;
  assign g4100 = g36;
  assign g4101 = g37;
  assign g4102 = g38;
  assign g4103 = g39;
  assign g4104 = g22;
  assign g4105 = g40;
  assign g4106 = g42;
  assign g4107 = g44;
  assign g4108 = g45;
  assign g4109 = g46;
  assign g4110 = g41;
  assign g4112 = g47;
  assign g4122 = \DFF_19.D ;
  assign g4123 = \DFF_140.D ;
  assign g4124 = \DFF_144.D ;
  assign g4125 = g42;
  assign g4126 = g42;
  assign g4127 = g45;
  assign g4128 = g46;
  assign g4129 = \DFF_209.Q ;
  assign g4130 = \DFF_117.Q ;
  assign g4131 = \DFF_98.Q ;
  assign g4132 = \DFF_127.Q ;
  assign g4133 = \DFF_128.Q ;
  assign g4134 = \DFF_6.Q ;
  assign g4135 = \DFF_10.Q ;
  assign g4136 = \DFF_123.Q ;
  assign g4137 = g32;
  assign g4138 = g36;
  assign g4139 = g37;
  assign g414 = \DFF_195.Q ;
  assign g4140 = g38;
  assign g4141 = g39;
  assign g4142 = \DFF_209.Q ;
  assign g4143 = \DFF_117.Q ;
  assign g4144 = \DFF_98.Q ;
  assign g4145 = \DFF_127.Q ;
  assign g4146 = \DFF_128.Q ;
  assign g4147 = \DFF_6.Q ;
  assign g4148 = \DFF_10.Q ;
  assign g4149 = \DFF_123.Q ;
  assign g4150 = g40;
  assign g4152 = \DFF_191.D ;
  assign g4153 = \DFF_169.D ;
  assign g4157 = \DFF_36.D ;
  assign g418 = \DFF_73.Q ;
  assign g4194 = \DFF_197.D ;
  assign g4213 = \DFF_154.D ;
  assign g4219 = \DFF_28.D ;
  assign g422 = \DFF_163.Q ;
  assign g4228 = \DFF_126.D ;
  assign g4249 = \DFF_141.D ;
  assign g426 = \DFF_57.Q ;
  assign g4299 = \DFF_58.D ;
  assign g43 = \DFF_48.Q ;
  assign g430 = \DFF_78.Q ;
  assign g4307 = \DFF_190.Q ;
  assign g4308 = \DFF_190.Q ;
  assign g4320 = g4809;
  assign g4321 = \DFF_161.Q ;
  assign g4322 = \DFF_161.Q ;
  assign g434 = \DFF_196.Q ;
  assign g4343 = g4809;
  assign g4350 = \DFF_48.Q ;
  assign g437 = \DFF_42.Q ;
  assign g441 = \DFF_84.Q ;
  assign g4422 = g564;
  assign g4423 = \DFF_126.D ;
  assign g4424 = \DFF_58.D ;
  assign g4425 = \DFF_169.D ;
  assign g4426 = \DFF_191.D ;
  assign g4430 = \DFF_84.D ;
  assign g4433 = \DFF_42.D ;
  assign g4434 = \DFF_78.D ;
  assign g4436 = \DFF_196.D ;
  assign g4438 = \DFF_74.D ;
  assign g4440 = \DFF_5.D ;
  assign g4441 = \DFF_175.D ;
  assign g4443 = \DFF_68.D ;
  assign g4444 = \DFF_77.D ;
  assign g4446 = \DFF_81.D ;
  assign g4447 = \DFF_195.D ;
  assign g445 = \DFF_96.Q ;
  assign g4450 = \DFF_53.D ;
  assign g4451 = \DFF_73.D ;
  assign g4454 = \DFF_96.D ;
  assign g4455 = \DFF_163.D ;
  assign g4458 = \DFF_57.D ;
  assign g4460 = \DFF_15.D ;
  assign g449 = \DFF_53.Q ;
  assign g4492 = \DFF_36.D ;
  assign g4501 = \DFF_30.D ;
  assign g4514 = \DFF_197.D ;
  assign g4519 = \DFF_154.D ;
  assign g453 = \DFF_81.Q ;
  assign g4562 = \DFF_28.D ;
  assign g457 = \DFF_68.Q ;
  assign g4603 = g4809;
  assign g4609 = \DFF_141.D ;
  assign g461 = \DFF_5.Q ;
  assign g4644 = \DFF_48.Q ;
  assign g465 = \DFF_11.Q ;
  assign g4657 = \DFF_154.D ;
  assign g4658 = \DFF_141.D ;
  assign g4659 = \DFF_197.D ;
  assign g4687 = \DFF_40.D ;
  assign g4692 = \DFF_84.D ;
  assign g4699 = \DFF_42.D ;
  assign g4700 = \DFF_78.D ;
  assign g4702 = \DFF_196.D ;
  assign g4703 = \DFF_74.D ;
  assign g4704 = \DFF_5.D ;
  assign g4705 = \DFF_175.D ;
  assign g4706 = \DFF_68.D ;
  assign g4707 = \DFF_77.D ;
  assign g471 = \DFF_70.Q ;
  assign g4711 = \DFF_81.D ;
  assign g4712 = \DFF_195.D ;
  assign g4714 = \DFF_53.D ;
  assign g4715 = \DFF_73.D ;
  assign g4718 = \DFF_96.D ;
  assign g4719 = \DFF_163.D ;
  assign g4721 = \DFF_57.D ;
  assign g4758 = \DFF_15.D ;
  assign g4761 = \DFF_170.D ;
  assign g4765 = \DFF_36.D ;
  assign g478 = \DFF_148.Q ;
  assign g4781 = \DFF_30.D ;
  assign g4798 = \DFF_28.D ;
  assign g48 = \DFF_23.Q ;
  assign g4810 = g4809;
  assign g4822 = \DFF_190.Q ;
  assign g4823 = \DFF_48.Q ;
  assign g4824 = \DFF_161.Q ;
  assign g4841 = \DFF_5.D ;
  assign g4842 = \DFF_68.D ;
  assign g4843 = \DFF_81.D ;
  assign g4844 = \DFF_53.D ;
  assign g4845 = \DFF_96.D ;
  assign g4846 = \DFF_84.D ;
  assign g4847 = \DFF_42.D ;
  assign g4848 = \DFF_196.D ;
  assign g4849 = \DFF_74.D ;
  assign g485 = \DFF_190.Q ;
  assign g4850 = \DFF_175.D ;
  assign g4851 = \DFF_77.D ;
  assign g4852 = \DFF_195.D ;
  assign g4853 = \DFF_73.D ;
  assign g4854 = \DFF_163.D ;
  assign g4855 = \DFF_57.D ;
  assign g4856 = \DFF_78.D ;
  assign g4857 = \DFF_28.D ;
  assign g4858 = \DFF_36.D ;
  assign g486 = \DFF_69.Q ;
  assign g4871 = \DFF_48.Q ;
  assign g4872 = \DFF_121.D ;
  assign g489 = \DFF_153.Q ;
  assign g492 = \DFF_135.Q ;
  assign g496 = \DFF_21.Q ;
  assign g500 = \DFF_177.Q ;
  assign g5010 = \DFF_40.D ;
  assign g5017 = \DFF_93.D ;
  assign g5019 = \DFF_14.D ;
  assign g504 = \DFF_102.Q ;
  assign g5051 = \DFF_15.D ;
  assign g508 = \DFF_172.Q ;
  assign g5089 = \DFF_170.D ;
  assign g5110 = \DFF_30.D ;
  assign g512 = \DFF_204.Q ;
  assign g5135 = \DFF_190.Q ;
  assign g5136 = \DFF_161.Q ;
  assign g5137 = \DFF_48.Q ;
  assign g5147 = \DFF_15.D ;
  assign g5148 = \DFF_30.D ;
  assign g5149 = \DFF_89.D ;
  assign g5151 = \DFF_14.D ;
  assign g516 = \DFF_109.Q ;
  assign g5167 = \DFF_64.D ;
  assign g520 = \DFF_60.Q ;
  assign g5219 = \DFF_121.D ;
  assign g5230 = \DFF_40.D ;
  assign g5231 = \DFF_131.D ;
  assign g524 = \DFF_182.Q ;
  assign g5273 = \DFF_93.D ;
  assign g528 = \DFF_55.Q ;
  assign g5307 = \DFF_170.D ;
  assign g5314 = \DFF_190.Q ;
  assign g5315 = g4809;
  assign g5316 = \DFF_161.Q ;
  assign g532 = \DFF_205.Q ;
  assign g5328 = \DFF_40.D ;
  assign g5329 = \DFF_170.D ;
  assign g5330 = \DFF_14.D ;
  assign g5355 = \DFF_190.Q ;
  assign g5358 = \DFF_161.Q ;
  assign g536 = \DFF_110.Q ;
  assign g5375 = \DFF_89.D ;
  assign g5383 = \DFF_64.D ;
  assign g5385 = g6282;
  assign g5386 = \DFF_59.D ;
  assign g5387 = \DFF_121.D ;
  assign g541 = \DFF_105.Q ;
  assign g5432 = \DFF_93.D ;
  assign g545 = \DFF_113.Q ;
  assign g5466 = \DFF_131.D ;
  assign g5468 = \DFF_190.Q ;
  assign g5469 = \DFF_161.Q ;
  assign g548 = \DFF_173.Q ;
  assign g5489 = \DFF_121.D ;
  assign g5490 = \DFF_93.D ;
  assign g5491 = \DFF_131.D ;
  assign g551 = \DFF_25.Q ;
  assign g5531 = \DFF_168.D ;
  assign g5532 = \DFF_43.D ;
  assign g5533 = \DFF_37.D ;
  assign g5534 = \DFF_89.D ;
  assign g5535 = \DFF_142.D ;
  assign g554 = \DFF_20.Q ;
  assign g5540 = \DFF_64.D ;
  assign g5579 = \DFF_59.D ;
  assign g5580 = \DFF_89.D ;
  assign g5581 = \DFF_64.D ;
  assign g5582 = \DFF_59.D ;
  assign g5584 = \DFF_168.D ;
  assign g5587 = \DFF_43.D ;
  assign g5590 = \DFF_37.D ;
  assign g5593 = \DFF_142.D ;
  assign g5622 = \DFF_178.D ;
  assign g5624 = \DFF_52.D ;
  assign g5625 = \DFF_201.D ;
  assign g5626 = \DFF_3.D ;
  assign g5627 = \DFF_17.D ;
  assign g5628 = \DFF_134.D ;
  assign g5629 = \DFF_146.D ;
  assign g5630 = \DFF_61.D ;
  assign g5645 = g6282;
  assign g5692 = 1'b0;
  assign g5702 = \DFF_178.D ;
  assign g5705 = \DFF_52.D ;
  assign g5708 = \DFF_201.D ;
  assign g571 = \DFF_89.Q ;
  assign g5711 = \DFF_3.D ;
  assign g5714 = \DFF_17.D ;
  assign g5717 = \DFF_134.D ;
  assign g5720 = \DFF_146.D ;
  assign g5723 = \DFF_61.D ;
  assign g574 = \DFF_83.Q ;
  assign g5751 = \DFF_168.D ;
  assign g5752 = \DFF_43.D ;
  assign g5773 = \DFF_37.D ;
  assign g5774 = \DFF_142.D ;
  assign g578 = \DFF_158.Q ;
  assign g582 = \DFF_189.Q ;
  assign g586 = \DFF_88.Q ;
  assign g5875 = \DFF_168.D ;
  assign g5876 = \DFF_37.D ;
  assign g5877 = \DFF_43.D ;
  assign g5878 = \DFF_142.D ;
  assign g5879 = g6282;
  assign g590 = \DFF_24.Q ;
  assign g5917 = \DFF_178.D ;
  assign g5918 = \DFF_52.D ;
  assign g5919 = \DFF_201.D ;
  assign g5920 = \DFF_3.D ;
  assign g5921 = \DFF_17.D ;
  assign g5922 = \DFF_134.D ;
  assign g5923 = \DFF_146.D ;
  assign g5924 = \DFF_61.D ;
  assign g594 = \DFF_151.Q ;
  assign g598 = \DFF_19.Q ;
  assign g6 = \DFF_98.Q ;
  assign g602 = \DFF_140.Q ;
  assign g6032 = g6282;
  assign g606 = \DFF_28.Q ;
  assign g610 = \DFF_144.Q ;
  assign g6100 = \DFF_178.D ;
  assign g6101 = \DFF_52.D ;
  assign g6102 = \DFF_3.D ;
  assign g6103 = \DFF_146.D ;
  assign g6104 = \DFF_201.D ;
  assign g6105 = \DFF_17.D ;
  assign g6106 = \DFF_134.D ;
  assign g6107 = \DFF_61.D ;
  assign g6110 = g6284;
  assign g613 = \DFF_126.Q ;
  assign g6137 = g6282;
  assign g6142 = \DFF_48.D ;
  assign g616 = \DFF_154.Q ;
  assign g6167 = g6364;
  assign g6170 = g6368;
  assign g6173 = g6370;
  assign g6176 = g6372;
  assign g6179 = g6374;
  assign g6182 = g6360;
  assign g6185 = g6362;
  assign g6189 = g6366;
  assign g619 = \DFF_36.Q ;
  assign g622 = \DFF_15.Q ;
  assign g625 = \DFF_40.Q ;
  assign g628 = \DFF_121.Q ;
  assign g6283 = g6282;
  assign g6285 = g6284;
  assign g6286 = \DFF_55.D ;
  assign g6287 = \DFF_179.D ;
  assign g6289 = \DFF_105.D ;
  assign g6290 = \DFF_82.D ;
  assign g6291 = \DFF_158.D ;
  assign g6292 = \DFF_177.D ;
  assign g6293 = \DFF_110.D ;
  assign g6294 = \DFF_94.D ;
  assign g6295 = \DFF_189.D ;
  assign g6296 = \DFF_102.D ;
  assign g6297 = \DFF_11.D ;
  assign g6298 = \DFF_75.D ;
  assign g6299 = \DFF_88.D ;
  assign g6300 = \DFF_172.D ;
  assign g6301 = \DFF_205.D ;
  assign g6303 = \DFF_204.D ;
  assign g6304 = \DFF_151.D ;
  assign g6307 = \DFF_109.D ;
  assign g6309 = \DFF_60.D ;
  assign g631 = \DFF_64.Q ;
  assign g6310 = \DFF_182.D ;
  assign g6312 = \DFF_48.D ;
  assign g634 = \DFF_58.Q ;
  assign g6361 = g6360;
  assign g6363 = g6362;
  assign g6365 = g6364;
  assign g6367 = g6366;
  assign g6369 = g6368;
  assign g6371 = g6370;
  assign g6373 = g6372;
  assign g6375 = g6374;
  assign g638 = \DFF_139.Q ;
  assign g6407 = \DFF_48.D ;
  assign g6410 = \DFF_179.D ;
  assign g6411 = \DFF_55.D ;
  assign g6412 = \DFF_82.D ;
  assign g6413 = \DFF_105.D ;
  assign g6414 = \DFF_94.D ;
  assign g6415 = \DFF_177.D ;
  assign g6416 = \DFF_110.D ;
  assign g6417 = \DFF_75.D ;
  assign g6418 = \DFF_102.D ;
  assign g6419 = \DFF_11.D ;
  assign g642 = \DFF_141.Q ;
  assign g6420 = \DFF_172.D ;
  assign g6421 = \DFF_205.D ;
  assign g6422 = \DFF_204.D ;
  assign g6423 = \DFF_109.D ;
  assign g6424 = \DFF_60.D ;
  assign g6425 = \DFF_182.D ;
  assign g6426 = \DFF_83.D ;
  assign g6428 = \DFF_158.D ;
  assign g6431 = \DFF_189.D ;
  assign g6434 = \DFF_88.D ;
  assign g6437 = \DFF_24.D ;
  assign g6441 = \DFF_151.D ;
  assign g646 = \DFF_30.Q ;
  assign g6479 = \DFF_44.D ;
  assign g6480 = \DFF_186.D ;
  assign g6481 = \DFF_27.D ;
  assign g6482 = \DFF_63.D ;
  assign g6483 = \DFF_187.D ;
  assign g6485 = \DFF_167.D ;
  assign g6497 = \DFF_177.D ;
  assign g6498 = \DFF_102.D ;
  assign g6499 = \DFF_172.D ;
  assign g650 = \DFF_170.Q ;
  assign g6500 = \DFF_204.D ;
  assign g6501 = \DFF_109.D ;
  assign g6502 = \DFF_60.D ;
  assign g6503 = \DFF_182.D ;
  assign g6504 = \DFF_55.D ;
  assign g6505 = \DFF_105.D ;
  assign g6506 = \DFF_110.D ;
  assign g6507 = \DFF_11.D ;
  assign g6508 = \DFF_205.D ;
  assign g6509 = \DFF_179.D ;
  assign g6510 = \DFF_82.D ;
  assign g6511 = \DFF_94.D ;
  assign g6512 = \DFF_75.D ;
  assign g6515 = g6282;
  assign g6516 = g6284;
  assign g6519 = \DFF_167.D ;
  assign g6521 = \DFF_63.D ;
  assign g6523 = \DFF_44.D ;
  assign g6524 = \DFF_83.D ;
  assign g6525 = \DFF_186.D ;
  assign g6526 = \DFF_158.D ;
  assign g6527 = \DFF_27.D ;
  assign g6528 = \DFF_189.D ;
  assign g6529 = \DFF_88.D ;
  assign g6530 = \DFF_187.D ;
  assign g6531 = \DFF_24.D ;
  assign g6532 = \DFF_151.D ;
  assign g654 = \DFF_93.Q ;
  assign g6574 = g6360;
  assign g6575 = g6362;
  assign g6576 = g6364;
  assign g6577 = g6366;
  assign g6578 = g6368;
  assign g6579 = g6370;
  assign g658 = \DFF_169.Q ;
  assign g6580 = g6372;
  assign g6581 = g6374;
  assign g6591 = \DFF_83.D ;
  assign g6592 = \DFF_158.D ;
  assign g6593 = \DFF_189.D ;
  assign g6594 = \DFF_88.D ;
  assign g6595 = \DFF_24.D ;
  assign g6596 = \DFF_151.D ;
  assign g6597 = \DFF_44.D ;
  assign g6598 = \DFF_186.D ;
  assign g6599 = \DFF_27.D ;
  assign g6600 = \DFF_187.D ;
  assign g6601 = \DFF_167.D ;
  assign g6602 = \DFF_63.D ;
  assign g662 = \DFF_80.Q ;
  assign g663 = \DFF_143.Q ;
  assign g664 = \DFF_148.Q ;
  assign g665 = \DFF_143.Q ;
  assign g6658 = \DFF_23.D ;
  assign g666 = \DFF_180.Q ;
  assign g667 = \DFF_132.Q ;
  assign g668 = \DFF_161.Q ;
  assign g6684 = \DFF_6.D ;
  assign g6685 = \DFF_10.D ;
  assign g6686 = \DFF_209.D ;
  assign g6687 = \DFF_123.D ;
  assign g6688 = \DFF_117.D ;
  assign g6689 = \DFF_98.D ;
  assign g669 = \DFF_59.Q ;
  assign g6690 = \DFF_127.D ;
  assign g6691 = \DFF_128.D ;
  assign g6694 = \DFF_6.D ;
  assign g6695 = \DFF_10.D ;
  assign g6696 = \DFF_209.D ;
  assign g6697 = \DFF_123.D ;
  assign g6698 = \DFF_117.D ;
  assign g6699 = \DFF_98.D ;
  assign g6700 = \DFF_127.D ;
  assign g6701 = \DFF_128.D ;
  assign g6702 = \DFF_21.D ;
  assign g6704 = \DFF_135.D ;
  assign g6711 = \DFF_23.D ;
  assign g672 = \DFF_131.Q ;
  assign g6720 = \DFF_209.D ;
  assign g6721 = \DFF_117.D ;
  assign g6722 = \DFF_98.D ;
  assign g6723 = \DFF_127.D ;
  assign g6724 = \DFF_128.D ;
  assign g6725 = \DFF_6.D ;
  assign g6726 = \DFF_10.D ;
  assign g6727 = \DFF_123.D ;
  assign g6728 = 1'b0;
  assign g6729 = \DFF_23.D ;
  assign g6730 = \DFF_135.D ;
  assign g6743 = \DFF_21.D ;
  assign g6744 = \DFF_135.D ;
  assign g6745 = \DFF_21.D ;
  assign g675 = \DFF_147.Q ;
  assign g676 = \DFF_14.Q ;
  assign g677 = \DFF_188.Q ;
  assign g6774 = \DFF_161.D ;
  assign g6778 = \DFF_190.D ;
  assign g678 = \DFF_208.Q ;
  assign g6785 = \DFF_161.D ;
  assign g6786 = \DFF_190.D ;
  assign g6787 = \DFF_113.D ;
  assign g6788 = \DFF_173.D ;
  assign g6789 = \DFF_25.D ;
  assign g679 = \DFF_200.Q ;
  assign g6790 = \DFF_20.D ;
  assign g6791 = \DFF_164.D ;
  assign g6792 = \DFF_87.D ;
  assign g6793 = \DFF_50.D ;
  assign g6794 = \DFF_125.D ;
  assign g6796 = \DFF_161.D ;
  assign g6797 = \DFF_190.D ;
  assign g680 = \DFF_129.Q ;
  assign g6800 = \DFF_161.D ;
  assign g6801 = \DFF_190.D ;
  assign g6803 = \DFF_164.D ;
  assign g6806 = \DFF_87.D ;
  assign g6809 = \DFF_50.D ;
  assign g681 = \DFF_207.Q ;
  assign g6812 = \DFF_125.D ;
  assign g6817 = \DFF_113.D ;
  assign g6818 = \DFF_173.D ;
  assign g6819 = \DFF_25.D ;
  assign g682 = \DFF_26.Q ;
  assign g6820 = \DFF_20.D ;
  assign g6824 = \DFF_113.D ;
  assign g6825 = \DFF_173.D ;
  assign g6826 = \DFF_25.D ;
  assign g6827 = \DFF_20.D ;
  assign g683 = \DFF_111.Q ;
  assign g6832 = \DFF_125.D ;
  assign g6833 = \DFF_164.D ;
  assign g6834 = \DFF_161.D ;
  assign g6835 = \DFF_87.D ;
  assign g6836 = \DFF_50.D ;
  assign g6837 = \DFF_190.D ;
  assign g6838 = \DFF_125.D ;
  assign g6839 = \DFF_164.D ;
  assign g684 = \DFF_51.Q ;
  assign g6840 = \DFF_87.D ;
  assign g6841 = \DFF_50.D ;
  assign g6842 = \DFF_125.D ;
  assign g6844 = \DFF_90.D ;
  assign g6845 = \DFF_79.D ;
  assign g6849 = \DFF_90.D ;
  assign g685 = \DFF_47.Q ;
  assign g6850 = \DFF_79.D ;
  assign g6853 = \DFF_90.D ;
  assign g6854 = \DFF_79.D ;
  assign g687 = \DFF_99.Q ;
  assign g688 = \DFF_124.Q ;
  assign g689 = \DFF_9.Q ;
  assign g690 = \DFF_188.Q ;
  assign g691 = \DFF_208.Q ;
  assign g692 = \DFF_200.Q ;
  assign g693 = \DFF_129.Q ;
  assign g694 = \DFF_207.Q ;
  assign g695 = \DFF_26.Q ;
  assign g696 = \DFF_111.Q ;
  assign g697 = \DFF_51.Q ;
  assign g698 = \DFF_92.Q ;
  assign g699 = \DFF_191.Q ;
  assign g7 = \DFF_186.Q ;
  assign g719 = \DFF_178.Q ;
  assign g729 = \DFF_52.Q ;
  assign g736 = \DFF_3.Q ;
  assign g743 = \DFF_37.Q ;
  assign g749 = \DFF_146.Q ;
  assign g754 = \DFF_164.Q ;
  assign g760 = \DFF_87.Q ;
  assign g766 = \DFF_168.Q ;
  assign g774 = \DFF_201.Q ;
  assign g784 = \DFF_17.Q ;
  assign g791 = \DFF_134.Q ;
  assign g798 = \DFF_142.Q ;
  assign g804 = \DFF_61.Q ;
  assign g809 = \DFF_50.Q ;
  assign g815 = \DFF_125.Q ;
  assign g821 = \DFF_43.Q ;
  assign g894 = \DFF_23.Q ;
  assign g898 = \DFF_191.D ;
  assign g899 = \DFF_143.Q ;
  assign g900 = \DFF_143.Q ;
  assign g908 = \DFF_132.Q ;
  assign g909 = \DFF_180.Q ;
  assign g917 = \DFF_148.Q ;
  assign g922 = \DFF_191.Q ;
  assign g927 = g702;
  assign g952 = \DFF_188.Q ;
  assign g965 = \DFF_208.Q ;
  assign g980 = \DFF_200.Q ;
  assign g996 = \DFF_129.Q ;
endmodule
