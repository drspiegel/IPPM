
module s38584(GND, VDD, CK, g100, g10122, g10306, g10500, g10527, g113, g11349, g11388, g114, g11418, g11447, g115, g116, g11678, g11770, g120, g12184, g12238, g12300, g12350, g12368, g124, g12422, g12470, g125, g126, g127, g12832, g12833, g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259, g13272, g134, g135, g13865, g13881, g13895, g13906, g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624, g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744, g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320, g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607, g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711, g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787, g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096, g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612, g23652, g23683, g23759, g24151, g24161, g24162, g24163, g24164, g24165, g24166, g24167, g24168, g24169, g24170, g24171, g24172, g24173, g24174, g24175, g24176, g24177, g24178, g24179, g24180, g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219, g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041, g28042, g28753, g29210, g29211, g29212, g29213, g29214, g29215, g29216, g29217, g29218, g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945, g33946, g33947, g33948, g33949, g33950, g33959, g34201, g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238, g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925, g34927, g34956, g34972, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, g7243, g7245, g7257, g7260, g73, g7540, g7916, g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, g8398, g84, g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, g8920, g90, g9019, g9048, g91, g92, g9251, g9497, g9553, g9555, g9615, g9617, g9680, g9682, g9741, g9743, g9817, g99);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  input CK;
  wire \DFF_0.CK ;
  wire \DFF_0.D ;
  wire \DFF_0.Q ;
  wire \DFF_1.CK ;
  wire \DFF_1.D ;
  wire \DFF_1.Q ;
  wire \DFF_10.CK ;
  wire \DFF_10.D ;
  wire \DFF_10.Q ;
  wire \DFF_100.CK ;
  wire \DFF_100.D ;
  wire \DFF_100.Q ;
  wire \DFF_1000.CK ;
  wire \DFF_1000.D ;
  wire \DFF_1000.Q ;
  wire \DFF_1001.CK ;
  wire \DFF_1001.D ;
  wire \DFF_1001.Q ;
  wire \DFF_1002.CK ;
  wire \DFF_1002.D ;
  wire \DFF_1002.Q ;
  wire \DFF_1003.CK ;
  wire \DFF_1003.D ;
  wire \DFF_1003.Q ;
  wire \DFF_1004.CK ;
  wire \DFF_1004.D ;
  wire \DFF_1004.Q ;
  wire \DFF_1005.CK ;
  wire \DFF_1005.D ;
  wire \DFF_1005.Q ;
  wire \DFF_1006.CK ;
  wire \DFF_1006.D ;
  wire \DFF_1006.Q ;
  wire \DFF_1007.CK ;
  wire \DFF_1007.D ;
  wire \DFF_1007.Q ;
  wire \DFF_1008.CK ;
  wire \DFF_1008.D ;
  wire \DFF_1008.Q ;
  wire \DFF_1009.CK ;
  wire \DFF_1009.D ;
  wire \DFF_1009.Q ;
  wire \DFF_101.CK ;
  wire \DFF_101.D ;
  wire \DFF_101.Q ;
  wire \DFF_1010.CK ;
  wire \DFF_1010.D ;
  wire \DFF_1010.Q ;
  wire \DFF_1011.CK ;
  wire \DFF_1011.D ;
  wire \DFF_1011.Q ;
  wire \DFF_1012.CK ;
  wire \DFF_1012.D ;
  wire \DFF_1012.Q ;
  wire \DFF_1013.CK ;
  wire \DFF_1013.D ;
  wire \DFF_1013.Q ;
  wire \DFF_1014.CK ;
  wire \DFF_1014.D ;
  wire \DFF_1014.Q ;
  wire \DFF_1015.CK ;
  wire \DFF_1015.D ;
  wire \DFF_1015.Q ;
  wire \DFF_1016.CK ;
  wire \DFF_1016.D ;
  wire \DFF_1016.Q ;
  wire \DFF_1017.CK ;
  wire \DFF_1017.D ;
  wire \DFF_1017.Q ;
  wire \DFF_1018.CK ;
  wire \DFF_1018.D ;
  wire \DFF_1018.Q ;
  wire \DFF_1019.CK ;
  wire \DFF_1019.D ;
  wire \DFF_1019.Q ;
  wire \DFF_102.CK ;
  wire \DFF_102.D ;
  wire \DFF_102.Q ;
  wire \DFF_1020.CK ;
  wire \DFF_1020.D ;
  wire \DFF_1020.Q ;
  wire \DFF_1021.CK ;
  wire \DFF_1021.D ;
  wire \DFF_1021.Q ;
  wire \DFF_1022.CK ;
  wire \DFF_1022.D ;
  wire \DFF_1022.Q ;
  wire \DFF_1023.CK ;
  wire \DFF_1023.D ;
  wire \DFF_1023.Q ;
  wire \DFF_1024.CK ;
  wire \DFF_1024.D ;
  wire \DFF_1024.Q ;
  wire \DFF_1025.CK ;
  wire \DFF_1025.D ;
  wire \DFF_1025.Q ;
  wire \DFF_1026.CK ;
  wire \DFF_1026.D ;
  wire \DFF_1026.Q ;
  wire \DFF_1027.CK ;
  wire \DFF_1027.D ;
  wire \DFF_1027.Q ;
  wire \DFF_1028.CK ;
  wire \DFF_1028.D ;
  wire \DFF_1028.Q ;
  wire \DFF_1029.CK ;
  wire \DFF_1029.D ;
  wire \DFF_1029.Q ;
  wire \DFF_103.CK ;
  wire \DFF_103.D ;
  wire \DFF_103.Q ;
  wire \DFF_1030.CK ;
  wire \DFF_1030.D ;
  wire \DFF_1030.Q ;
  wire \DFF_1031.CK ;
  wire \DFF_1031.D ;
  wire \DFF_1031.Q ;
  wire \DFF_1032.CK ;
  wire \DFF_1032.D ;
  wire \DFF_1032.Q ;
  wire \DFF_1033.CK ;
  wire \DFF_1033.D ;
  wire \DFF_1033.Q ;
  wire \DFF_1034.CK ;
  wire \DFF_1034.D ;
  wire \DFF_1034.Q ;
  wire \DFF_1035.CK ;
  wire \DFF_1035.D ;
  wire \DFF_1035.Q ;
  wire \DFF_1036.CK ;
  wire \DFF_1036.D ;
  wire \DFF_1036.Q ;
  wire \DFF_1037.CK ;
  wire \DFF_1037.D ;
  wire \DFF_1037.Q ;
  wire \DFF_1038.CK ;
  wire \DFF_1038.D ;
  wire \DFF_1038.Q ;
  wire \DFF_1039.CK ;
  wire \DFF_1039.D ;
  wire \DFF_1039.Q ;
  wire \DFF_104.CK ;
  wire \DFF_104.D ;
  wire \DFF_104.Q ;
  wire \DFF_1040.CK ;
  wire \DFF_1040.D ;
  wire \DFF_1040.Q ;
  wire \DFF_1041.CK ;
  wire \DFF_1041.D ;
  wire \DFF_1041.Q ;
  wire \DFF_1042.CK ;
  wire \DFF_1042.D ;
  wire \DFF_1042.Q ;
  wire \DFF_1043.CK ;
  wire \DFF_1043.D ;
  wire \DFF_1043.Q ;
  wire \DFF_1044.CK ;
  wire \DFF_1044.D ;
  wire \DFF_1044.Q ;
  wire \DFF_1045.CK ;
  wire \DFF_1045.D ;
  wire \DFF_1045.Q ;
  wire \DFF_1046.CK ;
  wire \DFF_1046.D ;
  wire \DFF_1046.Q ;
  wire \DFF_1047.CK ;
  wire \DFF_1047.D ;
  wire \DFF_1047.Q ;
  wire \DFF_1048.CK ;
  wire \DFF_1048.D ;
  wire \DFF_1048.Q ;
  wire \DFF_1049.CK ;
  wire \DFF_1049.D ;
  wire \DFF_1049.Q ;
  wire \DFF_105.CK ;
  wire \DFF_105.D ;
  wire \DFF_105.Q ;
  wire \DFF_1050.CK ;
  wire \DFF_1050.D ;
  wire \DFF_1050.Q ;
  wire \DFF_1051.CK ;
  wire \DFF_1051.D ;
  wire \DFF_1051.Q ;
  wire \DFF_1052.CK ;
  wire \DFF_1052.D ;
  wire \DFF_1052.Q ;
  wire \DFF_1053.CK ;
  wire \DFF_1053.D ;
  wire \DFF_1053.Q ;
  wire \DFF_1054.CK ;
  wire \DFF_1054.D ;
  wire \DFF_1054.Q ;
  wire \DFF_1055.CK ;
  wire \DFF_1055.D ;
  wire \DFF_1055.Q ;
  wire \DFF_1056.CK ;
  wire \DFF_1056.D ;
  wire \DFF_1056.Q ;
  wire \DFF_1057.CK ;
  wire \DFF_1057.D ;
  wire \DFF_1057.Q ;
  wire \DFF_1058.CK ;
  wire \DFF_1058.D ;
  wire \DFF_1058.Q ;
  wire \DFF_1059.CK ;
  wire \DFF_1059.D ;
  wire \DFF_1059.Q ;
  wire \DFF_106.CK ;
  wire \DFF_106.D ;
  wire \DFF_106.Q ;
  wire \DFF_1060.CK ;
  wire \DFF_1060.D ;
  wire \DFF_1060.Q ;
  wire \DFF_1061.CK ;
  wire \DFF_1061.D ;
  wire \DFF_1061.Q ;
  wire \DFF_1062.CK ;
  wire \DFF_1062.D ;
  wire \DFF_1062.Q ;
  wire \DFF_1063.CK ;
  wire \DFF_1063.D ;
  wire \DFF_1063.Q ;
  wire \DFF_1064.CK ;
  wire \DFF_1064.D ;
  wire \DFF_1064.Q ;
  wire \DFF_1065.CK ;
  wire \DFF_1065.D ;
  wire \DFF_1065.Q ;
  wire \DFF_1066.CK ;
  wire \DFF_1066.D ;
  wire \DFF_1066.Q ;
  wire \DFF_1067.CK ;
  wire \DFF_1067.D ;
  wire \DFF_1067.Q ;
  wire \DFF_1068.CK ;
  wire \DFF_1068.D ;
  wire \DFF_1068.Q ;
  wire \DFF_1069.CK ;
  wire \DFF_1069.D ;
  wire \DFF_1069.Q ;
  wire \DFF_107.CK ;
  wire \DFF_107.D ;
  wire \DFF_107.Q ;
  wire \DFF_1070.CK ;
  wire \DFF_1070.D ;
  wire \DFF_1070.Q ;
  wire \DFF_1071.CK ;
  wire \DFF_1071.D ;
  wire \DFF_1071.Q ;
  wire \DFF_1072.CK ;
  wire \DFF_1072.D ;
  wire \DFF_1072.Q ;
  wire \DFF_1073.CK ;
  wire \DFF_1073.D ;
  wire \DFF_1073.Q ;
  wire \DFF_1074.CK ;
  wire \DFF_1074.D ;
  wire \DFF_1074.Q ;
  wire \DFF_1075.CK ;
  wire \DFF_1075.D ;
  wire \DFF_1075.Q ;
  wire \DFF_1076.CK ;
  wire \DFF_1076.D ;
  wire \DFF_1076.Q ;
  wire \DFF_1077.CK ;
  wire \DFF_1077.D ;
  wire \DFF_1077.Q ;
  wire \DFF_1078.CK ;
  wire \DFF_1078.D ;
  wire \DFF_1078.Q ;
  wire \DFF_1079.CK ;
  wire \DFF_1079.D ;
  wire \DFF_1079.Q ;
  wire \DFF_108.CK ;
  wire \DFF_108.D ;
  wire \DFF_108.Q ;
  wire \DFF_1080.CK ;
  wire \DFF_1080.D ;
  wire \DFF_1080.Q ;
  wire \DFF_1081.CK ;
  wire \DFF_1081.D ;
  wire \DFF_1081.Q ;
  wire \DFF_1082.CK ;
  wire \DFF_1082.D ;
  wire \DFF_1082.Q ;
  wire \DFF_1083.CK ;
  wire \DFF_1083.D ;
  wire \DFF_1083.Q ;
  wire \DFF_1084.CK ;
  wire \DFF_1084.D ;
  wire \DFF_1084.Q ;
  wire \DFF_1085.CK ;
  wire \DFF_1085.D ;
  wire \DFF_1085.Q ;
  wire \DFF_1086.CK ;
  wire \DFF_1086.D ;
  wire \DFF_1086.Q ;
  wire \DFF_1087.CK ;
  wire \DFF_1087.D ;
  wire \DFF_1087.Q ;
  wire \DFF_1088.CK ;
  wire \DFF_1089.CK ;
  wire \DFF_1089.D ;
  wire \DFF_1089.Q ;
  wire \DFF_109.CK ;
  wire \DFF_109.D ;
  wire \DFF_109.Q ;
  wire \DFF_1090.CK ;
  wire \DFF_1090.D ;
  wire \DFF_1090.Q ;
  wire \DFF_1091.CK ;
  wire \DFF_1091.D ;
  wire \DFF_1091.Q ;
  wire \DFF_1092.CK ;
  wire \DFF_1092.D ;
  wire \DFF_1092.Q ;
  wire \DFF_1093.CK ;
  wire \DFF_1093.D ;
  wire \DFF_1093.Q ;
  wire \DFF_1094.CK ;
  wire \DFF_1094.D ;
  wire \DFF_1094.Q ;
  wire \DFF_1095.CK ;
  wire \DFF_1095.D ;
  wire \DFF_1095.Q ;
  wire \DFF_1096.CK ;
  wire \DFF_1096.D ;
  wire \DFF_1096.Q ;
  wire \DFF_1097.CK ;
  wire \DFF_1097.D ;
  wire \DFF_1097.Q ;
  wire \DFF_1098.CK ;
  wire \DFF_1098.D ;
  wire \DFF_1098.Q ;
  wire \DFF_1099.CK ;
  wire \DFF_1099.D ;
  wire \DFF_1099.Q ;
  wire \DFF_11.CK ;
  wire \DFF_11.D ;
  wire \DFF_11.Q ;
  wire \DFF_110.CK ;
  wire \DFF_110.D ;
  wire \DFF_110.Q ;
  wire \DFF_1100.CK ;
  wire \DFF_1100.D ;
  wire \DFF_1100.Q ;
  wire \DFF_1101.CK ;
  wire \DFF_1101.D ;
  wire \DFF_1101.Q ;
  wire \DFF_1102.CK ;
  wire \DFF_1102.D ;
  wire \DFF_1102.Q ;
  wire \DFF_1103.CK ;
  wire \DFF_1103.D ;
  wire \DFF_1103.Q ;
  wire \DFF_1104.CK ;
  wire \DFF_1104.D ;
  wire \DFF_1104.Q ;
  wire \DFF_1105.CK ;
  wire \DFF_1105.D ;
  wire \DFF_1105.Q ;
  wire \DFF_1106.CK ;
  wire \DFF_1106.D ;
  wire \DFF_1106.Q ;
  wire \DFF_1107.CK ;
  wire \DFF_1107.D ;
  wire \DFF_1107.Q ;
  wire \DFF_1108.CK ;
  wire \DFF_1108.D ;
  wire \DFF_1108.Q ;
  wire \DFF_1109.CK ;
  wire \DFF_1109.D ;
  wire \DFF_1109.Q ;
  wire \DFF_111.CK ;
  wire \DFF_111.D ;
  wire \DFF_111.Q ;
  wire \DFF_1110.CK ;
  wire \DFF_1110.D ;
  wire \DFF_1110.Q ;
  wire \DFF_1111.CK ;
  wire \DFF_1111.D ;
  wire \DFF_1111.Q ;
  wire \DFF_1112.CK ;
  wire \DFF_1112.D ;
  wire \DFF_1112.Q ;
  wire \DFF_1113.CK ;
  wire \DFF_1113.D ;
  wire \DFF_1113.Q ;
  wire \DFF_1114.CK ;
  wire \DFF_1114.D ;
  wire \DFF_1114.Q ;
  wire \DFF_1115.CK ;
  wire \DFF_1115.D ;
  wire \DFF_1115.Q ;
  wire \DFF_1116.CK ;
  wire \DFF_1116.D ;
  wire \DFF_1116.Q ;
  wire \DFF_1117.CK ;
  wire \DFF_1117.D ;
  wire \DFF_1117.Q ;
  wire \DFF_1118.CK ;
  wire \DFF_1118.D ;
  wire \DFF_1118.Q ;
  wire \DFF_1119.CK ;
  wire \DFF_1119.D ;
  wire \DFF_1119.Q ;
  wire \DFF_112.CK ;
  wire \DFF_112.D ;
  wire \DFF_112.Q ;
  wire \DFF_1120.CK ;
  wire \DFF_1120.D ;
  wire \DFF_1120.Q ;
  wire \DFF_1121.CK ;
  wire \DFF_1121.D ;
  wire \DFF_1121.Q ;
  wire \DFF_1122.CK ;
  wire \DFF_1122.D ;
  wire \DFF_1122.Q ;
  wire \DFF_1123.CK ;
  wire \DFF_1123.D ;
  wire \DFF_1123.Q ;
  wire \DFF_1124.CK ;
  wire \DFF_1124.D ;
  wire \DFF_1124.Q ;
  wire \DFF_1125.CK ;
  wire \DFF_1125.D ;
  wire \DFF_1125.Q ;
  wire \DFF_1126.CK ;
  wire \DFF_1126.D ;
  wire \DFF_1126.Q ;
  wire \DFF_1127.CK ;
  wire \DFF_1127.D ;
  wire \DFF_1127.Q ;
  wire \DFF_1128.CK ;
  wire \DFF_1128.D ;
  wire \DFF_1128.Q ;
  wire \DFF_1129.CK ;
  wire \DFF_1129.D ;
  wire \DFF_1129.Q ;
  wire \DFF_113.CK ;
  wire \DFF_113.D ;
  wire \DFF_113.Q ;
  wire \DFF_1130.CK ;
  wire \DFF_1130.D ;
  wire \DFF_1130.Q ;
  wire \DFF_1131.CK ;
  wire \DFF_1131.D ;
  wire \DFF_1131.Q ;
  wire \DFF_1132.CK ;
  wire \DFF_1132.D ;
  wire \DFF_1132.Q ;
  wire \DFF_1133.CK ;
  wire \DFF_1133.D ;
  wire \DFF_1133.Q ;
  wire \DFF_1134.CK ;
  wire \DFF_1134.D ;
  wire \DFF_1134.Q ;
  wire \DFF_1135.CK ;
  wire \DFF_1135.D ;
  wire \DFF_1135.Q ;
  wire \DFF_1136.CK ;
  wire \DFF_1136.D ;
  wire \DFF_1136.Q ;
  wire \DFF_1137.CK ;
  wire \DFF_1137.D ;
  wire \DFF_1137.Q ;
  wire \DFF_1138.CK ;
  wire \DFF_1138.D ;
  wire \DFF_1138.Q ;
  wire \DFF_1139.CK ;
  wire \DFF_1139.D ;
  wire \DFF_1139.Q ;
  wire \DFF_114.CK ;
  wire \DFF_114.D ;
  wire \DFF_114.Q ;
  wire \DFF_1140.CK ;
  wire \DFF_1140.D ;
  wire \DFF_1140.Q ;
  wire \DFF_1141.CK ;
  wire \DFF_1141.D ;
  wire \DFF_1141.Q ;
  wire \DFF_1142.CK ;
  wire \DFF_1142.D ;
  wire \DFF_1142.Q ;
  wire \DFF_1143.CK ;
  wire \DFF_1143.D ;
  wire \DFF_1143.Q ;
  wire \DFF_1144.CK ;
  wire \DFF_1144.D ;
  wire \DFF_1144.Q ;
  wire \DFF_1145.CK ;
  wire \DFF_1145.D ;
  wire \DFF_1145.Q ;
  wire \DFF_1146.CK ;
  wire \DFF_1146.D ;
  wire \DFF_1146.Q ;
  wire \DFF_1147.CK ;
  wire \DFF_1147.D ;
  wire \DFF_1147.Q ;
  wire \DFF_1148.CK ;
  wire \DFF_1148.D ;
  wire \DFF_1148.Q ;
  wire \DFF_1149.CK ;
  wire \DFF_1149.D ;
  wire \DFF_1149.Q ;
  wire \DFF_115.CK ;
  wire \DFF_115.D ;
  wire \DFF_115.Q ;
  wire \DFF_1150.CK ;
  wire \DFF_1150.D ;
  wire \DFF_1150.Q ;
  wire \DFF_1151.CK ;
  wire \DFF_1151.D ;
  wire \DFF_1151.Q ;
  wire \DFF_1152.CK ;
  wire \DFF_1152.D ;
  wire \DFF_1152.Q ;
  wire \DFF_1153.CK ;
  wire \DFF_1153.D ;
  wire \DFF_1153.Q ;
  wire \DFF_1154.CK ;
  wire \DFF_1154.D ;
  wire \DFF_1154.Q ;
  wire \DFF_1155.CK ;
  wire \DFF_1155.D ;
  wire \DFF_1155.Q ;
  wire \DFF_1156.CK ;
  wire \DFF_1156.D ;
  wire \DFF_1156.Q ;
  wire \DFF_1157.CK ;
  wire \DFF_1157.D ;
  wire \DFF_1157.Q ;
  wire \DFF_1158.CK ;
  wire \DFF_1158.D ;
  wire \DFF_1158.Q ;
  wire \DFF_1159.CK ;
  wire \DFF_1159.D ;
  wire \DFF_1159.Q ;
  wire \DFF_116.CK ;
  wire \DFF_116.D ;
  wire \DFF_116.Q ;
  wire \DFF_1160.CK ;
  wire \DFF_1160.D ;
  wire \DFF_1160.Q ;
  wire \DFF_1161.CK ;
  wire \DFF_1161.D ;
  wire \DFF_1161.Q ;
  wire \DFF_1162.CK ;
  wire \DFF_1162.D ;
  wire \DFF_1162.Q ;
  wire \DFF_1163.CK ;
  wire \DFF_1163.D ;
  wire \DFF_1163.Q ;
  wire \DFF_1164.CK ;
  wire \DFF_1164.D ;
  wire \DFF_1164.Q ;
  wire \DFF_1165.CK ;
  wire \DFF_1165.D ;
  wire \DFF_1165.Q ;
  wire \DFF_1166.CK ;
  wire \DFF_1166.D ;
  wire \DFF_1166.Q ;
  wire \DFF_1167.CK ;
  wire \DFF_1167.D ;
  wire \DFF_1167.Q ;
  wire \DFF_1168.CK ;
  wire \DFF_1168.D ;
  wire \DFF_1168.Q ;
  wire \DFF_1169.CK ;
  wire \DFF_1169.D ;
  wire \DFF_1169.Q ;
  wire \DFF_117.CK ;
  wire \DFF_117.D ;
  wire \DFF_117.Q ;
  wire \DFF_1170.CK ;
  wire \DFF_1170.D ;
  wire \DFF_1170.Q ;
  wire \DFF_1171.CK ;
  wire \DFF_1171.D ;
  wire \DFF_1171.Q ;
  wire \DFF_1172.CK ;
  wire \DFF_1172.D ;
  wire \DFF_1172.Q ;
  wire \DFF_1173.CK ;
  wire \DFF_1173.D ;
  wire \DFF_1173.Q ;
  wire \DFF_1174.CK ;
  wire \DFF_1174.D ;
  wire \DFF_1174.Q ;
  wire \DFF_1175.CK ;
  wire \DFF_1175.D ;
  wire \DFF_1175.Q ;
  wire \DFF_1176.CK ;
  wire \DFF_1176.D ;
  wire \DFF_1176.Q ;
  wire \DFF_1177.CK ;
  wire \DFF_1177.D ;
  wire \DFF_1177.Q ;
  wire \DFF_1178.CK ;
  wire \DFF_1178.D ;
  wire \DFF_1178.Q ;
  wire \DFF_1179.CK ;
  wire \DFF_1179.D ;
  wire \DFF_1179.Q ;
  wire \DFF_118.CK ;
  wire \DFF_118.D ;
  wire \DFF_118.Q ;
  wire \DFF_1180.CK ;
  wire \DFF_1180.D ;
  wire \DFF_1180.Q ;
  wire \DFF_1181.CK ;
  wire \DFF_1181.D ;
  wire \DFF_1181.Q ;
  wire \DFF_1182.CK ;
  wire \DFF_1182.D ;
  wire \DFF_1182.Q ;
  wire \DFF_1183.CK ;
  wire \DFF_1183.D ;
  wire \DFF_1183.Q ;
  wire \DFF_1184.CK ;
  wire \DFF_1184.D ;
  wire \DFF_1184.Q ;
  wire \DFF_1185.CK ;
  wire \DFF_1185.D ;
  wire \DFF_1185.Q ;
  wire \DFF_1186.CK ;
  wire \DFF_1186.D ;
  wire \DFF_1186.Q ;
  wire \DFF_1187.CK ;
  wire \DFF_1187.D ;
  wire \DFF_1187.Q ;
  wire \DFF_1188.CK ;
  wire \DFF_1188.D ;
  wire \DFF_1188.Q ;
  wire \DFF_1189.CK ;
  wire \DFF_1189.D ;
  wire \DFF_1189.Q ;
  wire \DFF_119.CK ;
  wire \DFF_119.D ;
  wire \DFF_119.Q ;
  wire \DFF_1190.CK ;
  wire \DFF_1190.D ;
  wire \DFF_1190.Q ;
  wire \DFF_1191.CK ;
  wire \DFF_1191.D ;
  wire \DFF_1191.Q ;
  wire \DFF_1192.CK ;
  wire \DFF_1192.D ;
  wire \DFF_1192.Q ;
  wire \DFF_1193.CK ;
  wire \DFF_1193.D ;
  wire \DFF_1193.Q ;
  wire \DFF_1194.CK ;
  wire \DFF_1194.D ;
  wire \DFF_1194.Q ;
  wire \DFF_1195.CK ;
  wire \DFF_1195.D ;
  wire \DFF_1195.Q ;
  wire \DFF_1196.CK ;
  wire \DFF_1196.D ;
  wire \DFF_1196.Q ;
  wire \DFF_1197.CK ;
  wire \DFF_1197.D ;
  wire \DFF_1197.Q ;
  wire \DFF_1198.CK ;
  wire \DFF_1198.D ;
  wire \DFF_1198.Q ;
  wire \DFF_1199.CK ;
  wire \DFF_1199.D ;
  wire \DFF_1199.Q ;
  wire \DFF_12.CK ;
  wire \DFF_12.D ;
  wire \DFF_12.Q ;
  wire \DFF_120.CK ;
  wire \DFF_120.D ;
  wire \DFF_120.Q ;
  wire \DFF_1200.CK ;
  wire \DFF_1200.D ;
  wire \DFF_1200.Q ;
  wire \DFF_1201.CK ;
  wire \DFF_1201.D ;
  wire \DFF_1201.Q ;
  wire \DFF_1202.CK ;
  wire \DFF_1202.D ;
  wire \DFF_1202.Q ;
  wire \DFF_1203.CK ;
  wire \DFF_1203.D ;
  wire \DFF_1203.Q ;
  wire \DFF_1204.CK ;
  wire \DFF_1204.D ;
  wire \DFF_1204.Q ;
  wire \DFF_1205.CK ;
  wire \DFF_1205.D ;
  wire \DFF_1205.Q ;
  wire \DFF_1206.CK ;
  wire \DFF_1206.D ;
  wire \DFF_1206.Q ;
  wire \DFF_1207.CK ;
  wire \DFF_1207.D ;
  wire \DFF_1207.Q ;
  wire \DFF_1208.CK ;
  wire \DFF_1208.D ;
  wire \DFF_1208.Q ;
  wire \DFF_1209.CK ;
  wire \DFF_1209.D ;
  wire \DFF_1209.Q ;
  wire \DFF_121.CK ;
  wire \DFF_121.D ;
  wire \DFF_121.Q ;
  wire \DFF_1210.CK ;
  wire \DFF_1210.D ;
  wire \DFF_1210.Q ;
  wire \DFF_1211.CK ;
  wire \DFF_1211.D ;
  wire \DFF_1211.Q ;
  wire \DFF_1212.CK ;
  wire \DFF_1212.D ;
  wire \DFF_1212.Q ;
  wire \DFF_1213.CK ;
  wire \DFF_1213.D ;
  wire \DFF_1213.Q ;
  wire \DFF_1214.CK ;
  wire \DFF_1214.D ;
  wire \DFF_1214.Q ;
  wire \DFF_1215.CK ;
  wire \DFF_1215.D ;
  wire \DFF_1215.Q ;
  wire \DFF_1216.CK ;
  wire \DFF_1216.D ;
  wire \DFF_1216.Q ;
  wire \DFF_1217.CK ;
  wire \DFF_1217.D ;
  wire \DFF_1217.Q ;
  wire \DFF_1218.CK ;
  wire \DFF_1218.D ;
  wire \DFF_1218.Q ;
  wire \DFF_1219.CK ;
  wire \DFF_1219.D ;
  wire \DFF_1219.Q ;
  wire \DFF_122.CK ;
  wire \DFF_122.D ;
  wire \DFF_122.Q ;
  wire \DFF_1220.CK ;
  wire \DFF_1220.D ;
  wire \DFF_1220.Q ;
  wire \DFF_1221.CK ;
  wire \DFF_1221.D ;
  wire \DFF_1221.Q ;
  wire \DFF_1222.CK ;
  wire \DFF_1222.D ;
  wire \DFF_1222.Q ;
  wire \DFF_1223.CK ;
  wire \DFF_1223.D ;
  wire \DFF_1223.Q ;
  wire \DFF_1224.CK ;
  wire \DFF_1224.D ;
  wire \DFF_1224.Q ;
  wire \DFF_1225.CK ;
  wire \DFF_1225.D ;
  wire \DFF_1225.Q ;
  wire \DFF_1226.CK ;
  wire \DFF_1226.D ;
  wire \DFF_1226.Q ;
  wire \DFF_1227.CK ;
  wire \DFF_1227.D ;
  wire \DFF_1227.Q ;
  wire \DFF_1228.CK ;
  wire \DFF_1228.D ;
  wire \DFF_1228.Q ;
  wire \DFF_1229.CK ;
  wire \DFF_1229.D ;
  wire \DFF_1229.Q ;
  wire \DFF_123.CK ;
  wire \DFF_123.D ;
  wire \DFF_123.Q ;
  wire \DFF_1230.CK ;
  wire \DFF_1230.D ;
  wire \DFF_1230.Q ;
  wire \DFF_1231.CK ;
  wire \DFF_1231.D ;
  wire \DFF_1231.Q ;
  wire \DFF_1232.CK ;
  wire \DFF_1232.D ;
  wire \DFF_1232.Q ;
  wire \DFF_1233.CK ;
  wire \DFF_1233.D ;
  wire \DFF_1233.Q ;
  wire \DFF_1234.CK ;
  wire \DFF_1234.D ;
  wire \DFF_1234.Q ;
  wire \DFF_1235.CK ;
  wire \DFF_1235.D ;
  wire \DFF_1235.Q ;
  wire \DFF_1236.CK ;
  wire \DFF_1236.D ;
  wire \DFF_1236.Q ;
  wire \DFF_1237.CK ;
  wire \DFF_1237.D ;
  wire \DFF_1237.Q ;
  wire \DFF_1238.CK ;
  wire \DFF_1238.D ;
  wire \DFF_1238.Q ;
  wire \DFF_1239.CK ;
  wire \DFF_1239.D ;
  wire \DFF_1239.Q ;
  wire \DFF_124.CK ;
  wire \DFF_124.D ;
  wire \DFF_124.Q ;
  wire \DFF_1240.CK ;
  wire \DFF_1240.D ;
  wire \DFF_1240.Q ;
  wire \DFF_1241.CK ;
  wire \DFF_1241.D ;
  wire \DFF_1241.Q ;
  wire \DFF_1242.CK ;
  wire \DFF_1242.D ;
  wire \DFF_1242.Q ;
  wire \DFF_1243.CK ;
  wire \DFF_1243.D ;
  wire \DFF_1243.Q ;
  wire \DFF_1244.CK ;
  wire \DFF_1244.D ;
  wire \DFF_1244.Q ;
  wire \DFF_1245.CK ;
  wire \DFF_1245.D ;
  wire \DFF_1245.Q ;
  wire \DFF_1246.CK ;
  wire \DFF_1246.D ;
  wire \DFF_1246.Q ;
  wire \DFF_1247.CK ;
  wire \DFF_1247.D ;
  wire \DFF_1247.Q ;
  wire \DFF_1248.CK ;
  wire \DFF_1248.D ;
  wire \DFF_1248.Q ;
  wire \DFF_1249.CK ;
  wire \DFF_1249.D ;
  wire \DFF_1249.Q ;
  wire \DFF_125.CK ;
  wire \DFF_125.D ;
  wire \DFF_125.Q ;
  wire \DFF_1250.CK ;
  wire \DFF_1250.D ;
  wire \DFF_1250.Q ;
  wire \DFF_1251.CK ;
  wire \DFF_1251.D ;
  wire \DFF_1251.Q ;
  wire \DFF_1252.CK ;
  wire \DFF_1252.D ;
  wire \DFF_1252.Q ;
  wire \DFF_1253.CK ;
  wire \DFF_1253.D ;
  wire \DFF_1253.Q ;
  wire \DFF_1254.CK ;
  wire \DFF_1254.D ;
  wire \DFF_1254.Q ;
  wire \DFF_1255.CK ;
  wire \DFF_1255.D ;
  wire \DFF_1255.Q ;
  wire \DFF_1256.CK ;
  wire \DFF_1256.D ;
  wire \DFF_1256.Q ;
  wire \DFF_1257.CK ;
  wire \DFF_1257.D ;
  wire \DFF_1257.Q ;
  wire \DFF_1258.CK ;
  wire \DFF_1258.D ;
  wire \DFF_1258.Q ;
  wire \DFF_1259.CK ;
  wire \DFF_1259.D ;
  wire \DFF_1259.Q ;
  wire \DFF_126.CK ;
  wire \DFF_126.D ;
  wire \DFF_126.Q ;
  wire \DFF_1260.CK ;
  wire \DFF_1260.D ;
  wire \DFF_1260.Q ;
  wire \DFF_1261.CK ;
  wire \DFF_1261.D ;
  wire \DFF_1261.Q ;
  wire \DFF_1262.CK ;
  wire \DFF_1262.D ;
  wire \DFF_1262.Q ;
  wire \DFF_1263.CK ;
  wire \DFF_1263.D ;
  wire \DFF_1263.Q ;
  wire \DFF_1264.CK ;
  wire \DFF_1264.D ;
  wire \DFF_1264.Q ;
  wire \DFF_1265.CK ;
  wire \DFF_1265.D ;
  wire \DFF_1265.Q ;
  wire \DFF_1266.CK ;
  wire \DFF_1266.D ;
  wire \DFF_1266.Q ;
  wire \DFF_1267.CK ;
  wire \DFF_1267.D ;
  wire \DFF_1267.Q ;
  wire \DFF_1268.CK ;
  wire \DFF_1268.D ;
  wire \DFF_1268.Q ;
  wire \DFF_1269.CK ;
  wire \DFF_1269.D ;
  wire \DFF_1269.Q ;
  wire \DFF_127.CK ;
  wire \DFF_127.D ;
  wire \DFF_127.Q ;
  wire \DFF_1270.CK ;
  wire \DFF_1270.D ;
  wire \DFF_1270.Q ;
  wire \DFF_1271.CK ;
  wire \DFF_1271.D ;
  wire \DFF_1271.Q ;
  wire \DFF_1272.CK ;
  wire \DFF_1272.D ;
  wire \DFF_1272.Q ;
  wire \DFF_1273.CK ;
  wire \DFF_1273.D ;
  wire \DFF_1273.Q ;
  wire \DFF_1274.CK ;
  wire \DFF_1274.D ;
  wire \DFF_1274.Q ;
  wire \DFF_1275.CK ;
  wire \DFF_1275.D ;
  wire \DFF_1275.Q ;
  wire \DFF_1276.CK ;
  wire \DFF_1276.D ;
  wire \DFF_1276.Q ;
  wire \DFF_1277.CK ;
  wire \DFF_1277.D ;
  wire \DFF_1277.Q ;
  wire \DFF_1278.CK ;
  wire \DFF_1278.D ;
  wire \DFF_1278.Q ;
  wire \DFF_1279.CK ;
  wire \DFF_1279.D ;
  wire \DFF_1279.Q ;
  wire \DFF_128.CK ;
  wire \DFF_128.D ;
  wire \DFF_128.Q ;
  wire \DFF_1280.CK ;
  wire \DFF_1280.D ;
  wire \DFF_1280.Q ;
  wire \DFF_1281.CK ;
  wire \DFF_1281.D ;
  wire \DFF_1281.Q ;
  wire \DFF_1282.CK ;
  wire \DFF_1282.D ;
  wire \DFF_1282.Q ;
  wire \DFF_1283.CK ;
  wire \DFF_1283.D ;
  wire \DFF_1283.Q ;
  wire \DFF_1284.CK ;
  wire \DFF_1284.D ;
  wire \DFF_1284.Q ;
  wire \DFF_1285.CK ;
  wire \DFF_1285.D ;
  wire \DFF_1285.Q ;
  wire \DFF_1286.CK ;
  wire \DFF_1286.D ;
  wire \DFF_1286.Q ;
  wire \DFF_1287.CK ;
  wire \DFF_1287.D ;
  wire \DFF_1287.Q ;
  wire \DFF_1288.CK ;
  wire \DFF_1288.D ;
  wire \DFF_1288.Q ;
  wire \DFF_1289.CK ;
  wire \DFF_1289.D ;
  wire \DFF_1289.Q ;
  wire \DFF_129.CK ;
  wire \DFF_129.D ;
  wire \DFF_129.Q ;
  wire \DFF_1290.CK ;
  wire \DFF_1290.D ;
  wire \DFF_1290.Q ;
  wire \DFF_1291.CK ;
  wire \DFF_1291.D ;
  wire \DFF_1291.Q ;
  wire \DFF_1292.CK ;
  wire \DFF_1292.D ;
  wire \DFF_1292.Q ;
  wire \DFF_1293.CK ;
  wire \DFF_1293.D ;
  wire \DFF_1293.Q ;
  wire \DFF_1294.CK ;
  wire \DFF_1294.D ;
  wire \DFF_1294.Q ;
  wire \DFF_1295.CK ;
  wire \DFF_1295.D ;
  wire \DFF_1295.Q ;
  wire \DFF_1296.CK ;
  wire \DFF_1296.D ;
  wire \DFF_1296.Q ;
  wire \DFF_1297.CK ;
  wire \DFF_1297.D ;
  wire \DFF_1297.Q ;
  wire \DFF_1298.CK ;
  wire \DFF_1298.D ;
  wire \DFF_1298.Q ;
  wire \DFF_1299.CK ;
  wire \DFF_1299.D ;
  wire \DFF_1299.Q ;
  wire \DFF_13.CK ;
  wire \DFF_13.D ;
  wire \DFF_13.Q ;
  wire \DFF_130.CK ;
  wire \DFF_130.D ;
  wire \DFF_130.Q ;
  wire \DFF_1300.CK ;
  wire \DFF_1300.D ;
  wire \DFF_1300.Q ;
  wire \DFF_1301.CK ;
  wire \DFF_1301.D ;
  wire \DFF_1301.Q ;
  wire \DFF_1302.CK ;
  wire \DFF_1302.D ;
  wire \DFF_1302.Q ;
  wire \DFF_1303.CK ;
  wire \DFF_1303.D ;
  wire \DFF_1303.Q ;
  wire \DFF_1304.CK ;
  wire \DFF_1304.D ;
  wire \DFF_1304.Q ;
  wire \DFF_1305.CK ;
  wire \DFF_1305.D ;
  wire \DFF_1305.Q ;
  wire \DFF_1306.CK ;
  wire \DFF_1306.D ;
  wire \DFF_1306.Q ;
  wire \DFF_1307.CK ;
  wire \DFF_1307.D ;
  wire \DFF_1307.Q ;
  wire \DFF_1308.CK ;
  wire \DFF_1308.D ;
  wire \DFF_1308.Q ;
  wire \DFF_1309.CK ;
  wire \DFF_1309.D ;
  wire \DFF_1309.Q ;
  wire \DFF_131.CK ;
  wire \DFF_131.D ;
  wire \DFF_131.Q ;
  wire \DFF_1310.CK ;
  wire \DFF_1310.D ;
  wire \DFF_1310.Q ;
  wire \DFF_1311.CK ;
  wire \DFF_1311.D ;
  wire \DFF_1311.Q ;
  wire \DFF_1312.CK ;
  wire \DFF_1312.D ;
  wire \DFF_1312.Q ;
  wire \DFF_1313.CK ;
  wire \DFF_1313.D ;
  wire \DFF_1313.Q ;
  wire \DFF_1314.CK ;
  wire \DFF_1314.D ;
  wire \DFF_1314.Q ;
  wire \DFF_1315.CK ;
  wire \DFF_1315.D ;
  wire \DFF_1315.Q ;
  wire \DFF_1316.CK ;
  wire \DFF_1316.D ;
  wire \DFF_1316.Q ;
  wire \DFF_1317.CK ;
  wire \DFF_1317.D ;
  wire \DFF_1317.Q ;
  wire \DFF_1318.CK ;
  wire \DFF_1318.D ;
  wire \DFF_1318.Q ;
  wire \DFF_1319.CK ;
  wire \DFF_1319.D ;
  wire \DFF_1319.Q ;
  wire \DFF_132.CK ;
  wire \DFF_132.D ;
  wire \DFF_132.Q ;
  wire \DFF_1320.CK ;
  wire \DFF_1320.D ;
  wire \DFF_1320.Q ;
  wire \DFF_1321.CK ;
  wire \DFF_1321.D ;
  wire \DFF_1321.Q ;
  wire \DFF_1322.CK ;
  wire \DFF_1322.D ;
  wire \DFF_1322.Q ;
  wire \DFF_1323.CK ;
  wire \DFF_1323.D ;
  wire \DFF_1323.Q ;
  wire \DFF_1324.CK ;
  wire \DFF_1324.D ;
  wire \DFF_1324.Q ;
  wire \DFF_1325.CK ;
  wire \DFF_1325.D ;
  wire \DFF_1325.Q ;
  wire \DFF_1326.CK ;
  wire \DFF_1326.D ;
  wire \DFF_1326.Q ;
  wire \DFF_1327.CK ;
  wire \DFF_1327.D ;
  wire \DFF_1327.Q ;
  wire \DFF_1328.CK ;
  wire \DFF_1328.D ;
  wire \DFF_1328.Q ;
  wire \DFF_1329.CK ;
  wire \DFF_1329.D ;
  wire \DFF_1329.Q ;
  wire \DFF_133.CK ;
  wire \DFF_133.D ;
  wire \DFF_133.Q ;
  wire \DFF_1330.CK ;
  wire \DFF_1330.D ;
  wire \DFF_1330.Q ;
  wire \DFF_1331.CK ;
  wire \DFF_1331.D ;
  wire \DFF_1331.Q ;
  wire \DFF_1332.CK ;
  wire \DFF_1332.D ;
  wire \DFF_1332.Q ;
  wire \DFF_1333.CK ;
  wire \DFF_1333.D ;
  wire \DFF_1333.Q ;
  wire \DFF_1334.CK ;
  wire \DFF_1334.D ;
  wire \DFF_1334.Q ;
  wire \DFF_1335.CK ;
  wire \DFF_1335.D ;
  wire \DFF_1335.Q ;
  wire \DFF_1336.CK ;
  wire \DFF_1336.D ;
  wire \DFF_1336.Q ;
  wire \DFF_1337.CK ;
  wire \DFF_1337.D ;
  wire \DFF_1337.Q ;
  wire \DFF_1338.CK ;
  wire \DFF_1338.D ;
  wire \DFF_1338.Q ;
  wire \DFF_1339.CK ;
  wire \DFF_1339.D ;
  wire \DFF_1339.Q ;
  wire \DFF_134.CK ;
  wire \DFF_134.D ;
  wire \DFF_134.Q ;
  wire \DFF_1340.CK ;
  wire \DFF_1340.D ;
  wire \DFF_1340.Q ;
  wire \DFF_1341.CK ;
  wire \DFF_1341.D ;
  wire \DFF_1341.Q ;
  wire \DFF_1342.CK ;
  wire \DFF_1342.D ;
  wire \DFF_1342.Q ;
  wire \DFF_1343.CK ;
  wire \DFF_1343.D ;
  wire \DFF_1343.Q ;
  wire \DFF_1344.CK ;
  wire \DFF_1344.D ;
  wire \DFF_1344.Q ;
  wire \DFF_1345.CK ;
  wire \DFF_1345.D ;
  wire \DFF_1345.Q ;
  wire \DFF_1346.CK ;
  wire \DFF_1346.D ;
  wire \DFF_1346.Q ;
  wire \DFF_1347.CK ;
  wire \DFF_1347.D ;
  wire \DFF_1347.Q ;
  wire \DFF_1348.CK ;
  wire \DFF_1348.D ;
  wire \DFF_1348.Q ;
  wire \DFF_1349.CK ;
  wire \DFF_1349.D ;
  wire \DFF_1349.Q ;
  wire \DFF_135.CK ;
  wire \DFF_135.D ;
  wire \DFF_135.Q ;
  wire \DFF_1350.CK ;
  wire \DFF_1350.D ;
  wire \DFF_1350.Q ;
  wire \DFF_1351.CK ;
  wire \DFF_1351.D ;
  wire \DFF_1351.Q ;
  wire \DFF_1352.CK ;
  wire \DFF_1352.D ;
  wire \DFF_1352.Q ;
  wire \DFF_1353.CK ;
  wire \DFF_1353.D ;
  wire \DFF_1353.Q ;
  wire \DFF_1354.CK ;
  wire \DFF_1354.D ;
  wire \DFF_1354.Q ;
  wire \DFF_1355.CK ;
  wire \DFF_1355.D ;
  wire \DFF_1355.Q ;
  wire \DFF_1356.CK ;
  wire \DFF_1356.D ;
  wire \DFF_1356.Q ;
  wire \DFF_1357.CK ;
  wire \DFF_1357.D ;
  wire \DFF_1357.Q ;
  wire \DFF_1358.CK ;
  wire \DFF_1358.D ;
  wire \DFF_1358.Q ;
  wire \DFF_1359.CK ;
  wire \DFF_1359.D ;
  wire \DFF_1359.Q ;
  wire \DFF_136.CK ;
  wire \DFF_136.D ;
  wire \DFF_136.Q ;
  wire \DFF_1360.CK ;
  wire \DFF_1360.D ;
  wire \DFF_1360.Q ;
  wire \DFF_1361.CK ;
  wire \DFF_1361.D ;
  wire \DFF_1361.Q ;
  wire \DFF_1362.CK ;
  wire \DFF_1362.D ;
  wire \DFF_1362.Q ;
  wire \DFF_1363.CK ;
  wire \DFF_1363.D ;
  wire \DFF_1363.Q ;
  wire \DFF_1364.CK ;
  wire \DFF_1364.D ;
  wire \DFF_1364.Q ;
  wire \DFF_1365.CK ;
  wire \DFF_1365.D ;
  wire \DFF_1365.Q ;
  wire \DFF_1366.CK ;
  wire \DFF_1366.D ;
  wire \DFF_1366.Q ;
  wire \DFF_1367.CK ;
  wire \DFF_1367.D ;
  wire \DFF_1367.Q ;
  wire \DFF_1368.CK ;
  wire \DFF_1368.D ;
  wire \DFF_1368.Q ;
  wire \DFF_1369.CK ;
  wire \DFF_1369.D ;
  wire \DFF_1369.Q ;
  wire \DFF_137.CK ;
  wire \DFF_137.D ;
  wire \DFF_137.Q ;
  wire \DFF_1370.CK ;
  wire \DFF_1370.D ;
  wire \DFF_1370.Q ;
  wire \DFF_1371.CK ;
  wire \DFF_1371.D ;
  wire \DFF_1371.Q ;
  wire \DFF_1372.CK ;
  wire \DFF_1372.D ;
  wire \DFF_1372.Q ;
  wire \DFF_1373.CK ;
  wire \DFF_1373.D ;
  wire \DFF_1373.Q ;
  wire \DFF_1374.CK ;
  wire \DFF_1374.D ;
  wire \DFF_1374.Q ;
  wire \DFF_1375.CK ;
  wire \DFF_1375.D ;
  wire \DFF_1375.Q ;
  wire \DFF_1376.CK ;
  wire \DFF_1376.D ;
  wire \DFF_1376.Q ;
  wire \DFF_1377.CK ;
  wire \DFF_1377.D ;
  wire \DFF_1377.Q ;
  wire \DFF_1378.CK ;
  wire \DFF_1378.D ;
  wire \DFF_1378.Q ;
  wire \DFF_1379.CK ;
  wire \DFF_1379.D ;
  wire \DFF_1379.Q ;
  wire \DFF_138.CK ;
  wire \DFF_138.D ;
  wire \DFF_138.Q ;
  wire \DFF_1380.CK ;
  wire \DFF_1380.D ;
  wire \DFF_1380.Q ;
  wire \DFF_1381.CK ;
  wire \DFF_1381.D ;
  wire \DFF_1381.Q ;
  wire \DFF_1382.CK ;
  wire \DFF_1382.D ;
  wire \DFF_1382.Q ;
  wire \DFF_1383.CK ;
  wire \DFF_1383.D ;
  wire \DFF_1383.Q ;
  wire \DFF_1384.CK ;
  wire \DFF_1384.D ;
  wire \DFF_1384.Q ;
  wire \DFF_1385.CK ;
  wire \DFF_1385.D ;
  wire \DFF_1385.Q ;
  wire \DFF_1386.CK ;
  wire \DFF_1386.D ;
  wire \DFF_1386.Q ;
  wire \DFF_1387.CK ;
  wire \DFF_1387.D ;
  wire \DFF_1387.Q ;
  wire \DFF_1388.CK ;
  wire \DFF_1388.D ;
  wire \DFF_1388.Q ;
  wire \DFF_1389.CK ;
  wire \DFF_1389.D ;
  wire \DFF_1389.Q ;
  wire \DFF_139.CK ;
  wire \DFF_139.D ;
  wire \DFF_139.Q ;
  wire \DFF_1390.CK ;
  wire \DFF_1390.D ;
  wire \DFF_1390.Q ;
  wire \DFF_1391.CK ;
  wire \DFF_1391.D ;
  wire \DFF_1391.Q ;
  wire \DFF_1392.CK ;
  wire \DFF_1392.D ;
  wire \DFF_1392.Q ;
  wire \DFF_1393.CK ;
  wire \DFF_1393.D ;
  wire \DFF_1393.Q ;
  wire \DFF_1394.CK ;
  wire \DFF_1394.D ;
  wire \DFF_1394.Q ;
  wire \DFF_1395.CK ;
  wire \DFF_1395.D ;
  wire \DFF_1395.Q ;
  wire \DFF_1396.CK ;
  wire \DFF_1396.D ;
  wire \DFF_1396.Q ;
  wire \DFF_1397.CK ;
  wire \DFF_1397.D ;
  wire \DFF_1397.Q ;
  wire \DFF_1398.CK ;
  wire \DFF_1398.D ;
  wire \DFF_1398.Q ;
  wire \DFF_1399.CK ;
  wire \DFF_1399.D ;
  wire \DFF_1399.Q ;
  wire \DFF_14.CK ;
  wire \DFF_14.D ;
  wire \DFF_14.Q ;
  wire \DFF_140.CK ;
  wire \DFF_140.D ;
  wire \DFF_140.Q ;
  wire \DFF_1400.CK ;
  wire \DFF_1400.D ;
  wire \DFF_1400.Q ;
  wire \DFF_1401.CK ;
  wire \DFF_1401.D ;
  wire \DFF_1401.Q ;
  wire \DFF_1402.CK ;
  wire \DFF_1402.D ;
  wire \DFF_1402.Q ;
  wire \DFF_1403.CK ;
  wire \DFF_1403.D ;
  wire \DFF_1403.Q ;
  wire \DFF_1404.CK ;
  wire \DFF_1404.D ;
  wire \DFF_1404.Q ;
  wire \DFF_1405.CK ;
  wire \DFF_1405.D ;
  wire \DFF_1405.Q ;
  wire \DFF_1406.CK ;
  wire \DFF_1406.D ;
  wire \DFF_1406.Q ;
  wire \DFF_1407.CK ;
  wire \DFF_1407.D ;
  wire \DFF_1407.Q ;
  wire \DFF_1408.CK ;
  wire \DFF_1408.D ;
  wire \DFF_1408.Q ;
  wire \DFF_1409.CK ;
  wire \DFF_1409.D ;
  wire \DFF_1409.Q ;
  wire \DFF_141.CK ;
  wire \DFF_141.D ;
  wire \DFF_141.Q ;
  wire \DFF_1410.CK ;
  wire \DFF_1410.D ;
  wire \DFF_1410.Q ;
  wire \DFF_1411.CK ;
  wire \DFF_1411.D ;
  wire \DFF_1411.Q ;
  wire \DFF_1412.CK ;
  wire \DFF_1412.D ;
  wire \DFF_1412.Q ;
  wire \DFF_1413.CK ;
  wire \DFF_1413.D ;
  wire \DFF_1413.Q ;
  wire \DFF_1414.CK ;
  wire \DFF_1414.D ;
  wire \DFF_1414.Q ;
  wire \DFF_1415.CK ;
  wire \DFF_1415.D ;
  wire \DFF_1415.Q ;
  wire \DFF_1416.CK ;
  wire \DFF_1416.D ;
  wire \DFF_1416.Q ;
  wire \DFF_1417.CK ;
  wire \DFF_1417.D ;
  wire \DFF_1417.Q ;
  wire \DFF_1418.CK ;
  wire \DFF_1418.D ;
  wire \DFF_1418.Q ;
  wire \DFF_1419.CK ;
  wire \DFF_1419.D ;
  wire \DFF_1419.Q ;
  wire \DFF_142.CK ;
  wire \DFF_142.D ;
  wire \DFF_142.Q ;
  wire \DFF_1420.CK ;
  wire \DFF_1420.D ;
  wire \DFF_1420.Q ;
  wire \DFF_1421.CK ;
  wire \DFF_1422.CK ;
  wire \DFF_1422.D ;
  wire \DFF_1422.Q ;
  wire \DFF_1423.CK ;
  wire \DFF_1423.D ;
  wire \DFF_1423.Q ;
  wire \DFF_1424.CK ;
  wire \DFF_1424.D ;
  wire \DFF_1424.Q ;
  wire \DFF_1425.CK ;
  wire \DFF_1425.D ;
  wire \DFF_1425.Q ;
  wire \DFF_143.CK ;
  wire \DFF_143.D ;
  wire \DFF_143.Q ;
  wire \DFF_144.CK ;
  wire \DFF_144.D ;
  wire \DFF_144.Q ;
  wire \DFF_145.CK ;
  wire \DFF_145.D ;
  wire \DFF_145.Q ;
  wire \DFF_146.CK ;
  wire \DFF_146.D ;
  wire \DFF_146.Q ;
  wire \DFF_147.CK ;
  wire \DFF_147.D ;
  wire \DFF_147.Q ;
  wire \DFF_148.CK ;
  wire \DFF_148.D ;
  wire \DFF_148.Q ;
  wire \DFF_149.CK ;
  wire \DFF_149.D ;
  wire \DFF_149.Q ;
  wire \DFF_15.CK ;
  wire \DFF_15.D ;
  wire \DFF_15.Q ;
  wire \DFF_150.CK ;
  wire \DFF_150.D ;
  wire \DFF_150.Q ;
  wire \DFF_151.CK ;
  wire \DFF_151.D ;
  wire \DFF_151.Q ;
  wire \DFF_152.CK ;
  wire \DFF_152.D ;
  wire \DFF_152.Q ;
  wire \DFF_153.CK ;
  wire \DFF_153.D ;
  wire \DFF_153.Q ;
  wire \DFF_154.CK ;
  wire \DFF_154.D ;
  wire \DFF_154.Q ;
  wire \DFF_155.CK ;
  wire \DFF_155.D ;
  wire \DFF_155.Q ;
  wire \DFF_156.CK ;
  wire \DFF_156.D ;
  wire \DFF_156.Q ;
  wire \DFF_157.CK ;
  wire \DFF_157.D ;
  wire \DFF_157.Q ;
  wire \DFF_158.CK ;
  wire \DFF_158.D ;
  wire \DFF_158.Q ;
  wire \DFF_159.CK ;
  wire \DFF_159.D ;
  wire \DFF_159.Q ;
  wire \DFF_16.CK ;
  wire \DFF_16.D ;
  wire \DFF_16.Q ;
  wire \DFF_160.CK ;
  wire \DFF_160.D ;
  wire \DFF_160.Q ;
  wire \DFF_161.CK ;
  wire \DFF_161.D ;
  wire \DFF_161.Q ;
  wire \DFF_162.CK ;
  wire \DFF_162.D ;
  wire \DFF_162.Q ;
  wire \DFF_163.CK ;
  wire \DFF_163.D ;
  wire \DFF_163.Q ;
  wire \DFF_164.CK ;
  wire \DFF_164.D ;
  wire \DFF_164.Q ;
  wire \DFF_165.CK ;
  wire \DFF_165.D ;
  wire \DFF_165.Q ;
  wire \DFF_166.CK ;
  wire \DFF_166.D ;
  wire \DFF_166.Q ;
  wire \DFF_167.CK ;
  wire \DFF_167.D ;
  wire \DFF_167.Q ;
  wire \DFF_168.CK ;
  wire \DFF_168.D ;
  wire \DFF_168.Q ;
  wire \DFF_169.CK ;
  wire \DFF_169.D ;
  wire \DFF_169.Q ;
  wire \DFF_17.CK ;
  wire \DFF_17.D ;
  wire \DFF_17.Q ;
  wire \DFF_170.CK ;
  wire \DFF_170.D ;
  wire \DFF_170.Q ;
  wire \DFF_171.CK ;
  wire \DFF_171.D ;
  wire \DFF_171.Q ;
  wire \DFF_172.CK ;
  wire \DFF_172.D ;
  wire \DFF_172.Q ;
  wire \DFF_173.CK ;
  wire \DFF_173.D ;
  wire \DFF_173.Q ;
  wire \DFF_174.CK ;
  wire \DFF_174.D ;
  wire \DFF_174.Q ;
  wire \DFF_175.CK ;
  wire \DFF_175.D ;
  wire \DFF_175.Q ;
  wire \DFF_176.CK ;
  wire \DFF_176.D ;
  wire \DFF_176.Q ;
  wire \DFF_177.CK ;
  wire \DFF_177.D ;
  wire \DFF_177.Q ;
  wire \DFF_178.CK ;
  wire \DFF_178.D ;
  wire \DFF_178.Q ;
  wire \DFF_179.CK ;
  wire \DFF_179.D ;
  wire \DFF_179.Q ;
  wire \DFF_18.CK ;
  wire \DFF_18.D ;
  wire \DFF_18.Q ;
  wire \DFF_180.CK ;
  wire \DFF_180.D ;
  wire \DFF_180.Q ;
  wire \DFF_181.CK ;
  wire \DFF_181.D ;
  wire \DFF_181.Q ;
  wire \DFF_182.CK ;
  wire \DFF_182.D ;
  wire \DFF_182.Q ;
  wire \DFF_183.CK ;
  wire \DFF_183.D ;
  wire \DFF_183.Q ;
  wire \DFF_184.CK ;
  wire \DFF_184.D ;
  wire \DFF_184.Q ;
  wire \DFF_185.CK ;
  wire \DFF_185.D ;
  wire \DFF_185.Q ;
  wire \DFF_186.CK ;
  wire \DFF_186.D ;
  wire \DFF_186.Q ;
  wire \DFF_187.CK ;
  wire \DFF_187.D ;
  wire \DFF_187.Q ;
  wire \DFF_188.CK ;
  wire \DFF_188.D ;
  wire \DFF_188.Q ;
  wire \DFF_189.CK ;
  wire \DFF_189.D ;
  wire \DFF_189.Q ;
  wire \DFF_19.CK ;
  wire \DFF_19.D ;
  wire \DFF_19.Q ;
  wire \DFF_190.CK ;
  wire \DFF_190.D ;
  wire \DFF_190.Q ;
  wire \DFF_191.CK ;
  wire \DFF_191.D ;
  wire \DFF_191.Q ;
  wire \DFF_192.CK ;
  wire \DFF_192.D ;
  wire \DFF_192.Q ;
  wire \DFF_193.CK ;
  wire \DFF_193.D ;
  wire \DFF_193.Q ;
  wire \DFF_194.CK ;
  wire \DFF_194.D ;
  wire \DFF_194.Q ;
  wire \DFF_195.CK ;
  wire \DFF_195.D ;
  wire \DFF_195.Q ;
  wire \DFF_196.CK ;
  wire \DFF_196.D ;
  wire \DFF_196.Q ;
  wire \DFF_197.CK ;
  wire \DFF_197.D ;
  wire \DFF_197.Q ;
  wire \DFF_198.CK ;
  wire \DFF_198.D ;
  wire \DFF_198.Q ;
  wire \DFF_199.CK ;
  wire \DFF_199.D ;
  wire \DFF_199.Q ;
  wire \DFF_2.CK ;
  wire \DFF_2.D ;
  wire \DFF_2.Q ;
  wire \DFF_20.CK ;
  wire \DFF_20.D ;
  wire \DFF_20.Q ;
  wire \DFF_200.CK ;
  wire \DFF_200.D ;
  wire \DFF_200.Q ;
  wire \DFF_201.CK ;
  wire \DFF_201.D ;
  wire \DFF_201.Q ;
  wire \DFF_202.CK ;
  wire \DFF_202.D ;
  wire \DFF_202.Q ;
  wire \DFF_203.CK ;
  wire \DFF_203.D ;
  wire \DFF_203.Q ;
  wire \DFF_204.CK ;
  wire \DFF_204.D ;
  wire \DFF_204.Q ;
  wire \DFF_205.CK ;
  wire \DFF_205.D ;
  wire \DFF_205.Q ;
  wire \DFF_206.CK ;
  wire \DFF_206.D ;
  wire \DFF_206.Q ;
  wire \DFF_207.CK ;
  wire \DFF_207.D ;
  wire \DFF_207.Q ;
  wire \DFF_208.CK ;
  wire \DFF_208.D ;
  wire \DFF_208.Q ;
  wire \DFF_209.CK ;
  wire \DFF_209.D ;
  wire \DFF_209.Q ;
  wire \DFF_21.CK ;
  wire \DFF_21.D ;
  wire \DFF_21.Q ;
  wire \DFF_210.CK ;
  wire \DFF_210.D ;
  wire \DFF_210.Q ;
  wire \DFF_211.CK ;
  wire \DFF_211.D ;
  wire \DFF_211.Q ;
  wire \DFF_212.CK ;
  wire \DFF_212.D ;
  wire \DFF_212.Q ;
  wire \DFF_213.CK ;
  wire \DFF_213.D ;
  wire \DFF_213.Q ;
  wire \DFF_214.CK ;
  wire \DFF_214.D ;
  wire \DFF_214.Q ;
  wire \DFF_215.CK ;
  wire \DFF_215.D ;
  wire \DFF_215.Q ;
  wire \DFF_216.CK ;
  wire \DFF_216.D ;
  wire \DFF_216.Q ;
  wire \DFF_217.CK ;
  wire \DFF_217.D ;
  wire \DFF_217.Q ;
  wire \DFF_218.CK ;
  wire \DFF_218.D ;
  wire \DFF_218.Q ;
  wire \DFF_219.CK ;
  wire \DFF_219.D ;
  wire \DFF_219.Q ;
  wire \DFF_22.CK ;
  wire \DFF_22.D ;
  wire \DFF_22.Q ;
  wire \DFF_220.CK ;
  wire \DFF_220.D ;
  wire \DFF_220.Q ;
  wire \DFF_221.CK ;
  wire \DFF_221.D ;
  wire \DFF_221.Q ;
  wire \DFF_222.CK ;
  wire \DFF_222.D ;
  wire \DFF_222.Q ;
  wire \DFF_223.CK ;
  wire \DFF_223.D ;
  wire \DFF_223.Q ;
  wire \DFF_224.CK ;
  wire \DFF_224.D ;
  wire \DFF_224.Q ;
  wire \DFF_225.CK ;
  wire \DFF_225.D ;
  wire \DFF_225.Q ;
  wire \DFF_226.CK ;
  wire \DFF_226.D ;
  wire \DFF_226.Q ;
  wire \DFF_227.CK ;
  wire \DFF_227.D ;
  wire \DFF_227.Q ;
  wire \DFF_228.CK ;
  wire \DFF_228.D ;
  wire \DFF_228.Q ;
  wire \DFF_229.CK ;
  wire \DFF_229.D ;
  wire \DFF_229.Q ;
  wire \DFF_23.CK ;
  wire \DFF_23.D ;
  wire \DFF_23.Q ;
  wire \DFF_230.CK ;
  wire \DFF_230.D ;
  wire \DFF_230.Q ;
  wire \DFF_231.CK ;
  wire \DFF_231.D ;
  wire \DFF_231.Q ;
  wire \DFF_232.CK ;
  wire \DFF_232.D ;
  wire \DFF_232.Q ;
  wire \DFF_233.CK ;
  wire \DFF_233.D ;
  wire \DFF_233.Q ;
  wire \DFF_234.CK ;
  wire \DFF_234.D ;
  wire \DFF_234.Q ;
  wire \DFF_235.CK ;
  wire \DFF_235.D ;
  wire \DFF_235.Q ;
  wire \DFF_236.CK ;
  wire \DFF_236.D ;
  wire \DFF_236.Q ;
  wire \DFF_237.CK ;
  wire \DFF_237.D ;
  wire \DFF_237.Q ;
  wire \DFF_238.CK ;
  wire \DFF_238.D ;
  wire \DFF_238.Q ;
  wire \DFF_239.CK ;
  wire \DFF_239.D ;
  wire \DFF_239.Q ;
  wire \DFF_24.CK ;
  wire \DFF_24.D ;
  wire \DFF_24.Q ;
  wire \DFF_240.CK ;
  wire \DFF_240.D ;
  wire \DFF_240.Q ;
  wire \DFF_241.CK ;
  wire \DFF_241.D ;
  wire \DFF_241.Q ;
  wire \DFF_242.CK ;
  wire \DFF_242.D ;
  wire \DFF_242.Q ;
  wire \DFF_243.CK ;
  wire \DFF_243.D ;
  wire \DFF_243.Q ;
  wire \DFF_244.CK ;
  wire \DFF_244.D ;
  wire \DFF_244.Q ;
  wire \DFF_245.CK ;
  wire \DFF_245.D ;
  wire \DFF_245.Q ;
  wire \DFF_246.CK ;
  wire \DFF_246.D ;
  wire \DFF_246.Q ;
  wire \DFF_247.CK ;
  wire \DFF_247.D ;
  wire \DFF_247.Q ;
  wire \DFF_248.CK ;
  wire \DFF_248.D ;
  wire \DFF_248.Q ;
  wire \DFF_249.CK ;
  wire \DFF_249.D ;
  wire \DFF_249.Q ;
  wire \DFF_25.CK ;
  wire \DFF_25.D ;
  wire \DFF_25.Q ;
  wire \DFF_250.CK ;
  wire \DFF_250.D ;
  wire \DFF_250.Q ;
  wire \DFF_251.CK ;
  wire \DFF_251.D ;
  wire \DFF_251.Q ;
  wire \DFF_252.CK ;
  wire \DFF_252.D ;
  wire \DFF_252.Q ;
  wire \DFF_253.CK ;
  wire \DFF_253.D ;
  wire \DFF_253.Q ;
  wire \DFF_254.CK ;
  wire \DFF_254.D ;
  wire \DFF_254.Q ;
  wire \DFF_255.CK ;
  wire \DFF_255.D ;
  wire \DFF_255.Q ;
  wire \DFF_256.CK ;
  wire \DFF_256.D ;
  wire \DFF_256.Q ;
  wire \DFF_257.CK ;
  wire \DFF_257.D ;
  wire \DFF_257.Q ;
  wire \DFF_258.CK ;
  wire \DFF_258.D ;
  wire \DFF_258.Q ;
  wire \DFF_259.CK ;
  wire \DFF_259.D ;
  wire \DFF_259.Q ;
  wire \DFF_26.CK ;
  wire \DFF_26.D ;
  wire \DFF_26.Q ;
  wire \DFF_260.CK ;
  wire \DFF_260.D ;
  wire \DFF_260.Q ;
  wire \DFF_261.CK ;
  wire \DFF_261.D ;
  wire \DFF_261.Q ;
  wire \DFF_262.CK ;
  wire \DFF_263.CK ;
  wire \DFF_263.D ;
  wire \DFF_263.Q ;
  wire \DFF_264.CK ;
  wire \DFF_264.D ;
  wire \DFF_264.Q ;
  wire \DFF_265.CK ;
  wire \DFF_265.D ;
  wire \DFF_265.Q ;
  wire \DFF_266.CK ;
  wire \DFF_266.D ;
  wire \DFF_266.Q ;
  wire \DFF_267.CK ;
  wire \DFF_267.D ;
  wire \DFF_267.Q ;
  wire \DFF_268.CK ;
  wire \DFF_268.D ;
  wire \DFF_268.Q ;
  wire \DFF_269.CK ;
  wire \DFF_269.D ;
  wire \DFF_269.Q ;
  wire \DFF_27.CK ;
  wire \DFF_27.D ;
  wire \DFF_27.Q ;
  wire \DFF_270.CK ;
  wire \DFF_270.D ;
  wire \DFF_270.Q ;
  wire \DFF_271.CK ;
  wire \DFF_271.D ;
  wire \DFF_271.Q ;
  wire \DFF_272.CK ;
  wire \DFF_272.D ;
  wire \DFF_272.Q ;
  wire \DFF_273.CK ;
  wire \DFF_273.D ;
  wire \DFF_273.Q ;
  wire \DFF_274.CK ;
  wire \DFF_274.D ;
  wire \DFF_274.Q ;
  wire \DFF_275.CK ;
  wire \DFF_275.D ;
  wire \DFF_275.Q ;
  wire \DFF_276.CK ;
  wire \DFF_276.D ;
  wire \DFF_276.Q ;
  wire \DFF_277.CK ;
  wire \DFF_277.D ;
  wire \DFF_277.Q ;
  wire \DFF_278.CK ;
  wire \DFF_278.D ;
  wire \DFF_278.Q ;
  wire \DFF_279.CK ;
  wire \DFF_279.D ;
  wire \DFF_279.Q ;
  wire \DFF_28.CK ;
  wire \DFF_28.D ;
  wire \DFF_28.Q ;
  wire \DFF_280.CK ;
  wire \DFF_280.D ;
  wire \DFF_280.Q ;
  wire \DFF_281.CK ;
  wire \DFF_281.D ;
  wire \DFF_281.Q ;
  wire \DFF_282.CK ;
  wire \DFF_282.D ;
  wire \DFF_282.Q ;
  wire \DFF_283.CK ;
  wire \DFF_283.D ;
  wire \DFF_283.Q ;
  wire \DFF_284.CK ;
  wire \DFF_284.D ;
  wire \DFF_284.Q ;
  wire \DFF_285.CK ;
  wire \DFF_285.D ;
  wire \DFF_285.Q ;
  wire \DFF_286.CK ;
  wire \DFF_286.D ;
  wire \DFF_286.Q ;
  wire \DFF_287.CK ;
  wire \DFF_287.D ;
  wire \DFF_287.Q ;
  wire \DFF_288.CK ;
  wire \DFF_288.D ;
  wire \DFF_288.Q ;
  wire \DFF_289.CK ;
  wire \DFF_289.D ;
  wire \DFF_289.Q ;
  wire \DFF_29.CK ;
  wire \DFF_29.D ;
  wire \DFF_29.Q ;
  wire \DFF_290.CK ;
  wire \DFF_290.D ;
  wire \DFF_290.Q ;
  wire \DFF_291.CK ;
  wire \DFF_291.D ;
  wire \DFF_291.Q ;
  wire \DFF_292.CK ;
  wire \DFF_292.D ;
  wire \DFF_292.Q ;
  wire \DFF_293.CK ;
  wire \DFF_293.D ;
  wire \DFF_293.Q ;
  wire \DFF_294.CK ;
  wire \DFF_294.D ;
  wire \DFF_294.Q ;
  wire \DFF_295.CK ;
  wire \DFF_295.D ;
  wire \DFF_295.Q ;
  wire \DFF_296.CK ;
  wire \DFF_296.D ;
  wire \DFF_296.Q ;
  wire \DFF_297.CK ;
  wire \DFF_297.D ;
  wire \DFF_297.Q ;
  wire \DFF_298.CK ;
  wire \DFF_298.D ;
  wire \DFF_298.Q ;
  wire \DFF_299.CK ;
  wire \DFF_299.D ;
  wire \DFF_299.Q ;
  wire \DFF_3.CK ;
  wire \DFF_3.D ;
  wire \DFF_3.Q ;
  wire \DFF_30.CK ;
  wire \DFF_30.D ;
  wire \DFF_30.Q ;
  wire \DFF_300.CK ;
  wire \DFF_300.D ;
  wire \DFF_300.Q ;
  wire \DFF_301.CK ;
  wire \DFF_301.D ;
  wire \DFF_301.Q ;
  wire \DFF_302.CK ;
  wire \DFF_302.D ;
  wire \DFF_302.Q ;
  wire \DFF_303.CK ;
  wire \DFF_303.D ;
  wire \DFF_303.Q ;
  wire \DFF_304.CK ;
  wire \DFF_304.D ;
  wire \DFF_304.Q ;
  wire \DFF_305.CK ;
  wire \DFF_305.D ;
  wire \DFF_305.Q ;
  wire \DFF_306.CK ;
  wire \DFF_306.D ;
  wire \DFF_306.Q ;
  wire \DFF_307.CK ;
  wire \DFF_307.D ;
  wire \DFF_307.Q ;
  wire \DFF_308.CK ;
  wire \DFF_308.D ;
  wire \DFF_308.Q ;
  wire \DFF_309.CK ;
  wire \DFF_309.D ;
  wire \DFF_309.Q ;
  wire \DFF_31.CK ;
  wire \DFF_31.D ;
  wire \DFF_31.Q ;
  wire \DFF_310.CK ;
  wire \DFF_310.D ;
  wire \DFF_310.Q ;
  wire \DFF_311.CK ;
  wire \DFF_311.D ;
  wire \DFF_311.Q ;
  wire \DFF_312.CK ;
  wire \DFF_312.D ;
  wire \DFF_312.Q ;
  wire \DFF_313.CK ;
  wire \DFF_313.D ;
  wire \DFF_313.Q ;
  wire \DFF_314.CK ;
  wire \DFF_314.D ;
  wire \DFF_314.Q ;
  wire \DFF_315.CK ;
  wire \DFF_315.D ;
  wire \DFF_315.Q ;
  wire \DFF_316.CK ;
  wire \DFF_316.D ;
  wire \DFF_316.Q ;
  wire \DFF_317.CK ;
  wire \DFF_317.D ;
  wire \DFF_317.Q ;
  wire \DFF_318.CK ;
  wire \DFF_318.D ;
  wire \DFF_318.Q ;
  wire \DFF_319.CK ;
  wire \DFF_319.D ;
  wire \DFF_319.Q ;
  wire \DFF_32.CK ;
  wire \DFF_32.D ;
  wire \DFF_32.Q ;
  wire \DFF_320.CK ;
  wire \DFF_320.D ;
  wire \DFF_320.Q ;
  wire \DFF_321.CK ;
  wire \DFF_321.D ;
  wire \DFF_321.Q ;
  wire \DFF_322.CK ;
  wire \DFF_322.D ;
  wire \DFF_322.Q ;
  wire \DFF_323.CK ;
  wire \DFF_323.D ;
  wire \DFF_323.Q ;
  wire \DFF_324.CK ;
  wire \DFF_324.D ;
  wire \DFF_324.Q ;
  wire \DFF_325.CK ;
  wire \DFF_325.D ;
  wire \DFF_325.Q ;
  wire \DFF_326.CK ;
  wire \DFF_326.D ;
  wire \DFF_326.Q ;
  wire \DFF_327.CK ;
  wire \DFF_327.D ;
  wire \DFF_327.Q ;
  wire \DFF_328.CK ;
  wire \DFF_328.D ;
  wire \DFF_328.Q ;
  wire \DFF_329.CK ;
  wire \DFF_329.D ;
  wire \DFF_329.Q ;
  wire \DFF_33.CK ;
  wire \DFF_33.D ;
  wire \DFF_33.Q ;
  wire \DFF_330.CK ;
  wire \DFF_330.D ;
  wire \DFF_330.Q ;
  wire \DFF_331.CK ;
  wire \DFF_331.D ;
  wire \DFF_331.Q ;
  wire \DFF_332.CK ;
  wire \DFF_332.D ;
  wire \DFF_332.Q ;
  wire \DFF_333.CK ;
  wire \DFF_333.D ;
  wire \DFF_333.Q ;
  wire \DFF_334.CK ;
  wire \DFF_334.D ;
  wire \DFF_334.Q ;
  wire \DFF_335.CK ;
  wire \DFF_335.D ;
  wire \DFF_335.Q ;
  wire \DFF_336.CK ;
  wire \DFF_336.D ;
  wire \DFF_336.Q ;
  wire \DFF_337.CK ;
  wire \DFF_337.D ;
  wire \DFF_337.Q ;
  wire \DFF_338.CK ;
  wire \DFF_338.D ;
  wire \DFF_338.Q ;
  wire \DFF_339.CK ;
  wire \DFF_339.D ;
  wire \DFF_339.Q ;
  wire \DFF_34.CK ;
  wire \DFF_34.D ;
  wire \DFF_34.Q ;
  wire \DFF_340.CK ;
  wire \DFF_340.D ;
  wire \DFF_340.Q ;
  wire \DFF_341.CK ;
  wire \DFF_341.D ;
  wire \DFF_341.Q ;
  wire \DFF_342.CK ;
  wire \DFF_342.D ;
  wire \DFF_342.Q ;
  wire \DFF_343.CK ;
  wire \DFF_343.D ;
  wire \DFF_343.Q ;
  wire \DFF_344.CK ;
  wire \DFF_344.D ;
  wire \DFF_344.Q ;
  wire \DFF_345.CK ;
  wire \DFF_345.D ;
  wire \DFF_345.Q ;
  wire \DFF_346.CK ;
  wire \DFF_346.D ;
  wire \DFF_346.Q ;
  wire \DFF_347.CK ;
  wire \DFF_347.D ;
  wire \DFF_347.Q ;
  wire \DFF_348.CK ;
  wire \DFF_348.D ;
  wire \DFF_348.Q ;
  wire \DFF_349.CK ;
  wire \DFF_349.D ;
  wire \DFF_349.Q ;
  wire \DFF_35.CK ;
  wire \DFF_35.D ;
  wire \DFF_35.Q ;
  wire \DFF_350.CK ;
  wire \DFF_350.D ;
  wire \DFF_350.Q ;
  wire \DFF_351.CK ;
  wire \DFF_351.D ;
  wire \DFF_351.Q ;
  wire \DFF_352.CK ;
  wire \DFF_352.D ;
  wire \DFF_352.Q ;
  wire \DFF_353.CK ;
  wire \DFF_353.D ;
  wire \DFF_353.Q ;
  wire \DFF_354.CK ;
  wire \DFF_354.D ;
  wire \DFF_354.Q ;
  wire \DFF_355.CK ;
  wire \DFF_355.D ;
  wire \DFF_355.Q ;
  wire \DFF_356.CK ;
  wire \DFF_356.D ;
  wire \DFF_356.Q ;
  wire \DFF_357.CK ;
  wire \DFF_357.D ;
  wire \DFF_357.Q ;
  wire \DFF_358.CK ;
  wire \DFF_358.D ;
  wire \DFF_358.Q ;
  wire \DFF_359.CK ;
  wire \DFF_359.D ;
  wire \DFF_359.Q ;
  wire \DFF_36.CK ;
  wire \DFF_36.D ;
  wire \DFF_36.Q ;
  wire \DFF_360.CK ;
  wire \DFF_360.D ;
  wire \DFF_360.Q ;
  wire \DFF_361.CK ;
  wire \DFF_361.D ;
  wire \DFF_361.Q ;
  wire \DFF_362.CK ;
  wire \DFF_362.D ;
  wire \DFF_362.Q ;
  wire \DFF_363.CK ;
  wire \DFF_363.D ;
  wire \DFF_363.Q ;
  wire \DFF_364.CK ;
  wire \DFF_364.D ;
  wire \DFF_364.Q ;
  wire \DFF_365.CK ;
  wire \DFF_365.D ;
  wire \DFF_365.Q ;
  wire \DFF_366.CK ;
  wire \DFF_366.D ;
  wire \DFF_366.Q ;
  wire \DFF_367.CK ;
  wire \DFF_367.D ;
  wire \DFF_367.Q ;
  wire \DFF_368.CK ;
  wire \DFF_368.D ;
  wire \DFF_368.Q ;
  wire \DFF_369.CK ;
  wire \DFF_369.D ;
  wire \DFF_369.Q ;
  wire \DFF_37.CK ;
  wire \DFF_37.D ;
  wire \DFF_37.Q ;
  wire \DFF_370.CK ;
  wire \DFF_370.D ;
  wire \DFF_370.Q ;
  wire \DFF_371.CK ;
  wire \DFF_371.D ;
  wire \DFF_371.Q ;
  wire \DFF_372.CK ;
  wire \DFF_372.D ;
  wire \DFF_372.Q ;
  wire \DFF_373.CK ;
  wire \DFF_373.D ;
  wire \DFF_373.Q ;
  wire \DFF_374.CK ;
  wire \DFF_374.D ;
  wire \DFF_374.Q ;
  wire \DFF_375.CK ;
  wire \DFF_375.D ;
  wire \DFF_375.Q ;
  wire \DFF_376.CK ;
  wire \DFF_376.D ;
  wire \DFF_376.Q ;
  wire \DFF_377.CK ;
  wire \DFF_377.D ;
  wire \DFF_377.Q ;
  wire \DFF_378.CK ;
  wire \DFF_378.D ;
  wire \DFF_378.Q ;
  wire \DFF_379.CK ;
  wire \DFF_379.D ;
  wire \DFF_379.Q ;
  wire \DFF_38.CK ;
  wire \DFF_38.D ;
  wire \DFF_38.Q ;
  wire \DFF_380.CK ;
  wire \DFF_380.D ;
  wire \DFF_380.Q ;
  wire \DFF_381.CK ;
  wire \DFF_381.D ;
  wire \DFF_381.Q ;
  wire \DFF_382.CK ;
  wire \DFF_382.D ;
  wire \DFF_382.Q ;
  wire \DFF_383.CK ;
  wire \DFF_383.D ;
  wire \DFF_383.Q ;
  wire \DFF_384.CK ;
  wire \DFF_384.D ;
  wire \DFF_384.Q ;
  wire \DFF_385.CK ;
  wire \DFF_385.D ;
  wire \DFF_385.Q ;
  wire \DFF_386.CK ;
  wire \DFF_386.D ;
  wire \DFF_386.Q ;
  wire \DFF_387.CK ;
  wire \DFF_387.D ;
  wire \DFF_387.Q ;
  wire \DFF_388.CK ;
  wire \DFF_388.D ;
  wire \DFF_388.Q ;
  wire \DFF_389.CK ;
  wire \DFF_389.D ;
  wire \DFF_389.Q ;
  wire \DFF_39.CK ;
  wire \DFF_39.D ;
  wire \DFF_39.Q ;
  wire \DFF_390.CK ;
  wire \DFF_390.D ;
  wire \DFF_390.Q ;
  wire \DFF_391.CK ;
  wire \DFF_391.D ;
  wire \DFF_391.Q ;
  wire \DFF_392.CK ;
  wire \DFF_392.D ;
  wire \DFF_392.Q ;
  wire \DFF_393.CK ;
  wire \DFF_393.D ;
  wire \DFF_393.Q ;
  wire \DFF_394.CK ;
  wire \DFF_394.D ;
  wire \DFF_394.Q ;
  wire \DFF_395.CK ;
  wire \DFF_395.D ;
  wire \DFF_395.Q ;
  wire \DFF_396.CK ;
  wire \DFF_396.D ;
  wire \DFF_396.Q ;
  wire \DFF_397.CK ;
  wire \DFF_397.D ;
  wire \DFF_397.Q ;
  wire \DFF_398.CK ;
  wire \DFF_398.D ;
  wire \DFF_398.Q ;
  wire \DFF_399.CK ;
  wire \DFF_399.D ;
  wire \DFF_399.Q ;
  wire \DFF_4.CK ;
  wire \DFF_4.D ;
  wire \DFF_4.Q ;
  wire \DFF_40.CK ;
  wire \DFF_40.D ;
  wire \DFF_40.Q ;
  wire \DFF_400.CK ;
  wire \DFF_400.D ;
  wire \DFF_400.Q ;
  wire \DFF_401.CK ;
  wire \DFF_401.D ;
  wire \DFF_401.Q ;
  wire \DFF_402.CK ;
  wire \DFF_402.D ;
  wire \DFF_402.Q ;
  wire \DFF_403.CK ;
  wire \DFF_403.D ;
  wire \DFF_403.Q ;
  wire \DFF_404.CK ;
  wire \DFF_404.D ;
  wire \DFF_404.Q ;
  wire \DFF_405.CK ;
  wire \DFF_405.D ;
  wire \DFF_405.Q ;
  wire \DFF_406.CK ;
  wire \DFF_406.D ;
  wire \DFF_406.Q ;
  wire \DFF_407.CK ;
  wire \DFF_407.D ;
  wire \DFF_407.Q ;
  wire \DFF_408.CK ;
  wire \DFF_408.D ;
  wire \DFF_408.Q ;
  wire \DFF_409.CK ;
  wire \DFF_409.D ;
  wire \DFF_409.Q ;
  wire \DFF_41.CK ;
  wire \DFF_41.D ;
  wire \DFF_41.Q ;
  wire \DFF_410.CK ;
  wire \DFF_410.D ;
  wire \DFF_410.Q ;
  wire \DFF_411.CK ;
  wire \DFF_411.D ;
  wire \DFF_411.Q ;
  wire \DFF_412.CK ;
  wire \DFF_412.D ;
  wire \DFF_412.Q ;
  wire \DFF_413.CK ;
  wire \DFF_413.D ;
  wire \DFF_413.Q ;
  wire \DFF_414.CK ;
  wire \DFF_414.D ;
  wire \DFF_414.Q ;
  wire \DFF_415.CK ;
  wire \DFF_415.D ;
  wire \DFF_415.Q ;
  wire \DFF_416.CK ;
  wire \DFF_416.D ;
  wire \DFF_416.Q ;
  wire \DFF_417.CK ;
  wire \DFF_417.D ;
  wire \DFF_417.Q ;
  wire \DFF_418.CK ;
  wire \DFF_418.D ;
  wire \DFF_418.Q ;
  wire \DFF_419.CK ;
  wire \DFF_419.D ;
  wire \DFF_419.Q ;
  wire \DFF_42.CK ;
  wire \DFF_42.D ;
  wire \DFF_42.Q ;
  wire \DFF_420.CK ;
  wire \DFF_420.D ;
  wire \DFF_420.Q ;
  wire \DFF_421.CK ;
  wire \DFF_421.D ;
  wire \DFF_421.Q ;
  wire \DFF_422.CK ;
  wire \DFF_422.D ;
  wire \DFF_422.Q ;
  wire \DFF_423.CK ;
  wire \DFF_423.D ;
  wire \DFF_423.Q ;
  wire \DFF_424.CK ;
  wire \DFF_424.D ;
  wire \DFF_424.Q ;
  wire \DFF_425.CK ;
  wire \DFF_425.D ;
  wire \DFF_425.Q ;
  wire \DFF_426.CK ;
  wire \DFF_426.D ;
  wire \DFF_426.Q ;
  wire \DFF_427.CK ;
  wire \DFF_427.D ;
  wire \DFF_427.Q ;
  wire \DFF_428.CK ;
  wire \DFF_428.D ;
  wire \DFF_428.Q ;
  wire \DFF_429.CK ;
  wire \DFF_429.D ;
  wire \DFF_429.Q ;
  wire \DFF_43.CK ;
  wire \DFF_43.D ;
  wire \DFF_43.Q ;
  wire \DFF_430.CK ;
  wire \DFF_430.D ;
  wire \DFF_430.Q ;
  wire \DFF_431.CK ;
  wire \DFF_431.D ;
  wire \DFF_431.Q ;
  wire \DFF_432.CK ;
  wire \DFF_432.D ;
  wire \DFF_432.Q ;
  wire \DFF_433.CK ;
  wire \DFF_433.D ;
  wire \DFF_433.Q ;
  wire \DFF_434.CK ;
  wire \DFF_434.D ;
  wire \DFF_434.Q ;
  wire \DFF_435.CK ;
  wire \DFF_435.D ;
  wire \DFF_435.Q ;
  wire \DFF_436.CK ;
  wire \DFF_436.D ;
  wire \DFF_436.Q ;
  wire \DFF_437.CK ;
  wire \DFF_437.D ;
  wire \DFF_437.Q ;
  wire \DFF_438.CK ;
  wire \DFF_438.D ;
  wire \DFF_438.Q ;
  wire \DFF_439.CK ;
  wire \DFF_439.D ;
  wire \DFF_439.Q ;
  wire \DFF_44.CK ;
  wire \DFF_44.D ;
  wire \DFF_44.Q ;
  wire \DFF_440.CK ;
  wire \DFF_440.D ;
  wire \DFF_440.Q ;
  wire \DFF_441.CK ;
  wire \DFF_441.D ;
  wire \DFF_441.Q ;
  wire \DFF_442.CK ;
  wire \DFF_442.D ;
  wire \DFF_442.Q ;
  wire \DFF_443.CK ;
  wire \DFF_443.D ;
  wire \DFF_443.Q ;
  wire \DFF_444.CK ;
  wire \DFF_444.D ;
  wire \DFF_444.Q ;
  wire \DFF_445.CK ;
  wire \DFF_445.D ;
  wire \DFF_445.Q ;
  wire \DFF_446.CK ;
  wire \DFF_446.D ;
  wire \DFF_446.Q ;
  wire \DFF_447.CK ;
  wire \DFF_447.D ;
  wire \DFF_447.Q ;
  wire \DFF_448.CK ;
  wire \DFF_448.D ;
  wire \DFF_448.Q ;
  wire \DFF_449.CK ;
  wire \DFF_449.D ;
  wire \DFF_449.Q ;
  wire \DFF_45.CK ;
  wire \DFF_45.D ;
  wire \DFF_45.Q ;
  wire \DFF_450.CK ;
  wire \DFF_450.D ;
  wire \DFF_450.Q ;
  wire \DFF_451.CK ;
  wire \DFF_451.D ;
  wire \DFF_451.Q ;
  wire \DFF_452.CK ;
  wire \DFF_452.D ;
  wire \DFF_452.Q ;
  wire \DFF_453.CK ;
  wire \DFF_453.D ;
  wire \DFF_453.Q ;
  wire \DFF_454.CK ;
  wire \DFF_454.D ;
  wire \DFF_454.Q ;
  wire \DFF_455.CK ;
  wire \DFF_455.D ;
  wire \DFF_455.Q ;
  wire \DFF_456.CK ;
  wire \DFF_456.D ;
  wire \DFF_456.Q ;
  wire \DFF_457.CK ;
  wire \DFF_457.D ;
  wire \DFF_457.Q ;
  wire \DFF_458.CK ;
  wire \DFF_458.D ;
  wire \DFF_458.Q ;
  wire \DFF_459.CK ;
  wire \DFF_459.D ;
  wire \DFF_459.Q ;
  wire \DFF_46.CK ;
  wire \DFF_46.D ;
  wire \DFF_46.Q ;
  wire \DFF_460.CK ;
  wire \DFF_460.D ;
  wire \DFF_460.Q ;
  wire \DFF_461.CK ;
  wire \DFF_461.D ;
  wire \DFF_461.Q ;
  wire \DFF_462.CK ;
  wire \DFF_462.D ;
  wire \DFF_462.Q ;
  wire \DFF_463.CK ;
  wire \DFF_463.D ;
  wire \DFF_463.Q ;
  wire \DFF_464.CK ;
  wire \DFF_464.D ;
  wire \DFF_464.Q ;
  wire \DFF_465.CK ;
  wire \DFF_465.D ;
  wire \DFF_465.Q ;
  wire \DFF_466.CK ;
  wire \DFF_466.D ;
  wire \DFF_466.Q ;
  wire \DFF_467.CK ;
  wire \DFF_467.D ;
  wire \DFF_467.Q ;
  wire \DFF_468.CK ;
  wire \DFF_468.D ;
  wire \DFF_468.Q ;
  wire \DFF_469.CK ;
  wire \DFF_469.D ;
  wire \DFF_469.Q ;
  wire \DFF_47.CK ;
  wire \DFF_47.D ;
  wire \DFF_47.Q ;
  wire \DFF_470.CK ;
  wire \DFF_470.D ;
  wire \DFF_470.Q ;
  wire \DFF_471.CK ;
  wire \DFF_471.D ;
  wire \DFF_471.Q ;
  wire \DFF_472.CK ;
  wire \DFF_472.D ;
  wire \DFF_472.Q ;
  wire \DFF_473.CK ;
  wire \DFF_473.D ;
  wire \DFF_473.Q ;
  wire \DFF_474.CK ;
  wire \DFF_474.D ;
  wire \DFF_474.Q ;
  wire \DFF_475.CK ;
  wire \DFF_475.D ;
  wire \DFF_475.Q ;
  wire \DFF_476.CK ;
  wire \DFF_476.D ;
  wire \DFF_476.Q ;
  wire \DFF_477.CK ;
  wire \DFF_477.D ;
  wire \DFF_477.Q ;
  wire \DFF_478.CK ;
  wire \DFF_478.D ;
  wire \DFF_478.Q ;
  wire \DFF_479.CK ;
  wire \DFF_479.D ;
  wire \DFF_479.Q ;
  wire \DFF_48.CK ;
  wire \DFF_48.D ;
  wire \DFF_48.Q ;
  wire \DFF_480.CK ;
  wire \DFF_480.D ;
  wire \DFF_480.Q ;
  wire \DFF_481.CK ;
  wire \DFF_481.D ;
  wire \DFF_481.Q ;
  wire \DFF_482.CK ;
  wire \DFF_482.D ;
  wire \DFF_482.Q ;
  wire \DFF_483.CK ;
  wire \DFF_483.D ;
  wire \DFF_483.Q ;
  wire \DFF_484.CK ;
  wire \DFF_484.D ;
  wire \DFF_484.Q ;
  wire \DFF_485.CK ;
  wire \DFF_485.D ;
  wire \DFF_485.Q ;
  wire \DFF_486.CK ;
  wire \DFF_486.D ;
  wire \DFF_486.Q ;
  wire \DFF_487.CK ;
  wire \DFF_487.D ;
  wire \DFF_487.Q ;
  wire \DFF_488.CK ;
  wire \DFF_488.D ;
  wire \DFF_488.Q ;
  wire \DFF_489.CK ;
  wire \DFF_489.D ;
  wire \DFF_489.Q ;
  wire \DFF_49.CK ;
  wire \DFF_49.D ;
  wire \DFF_49.Q ;
  wire \DFF_490.CK ;
  wire \DFF_490.D ;
  wire \DFF_490.Q ;
  wire \DFF_491.CK ;
  wire \DFF_491.D ;
  wire \DFF_491.Q ;
  wire \DFF_492.CK ;
  wire \DFF_492.D ;
  wire \DFF_492.Q ;
  wire \DFF_493.CK ;
  wire \DFF_493.D ;
  wire \DFF_493.Q ;
  wire \DFF_494.CK ;
  wire \DFF_494.D ;
  wire \DFF_494.Q ;
  wire \DFF_495.CK ;
  wire \DFF_495.D ;
  wire \DFF_495.Q ;
  wire \DFF_496.CK ;
  wire \DFF_496.D ;
  wire \DFF_496.Q ;
  wire \DFF_497.CK ;
  wire \DFF_497.D ;
  wire \DFF_497.Q ;
  wire \DFF_498.CK ;
  wire \DFF_498.D ;
  wire \DFF_498.Q ;
  wire \DFF_499.CK ;
  wire \DFF_499.D ;
  wire \DFF_499.Q ;
  wire \DFF_5.CK ;
  wire \DFF_5.D ;
  wire \DFF_5.Q ;
  wire \DFF_50.CK ;
  wire \DFF_50.D ;
  wire \DFF_50.Q ;
  wire \DFF_500.CK ;
  wire \DFF_500.D ;
  wire \DFF_500.Q ;
  wire \DFF_501.CK ;
  wire \DFF_501.D ;
  wire \DFF_501.Q ;
  wire \DFF_502.CK ;
  wire \DFF_502.D ;
  wire \DFF_502.Q ;
  wire \DFF_503.CK ;
  wire \DFF_503.D ;
  wire \DFF_503.Q ;
  wire \DFF_504.CK ;
  wire \DFF_504.D ;
  wire \DFF_504.Q ;
  wire \DFF_505.CK ;
  wire \DFF_505.D ;
  wire \DFF_505.Q ;
  wire \DFF_506.CK ;
  wire \DFF_506.D ;
  wire \DFF_506.Q ;
  wire \DFF_507.CK ;
  wire \DFF_507.D ;
  wire \DFF_507.Q ;
  wire \DFF_508.CK ;
  wire \DFF_508.D ;
  wire \DFF_508.Q ;
  wire \DFF_509.CK ;
  wire \DFF_509.D ;
  wire \DFF_509.Q ;
  wire \DFF_51.CK ;
  wire \DFF_51.D ;
  wire \DFF_51.Q ;
  wire \DFF_510.CK ;
  wire \DFF_510.D ;
  wire \DFF_510.Q ;
  wire \DFF_511.CK ;
  wire \DFF_511.D ;
  wire \DFF_511.Q ;
  wire \DFF_512.CK ;
  wire \DFF_512.D ;
  wire \DFF_512.Q ;
  wire \DFF_513.CK ;
  wire \DFF_513.D ;
  wire \DFF_513.Q ;
  wire \DFF_514.CK ;
  wire \DFF_514.D ;
  wire \DFF_514.Q ;
  wire \DFF_515.CK ;
  wire \DFF_515.D ;
  wire \DFF_515.Q ;
  wire \DFF_516.CK ;
  wire \DFF_516.D ;
  wire \DFF_516.Q ;
  wire \DFF_517.CK ;
  wire \DFF_517.D ;
  wire \DFF_517.Q ;
  wire \DFF_518.CK ;
  wire \DFF_518.D ;
  wire \DFF_518.Q ;
  wire \DFF_519.CK ;
  wire \DFF_519.D ;
  wire \DFF_519.Q ;
  wire \DFF_52.CK ;
  wire \DFF_52.D ;
  wire \DFF_52.Q ;
  wire \DFF_520.CK ;
  wire \DFF_520.D ;
  wire \DFF_520.Q ;
  wire \DFF_521.CK ;
  wire \DFF_521.D ;
  wire \DFF_521.Q ;
  wire \DFF_522.CK ;
  wire \DFF_522.D ;
  wire \DFF_522.Q ;
  wire \DFF_523.CK ;
  wire \DFF_523.D ;
  wire \DFF_523.Q ;
  wire \DFF_524.CK ;
  wire \DFF_524.D ;
  wire \DFF_524.Q ;
  wire \DFF_525.CK ;
  wire \DFF_525.D ;
  wire \DFF_525.Q ;
  wire \DFF_526.CK ;
  wire \DFF_526.D ;
  wire \DFF_526.Q ;
  wire \DFF_527.CK ;
  wire \DFF_527.D ;
  wire \DFF_527.Q ;
  wire \DFF_528.CK ;
  wire \DFF_528.D ;
  wire \DFF_528.Q ;
  wire \DFF_529.CK ;
  wire \DFF_529.D ;
  wire \DFF_529.Q ;
  wire \DFF_53.CK ;
  wire \DFF_53.D ;
  wire \DFF_53.Q ;
  wire \DFF_530.CK ;
  wire \DFF_530.D ;
  wire \DFF_530.Q ;
  wire \DFF_531.CK ;
  wire \DFF_531.D ;
  wire \DFF_531.Q ;
  wire \DFF_532.CK ;
  wire \DFF_532.D ;
  wire \DFF_532.Q ;
  wire \DFF_533.CK ;
  wire \DFF_533.D ;
  wire \DFF_533.Q ;
  wire \DFF_534.CK ;
  wire \DFF_534.D ;
  wire \DFF_534.Q ;
  wire \DFF_535.CK ;
  wire \DFF_535.D ;
  wire \DFF_535.Q ;
  wire \DFF_536.CK ;
  wire \DFF_536.D ;
  wire \DFF_536.Q ;
  wire \DFF_537.CK ;
  wire \DFF_537.D ;
  wire \DFF_537.Q ;
  wire \DFF_538.CK ;
  wire \DFF_538.D ;
  wire \DFF_538.Q ;
  wire \DFF_539.CK ;
  wire \DFF_539.D ;
  wire \DFF_539.Q ;
  wire \DFF_54.CK ;
  wire \DFF_54.D ;
  wire \DFF_54.Q ;
  wire \DFF_540.CK ;
  wire \DFF_540.D ;
  wire \DFF_540.Q ;
  wire \DFF_541.CK ;
  wire \DFF_541.D ;
  wire \DFF_541.Q ;
  wire \DFF_542.CK ;
  wire \DFF_542.D ;
  wire \DFF_542.Q ;
  wire \DFF_543.CK ;
  wire \DFF_543.D ;
  wire \DFF_543.Q ;
  wire \DFF_544.CK ;
  wire \DFF_544.D ;
  wire \DFF_544.Q ;
  wire \DFF_545.CK ;
  wire \DFF_545.D ;
  wire \DFF_545.Q ;
  wire \DFF_546.CK ;
  wire \DFF_546.D ;
  wire \DFF_546.Q ;
  wire \DFF_547.CK ;
  wire \DFF_547.D ;
  wire \DFF_547.Q ;
  wire \DFF_548.CK ;
  wire \DFF_548.D ;
  wire \DFF_548.Q ;
  wire \DFF_549.CK ;
  wire \DFF_549.D ;
  wire \DFF_549.Q ;
  wire \DFF_55.CK ;
  wire \DFF_55.D ;
  wire \DFF_55.Q ;
  wire \DFF_550.CK ;
  wire \DFF_550.D ;
  wire \DFF_550.Q ;
  wire \DFF_551.CK ;
  wire \DFF_551.D ;
  wire \DFF_551.Q ;
  wire \DFF_552.CK ;
  wire \DFF_552.D ;
  wire \DFF_552.Q ;
  wire \DFF_553.CK ;
  wire \DFF_553.D ;
  wire \DFF_553.Q ;
  wire \DFF_554.CK ;
  wire \DFF_554.D ;
  wire \DFF_554.Q ;
  wire \DFF_555.CK ;
  wire \DFF_555.D ;
  wire \DFF_555.Q ;
  wire \DFF_556.CK ;
  wire \DFF_556.D ;
  wire \DFF_556.Q ;
  wire \DFF_557.CK ;
  wire \DFF_557.D ;
  wire \DFF_557.Q ;
  wire \DFF_558.CK ;
  wire \DFF_558.D ;
  wire \DFF_558.Q ;
  wire \DFF_559.CK ;
  wire \DFF_559.D ;
  wire \DFF_559.Q ;
  wire \DFF_56.CK ;
  wire \DFF_56.D ;
  wire \DFF_56.Q ;
  wire \DFF_560.CK ;
  wire \DFF_560.D ;
  wire \DFF_560.Q ;
  wire \DFF_561.CK ;
  wire \DFF_561.D ;
  wire \DFF_561.Q ;
  wire \DFF_562.CK ;
  wire \DFF_562.D ;
  wire \DFF_562.Q ;
  wire \DFF_563.CK ;
  wire \DFF_563.D ;
  wire \DFF_563.Q ;
  wire \DFF_564.CK ;
  wire \DFF_564.D ;
  wire \DFF_564.Q ;
  wire \DFF_565.CK ;
  wire \DFF_565.D ;
  wire \DFF_565.Q ;
  wire \DFF_566.CK ;
  wire \DFF_566.D ;
  wire \DFF_566.Q ;
  wire \DFF_567.CK ;
  wire \DFF_567.D ;
  wire \DFF_567.Q ;
  wire \DFF_568.CK ;
  wire \DFF_568.D ;
  wire \DFF_568.Q ;
  wire \DFF_569.CK ;
  wire \DFF_569.D ;
  wire \DFF_569.Q ;
  wire \DFF_57.CK ;
  wire \DFF_57.D ;
  wire \DFF_57.Q ;
  wire \DFF_570.CK ;
  wire \DFF_570.D ;
  wire \DFF_570.Q ;
  wire \DFF_571.CK ;
  wire \DFF_571.D ;
  wire \DFF_571.Q ;
  wire \DFF_572.CK ;
  wire \DFF_572.D ;
  wire \DFF_572.Q ;
  wire \DFF_573.CK ;
  wire \DFF_573.D ;
  wire \DFF_573.Q ;
  wire \DFF_574.CK ;
  wire \DFF_574.D ;
  wire \DFF_574.Q ;
  wire \DFF_575.CK ;
  wire \DFF_575.D ;
  wire \DFF_575.Q ;
  wire \DFF_576.CK ;
  wire \DFF_576.D ;
  wire \DFF_576.Q ;
  wire \DFF_577.CK ;
  wire \DFF_577.D ;
  wire \DFF_577.Q ;
  wire \DFF_578.CK ;
  wire \DFF_578.D ;
  wire \DFF_578.Q ;
  wire \DFF_579.CK ;
  wire \DFF_579.D ;
  wire \DFF_579.Q ;
  wire \DFF_58.CK ;
  wire \DFF_58.D ;
  wire \DFF_58.Q ;
  wire \DFF_580.CK ;
  wire \DFF_580.D ;
  wire \DFF_580.Q ;
  wire \DFF_581.CK ;
  wire \DFF_581.D ;
  wire \DFF_581.Q ;
  wire \DFF_582.CK ;
  wire \DFF_582.D ;
  wire \DFF_582.Q ;
  wire \DFF_583.CK ;
  wire \DFF_583.D ;
  wire \DFF_583.Q ;
  wire \DFF_584.CK ;
  wire \DFF_584.D ;
  wire \DFF_584.Q ;
  wire \DFF_585.CK ;
  wire \DFF_585.D ;
  wire \DFF_585.Q ;
  wire \DFF_586.CK ;
  wire \DFF_586.D ;
  wire \DFF_586.Q ;
  wire \DFF_587.CK ;
  wire \DFF_587.D ;
  wire \DFF_587.Q ;
  wire \DFF_588.CK ;
  wire \DFF_588.D ;
  wire \DFF_588.Q ;
  wire \DFF_589.CK ;
  wire \DFF_589.D ;
  wire \DFF_589.Q ;
  wire \DFF_59.CK ;
  wire \DFF_59.D ;
  wire \DFF_59.Q ;
  wire \DFF_590.CK ;
  wire \DFF_590.D ;
  wire \DFF_590.Q ;
  wire \DFF_591.CK ;
  wire \DFF_591.D ;
  wire \DFF_591.Q ;
  wire \DFF_592.CK ;
  wire \DFF_592.D ;
  wire \DFF_592.Q ;
  wire \DFF_593.CK ;
  wire \DFF_593.D ;
  wire \DFF_593.Q ;
  wire \DFF_594.CK ;
  wire \DFF_594.D ;
  wire \DFF_594.Q ;
  wire \DFF_595.CK ;
  wire \DFF_595.D ;
  wire \DFF_595.Q ;
  wire \DFF_596.CK ;
  wire \DFF_596.D ;
  wire \DFF_596.Q ;
  wire \DFF_597.CK ;
  wire \DFF_597.D ;
  wire \DFF_597.Q ;
  wire \DFF_598.CK ;
  wire \DFF_598.D ;
  wire \DFF_598.Q ;
  wire \DFF_599.CK ;
  wire \DFF_599.D ;
  wire \DFF_599.Q ;
  wire \DFF_6.CK ;
  wire \DFF_6.D ;
  wire \DFF_6.Q ;
  wire \DFF_60.CK ;
  wire \DFF_60.D ;
  wire \DFF_60.Q ;
  wire \DFF_600.CK ;
  wire \DFF_600.D ;
  wire \DFF_600.Q ;
  wire \DFF_601.CK ;
  wire \DFF_601.D ;
  wire \DFF_601.Q ;
  wire \DFF_602.CK ;
  wire \DFF_602.D ;
  wire \DFF_602.Q ;
  wire \DFF_603.CK ;
  wire \DFF_603.D ;
  wire \DFF_603.Q ;
  wire \DFF_604.CK ;
  wire \DFF_604.D ;
  wire \DFF_604.Q ;
  wire \DFF_605.CK ;
  wire \DFF_605.D ;
  wire \DFF_605.Q ;
  wire \DFF_606.CK ;
  wire \DFF_606.D ;
  wire \DFF_606.Q ;
  wire \DFF_607.CK ;
  wire \DFF_607.D ;
  wire \DFF_607.Q ;
  wire \DFF_608.CK ;
  wire \DFF_608.D ;
  wire \DFF_608.Q ;
  wire \DFF_609.CK ;
  wire \DFF_609.D ;
  wire \DFF_609.Q ;
  wire \DFF_61.CK ;
  wire \DFF_61.D ;
  wire \DFF_61.Q ;
  wire \DFF_610.CK ;
  wire \DFF_610.D ;
  wire \DFF_610.Q ;
  wire \DFF_611.CK ;
  wire \DFF_611.D ;
  wire \DFF_611.Q ;
  wire \DFF_612.CK ;
  wire \DFF_612.D ;
  wire \DFF_612.Q ;
  wire \DFF_613.CK ;
  wire \DFF_613.D ;
  wire \DFF_613.Q ;
  wire \DFF_614.CK ;
  wire \DFF_614.D ;
  wire \DFF_614.Q ;
  wire \DFF_615.CK ;
  wire \DFF_615.D ;
  wire \DFF_615.Q ;
  wire \DFF_616.CK ;
  wire \DFF_616.D ;
  wire \DFF_616.Q ;
  wire \DFF_617.CK ;
  wire \DFF_617.D ;
  wire \DFF_617.Q ;
  wire \DFF_618.CK ;
  wire \DFF_618.D ;
  wire \DFF_618.Q ;
  wire \DFF_619.CK ;
  wire \DFF_619.D ;
  wire \DFF_619.Q ;
  wire \DFF_62.CK ;
  wire \DFF_62.D ;
  wire \DFF_62.Q ;
  wire \DFF_620.CK ;
  wire \DFF_620.D ;
  wire \DFF_620.Q ;
  wire \DFF_621.CK ;
  wire \DFF_621.D ;
  wire \DFF_621.Q ;
  wire \DFF_622.CK ;
  wire \DFF_622.D ;
  wire \DFF_622.Q ;
  wire \DFF_623.CK ;
  wire \DFF_623.D ;
  wire \DFF_623.Q ;
  wire \DFF_624.CK ;
  wire \DFF_624.D ;
  wire \DFF_624.Q ;
  wire \DFF_625.CK ;
  wire \DFF_625.D ;
  wire \DFF_625.Q ;
  wire \DFF_626.CK ;
  wire \DFF_626.D ;
  wire \DFF_626.Q ;
  wire \DFF_627.CK ;
  wire \DFF_627.D ;
  wire \DFF_627.Q ;
  wire \DFF_628.CK ;
  wire \DFF_628.D ;
  wire \DFF_628.Q ;
  wire \DFF_629.CK ;
  wire \DFF_629.D ;
  wire \DFF_629.Q ;
  wire \DFF_63.CK ;
  wire \DFF_63.D ;
  wire \DFF_63.Q ;
  wire \DFF_630.CK ;
  wire \DFF_630.D ;
  wire \DFF_630.Q ;
  wire \DFF_631.CK ;
  wire \DFF_631.D ;
  wire \DFF_631.Q ;
  wire \DFF_632.CK ;
  wire \DFF_632.D ;
  wire \DFF_632.Q ;
  wire \DFF_633.CK ;
  wire \DFF_633.D ;
  wire \DFF_633.Q ;
  wire \DFF_634.CK ;
  wire \DFF_634.D ;
  wire \DFF_634.Q ;
  wire \DFF_635.CK ;
  wire \DFF_635.D ;
  wire \DFF_635.Q ;
  wire \DFF_636.CK ;
  wire \DFF_636.D ;
  wire \DFF_636.Q ;
  wire \DFF_637.CK ;
  wire \DFF_637.D ;
  wire \DFF_637.Q ;
  wire \DFF_638.CK ;
  wire \DFF_638.D ;
  wire \DFF_638.Q ;
  wire \DFF_639.CK ;
  wire \DFF_639.D ;
  wire \DFF_639.Q ;
  wire \DFF_64.CK ;
  wire \DFF_64.D ;
  wire \DFF_64.Q ;
  wire \DFF_640.CK ;
  wire \DFF_640.D ;
  wire \DFF_640.Q ;
  wire \DFF_641.CK ;
  wire \DFF_641.D ;
  wire \DFF_641.Q ;
  wire \DFF_642.CK ;
  wire \DFF_642.D ;
  wire \DFF_642.Q ;
  wire \DFF_643.CK ;
  wire \DFF_643.D ;
  wire \DFF_643.Q ;
  wire \DFF_644.CK ;
  wire \DFF_644.D ;
  wire \DFF_644.Q ;
  wire \DFF_645.CK ;
  wire \DFF_645.D ;
  wire \DFF_645.Q ;
  wire \DFF_646.CK ;
  wire \DFF_646.D ;
  wire \DFF_646.Q ;
  wire \DFF_647.CK ;
  wire \DFF_647.D ;
  wire \DFF_647.Q ;
  wire \DFF_648.CK ;
  wire \DFF_648.D ;
  wire \DFF_648.Q ;
  wire \DFF_649.CK ;
  wire \DFF_649.D ;
  wire \DFF_649.Q ;
  wire \DFF_65.CK ;
  wire \DFF_65.D ;
  wire \DFF_65.Q ;
  wire \DFF_650.CK ;
  wire \DFF_650.D ;
  wire \DFF_650.Q ;
  wire \DFF_651.CK ;
  wire \DFF_651.D ;
  wire \DFF_651.Q ;
  wire \DFF_652.CK ;
  wire \DFF_652.D ;
  wire \DFF_652.Q ;
  wire \DFF_653.CK ;
  wire \DFF_653.D ;
  wire \DFF_653.Q ;
  wire \DFF_654.CK ;
  wire \DFF_654.D ;
  wire \DFF_654.Q ;
  wire \DFF_655.CK ;
  wire \DFF_655.D ;
  wire \DFF_655.Q ;
  wire \DFF_656.CK ;
  wire \DFF_656.D ;
  wire \DFF_656.Q ;
  wire \DFF_657.CK ;
  wire \DFF_657.D ;
  wire \DFF_657.Q ;
  wire \DFF_658.CK ;
  wire \DFF_658.D ;
  wire \DFF_658.Q ;
  wire \DFF_659.CK ;
  wire \DFF_659.D ;
  wire \DFF_659.Q ;
  wire \DFF_66.CK ;
  wire \DFF_66.D ;
  wire \DFF_66.Q ;
  wire \DFF_660.CK ;
  wire \DFF_660.D ;
  wire \DFF_660.Q ;
  wire \DFF_661.CK ;
  wire \DFF_661.D ;
  wire \DFF_661.Q ;
  wire \DFF_662.CK ;
  wire \DFF_662.D ;
  wire \DFF_662.Q ;
  wire \DFF_663.CK ;
  wire \DFF_663.D ;
  wire \DFF_663.Q ;
  wire \DFF_664.CK ;
  wire \DFF_664.D ;
  wire \DFF_664.Q ;
  wire \DFF_665.CK ;
  wire \DFF_665.D ;
  wire \DFF_665.Q ;
  wire \DFF_666.CK ;
  wire \DFF_666.D ;
  wire \DFF_666.Q ;
  wire \DFF_667.CK ;
  wire \DFF_667.D ;
  wire \DFF_667.Q ;
  wire \DFF_668.CK ;
  wire \DFF_668.D ;
  wire \DFF_668.Q ;
  wire \DFF_669.CK ;
  wire \DFF_669.D ;
  wire \DFF_669.Q ;
  wire \DFF_67.CK ;
  wire \DFF_67.D ;
  wire \DFF_67.Q ;
  wire \DFF_670.CK ;
  wire \DFF_670.D ;
  wire \DFF_670.Q ;
  wire \DFF_671.CK ;
  wire \DFF_671.D ;
  wire \DFF_671.Q ;
  wire \DFF_672.CK ;
  wire \DFF_672.D ;
  wire \DFF_672.Q ;
  wire \DFF_673.CK ;
  wire \DFF_673.D ;
  wire \DFF_673.Q ;
  wire \DFF_674.CK ;
  wire \DFF_674.D ;
  wire \DFF_674.Q ;
  wire \DFF_675.CK ;
  wire \DFF_675.D ;
  wire \DFF_675.Q ;
  wire \DFF_676.CK ;
  wire \DFF_676.D ;
  wire \DFF_676.Q ;
  wire \DFF_677.CK ;
  wire \DFF_677.D ;
  wire \DFF_677.Q ;
  wire \DFF_678.CK ;
  wire \DFF_678.D ;
  wire \DFF_678.Q ;
  wire \DFF_679.CK ;
  wire \DFF_679.D ;
  wire \DFF_679.Q ;
  wire \DFF_68.CK ;
  wire \DFF_68.D ;
  wire \DFF_68.Q ;
  wire \DFF_680.CK ;
  wire \DFF_680.D ;
  wire \DFF_680.Q ;
  wire \DFF_681.CK ;
  wire \DFF_681.D ;
  wire \DFF_681.Q ;
  wire \DFF_682.CK ;
  wire \DFF_682.D ;
  wire \DFF_682.Q ;
  wire \DFF_683.CK ;
  wire \DFF_683.D ;
  wire \DFF_683.Q ;
  wire \DFF_684.CK ;
  wire \DFF_684.D ;
  wire \DFF_684.Q ;
  wire \DFF_685.CK ;
  wire \DFF_685.D ;
  wire \DFF_685.Q ;
  wire \DFF_686.CK ;
  wire \DFF_686.D ;
  wire \DFF_686.Q ;
  wire \DFF_687.CK ;
  wire \DFF_687.D ;
  wire \DFF_687.Q ;
  wire \DFF_688.CK ;
  wire \DFF_688.D ;
  wire \DFF_688.Q ;
  wire \DFF_689.CK ;
  wire \DFF_689.D ;
  wire \DFF_689.Q ;
  wire \DFF_69.CK ;
  wire \DFF_69.D ;
  wire \DFF_69.Q ;
  wire \DFF_690.CK ;
  wire \DFF_690.D ;
  wire \DFF_690.Q ;
  wire \DFF_691.CK ;
  wire \DFF_691.D ;
  wire \DFF_691.Q ;
  wire \DFF_692.CK ;
  wire \DFF_692.D ;
  wire \DFF_692.Q ;
  wire \DFF_693.CK ;
  wire \DFF_693.D ;
  wire \DFF_693.Q ;
  wire \DFF_694.CK ;
  wire \DFF_694.D ;
  wire \DFF_694.Q ;
  wire \DFF_695.CK ;
  wire \DFF_695.D ;
  wire \DFF_695.Q ;
  wire \DFF_696.CK ;
  wire \DFF_696.D ;
  wire \DFF_696.Q ;
  wire \DFF_697.CK ;
  wire \DFF_697.D ;
  wire \DFF_697.Q ;
  wire \DFF_698.CK ;
  wire \DFF_698.D ;
  wire \DFF_698.Q ;
  wire \DFF_699.CK ;
  wire \DFF_699.D ;
  wire \DFF_699.Q ;
  wire \DFF_7.CK ;
  wire \DFF_7.D ;
  wire \DFF_7.Q ;
  wire \DFF_70.CK ;
  wire \DFF_70.D ;
  wire \DFF_70.Q ;
  wire \DFF_700.CK ;
  wire \DFF_700.D ;
  wire \DFF_700.Q ;
  wire \DFF_701.CK ;
  wire \DFF_701.D ;
  wire \DFF_701.Q ;
  wire \DFF_702.CK ;
  wire \DFF_702.D ;
  wire \DFF_702.Q ;
  wire \DFF_703.CK ;
  wire \DFF_703.D ;
  wire \DFF_703.Q ;
  wire \DFF_704.CK ;
  wire \DFF_704.D ;
  wire \DFF_704.Q ;
  wire \DFF_705.CK ;
  wire \DFF_705.D ;
  wire \DFF_705.Q ;
  wire \DFF_706.CK ;
  wire \DFF_706.D ;
  wire \DFF_706.Q ;
  wire \DFF_707.CK ;
  wire \DFF_707.D ;
  wire \DFF_707.Q ;
  wire \DFF_708.CK ;
  wire \DFF_708.D ;
  wire \DFF_708.Q ;
  wire \DFF_709.CK ;
  wire \DFF_709.D ;
  wire \DFF_709.Q ;
  wire \DFF_71.CK ;
  wire \DFF_71.D ;
  wire \DFF_71.Q ;
  wire \DFF_710.CK ;
  wire \DFF_710.D ;
  wire \DFF_710.Q ;
  wire \DFF_711.CK ;
  wire \DFF_711.D ;
  wire \DFF_711.Q ;
  wire \DFF_712.CK ;
  wire \DFF_712.D ;
  wire \DFF_712.Q ;
  wire \DFF_713.CK ;
  wire \DFF_713.D ;
  wire \DFF_713.Q ;
  wire \DFF_714.CK ;
  wire \DFF_714.D ;
  wire \DFF_714.Q ;
  wire \DFF_715.CK ;
  wire \DFF_715.D ;
  wire \DFF_715.Q ;
  wire \DFF_716.CK ;
  wire \DFF_716.D ;
  wire \DFF_716.Q ;
  wire \DFF_717.CK ;
  wire \DFF_717.D ;
  wire \DFF_717.Q ;
  wire \DFF_718.CK ;
  wire \DFF_718.D ;
  wire \DFF_718.Q ;
  wire \DFF_719.CK ;
  wire \DFF_719.D ;
  wire \DFF_719.Q ;
  wire \DFF_72.CK ;
  wire \DFF_72.D ;
  wire \DFF_72.Q ;
  wire \DFF_720.CK ;
  wire \DFF_720.D ;
  wire \DFF_720.Q ;
  wire \DFF_721.CK ;
  wire \DFF_721.D ;
  wire \DFF_721.Q ;
  wire \DFF_722.CK ;
  wire \DFF_722.D ;
  wire \DFF_722.Q ;
  wire \DFF_723.CK ;
  wire \DFF_723.D ;
  wire \DFF_723.Q ;
  wire \DFF_724.CK ;
  wire \DFF_724.D ;
  wire \DFF_724.Q ;
  wire \DFF_725.CK ;
  wire \DFF_725.D ;
  wire \DFF_725.Q ;
  wire \DFF_726.CK ;
  wire \DFF_726.D ;
  wire \DFF_726.Q ;
  wire \DFF_727.CK ;
  wire \DFF_727.D ;
  wire \DFF_727.Q ;
  wire \DFF_728.CK ;
  wire \DFF_728.D ;
  wire \DFF_728.Q ;
  wire \DFF_729.CK ;
  wire \DFF_729.D ;
  wire \DFF_729.Q ;
  wire \DFF_73.CK ;
  wire \DFF_73.D ;
  wire \DFF_73.Q ;
  wire \DFF_730.CK ;
  wire \DFF_730.D ;
  wire \DFF_730.Q ;
  wire \DFF_731.CK ;
  wire \DFF_731.D ;
  wire \DFF_731.Q ;
  wire \DFF_732.CK ;
  wire \DFF_732.D ;
  wire \DFF_732.Q ;
  wire \DFF_733.CK ;
  wire \DFF_733.D ;
  wire \DFF_733.Q ;
  wire \DFF_734.CK ;
  wire \DFF_734.D ;
  wire \DFF_734.Q ;
  wire \DFF_735.CK ;
  wire \DFF_735.D ;
  wire \DFF_735.Q ;
  wire \DFF_736.CK ;
  wire \DFF_736.D ;
  wire \DFF_736.Q ;
  wire \DFF_737.CK ;
  wire \DFF_737.D ;
  wire \DFF_737.Q ;
  wire \DFF_738.CK ;
  wire \DFF_738.D ;
  wire \DFF_738.Q ;
  wire \DFF_739.CK ;
  wire \DFF_739.D ;
  wire \DFF_739.Q ;
  wire \DFF_74.CK ;
  wire \DFF_74.D ;
  wire \DFF_74.Q ;
  wire \DFF_740.CK ;
  wire \DFF_740.D ;
  wire \DFF_740.Q ;
  wire \DFF_741.CK ;
  wire \DFF_741.D ;
  wire \DFF_741.Q ;
  wire \DFF_742.CK ;
  wire \DFF_742.D ;
  wire \DFF_742.Q ;
  wire \DFF_743.CK ;
  wire \DFF_743.D ;
  wire \DFF_743.Q ;
  wire \DFF_744.CK ;
  wire \DFF_744.D ;
  wire \DFF_744.Q ;
  wire \DFF_745.CK ;
  wire \DFF_745.D ;
  wire \DFF_745.Q ;
  wire \DFF_746.CK ;
  wire \DFF_746.D ;
  wire \DFF_746.Q ;
  wire \DFF_747.CK ;
  wire \DFF_747.D ;
  wire \DFF_747.Q ;
  wire \DFF_748.CK ;
  wire \DFF_748.D ;
  wire \DFF_748.Q ;
  wire \DFF_749.CK ;
  wire \DFF_749.D ;
  wire \DFF_749.Q ;
  wire \DFF_75.CK ;
  wire \DFF_75.D ;
  wire \DFF_75.Q ;
  wire \DFF_750.CK ;
  wire \DFF_750.D ;
  wire \DFF_750.Q ;
  wire \DFF_751.CK ;
  wire \DFF_751.D ;
  wire \DFF_751.Q ;
  wire \DFF_752.CK ;
  wire \DFF_752.D ;
  wire \DFF_752.Q ;
  wire \DFF_753.CK ;
  wire \DFF_753.D ;
  wire \DFF_753.Q ;
  wire \DFF_754.CK ;
  wire \DFF_754.D ;
  wire \DFF_754.Q ;
  wire \DFF_755.CK ;
  wire \DFF_755.D ;
  wire \DFF_755.Q ;
  wire \DFF_756.CK ;
  wire \DFF_756.D ;
  wire \DFF_756.Q ;
  wire \DFF_757.CK ;
  wire \DFF_757.D ;
  wire \DFF_757.Q ;
  wire \DFF_758.CK ;
  wire \DFF_758.D ;
  wire \DFF_758.Q ;
  wire \DFF_759.CK ;
  wire \DFF_759.D ;
  wire \DFF_759.Q ;
  wire \DFF_76.CK ;
  wire \DFF_76.D ;
  wire \DFF_76.Q ;
  wire \DFF_760.CK ;
  wire \DFF_760.D ;
  wire \DFF_760.Q ;
  wire \DFF_761.CK ;
  wire \DFF_761.D ;
  wire \DFF_761.Q ;
  wire \DFF_762.CK ;
  wire \DFF_762.D ;
  wire \DFF_762.Q ;
  wire \DFF_763.CK ;
  wire \DFF_763.D ;
  wire \DFF_763.Q ;
  wire \DFF_764.CK ;
  wire \DFF_764.D ;
  wire \DFF_764.Q ;
  wire \DFF_765.CK ;
  wire \DFF_765.D ;
  wire \DFF_765.Q ;
  wire \DFF_766.CK ;
  wire \DFF_766.D ;
  wire \DFF_766.Q ;
  wire \DFF_767.CK ;
  wire \DFF_767.D ;
  wire \DFF_767.Q ;
  wire \DFF_768.CK ;
  wire \DFF_768.D ;
  wire \DFF_768.Q ;
  wire \DFF_769.CK ;
  wire \DFF_769.D ;
  wire \DFF_769.Q ;
  wire \DFF_77.CK ;
  wire \DFF_77.D ;
  wire \DFF_77.Q ;
  wire \DFF_770.CK ;
  wire \DFF_770.D ;
  wire \DFF_770.Q ;
  wire \DFF_771.CK ;
  wire \DFF_771.D ;
  wire \DFF_771.Q ;
  wire \DFF_772.CK ;
  wire \DFF_772.D ;
  wire \DFF_772.Q ;
  wire \DFF_773.CK ;
  wire \DFF_773.D ;
  wire \DFF_773.Q ;
  wire \DFF_774.CK ;
  wire \DFF_774.D ;
  wire \DFF_774.Q ;
  wire \DFF_775.CK ;
  wire \DFF_775.D ;
  wire \DFF_775.Q ;
  wire \DFF_776.CK ;
  wire \DFF_776.D ;
  wire \DFF_776.Q ;
  wire \DFF_777.CK ;
  wire \DFF_777.D ;
  wire \DFF_777.Q ;
  wire \DFF_778.CK ;
  wire \DFF_778.D ;
  wire \DFF_778.Q ;
  wire \DFF_779.CK ;
  wire \DFF_779.D ;
  wire \DFF_779.Q ;
  wire \DFF_78.CK ;
  wire \DFF_78.D ;
  wire \DFF_78.Q ;
  wire \DFF_780.CK ;
  wire \DFF_780.D ;
  wire \DFF_780.Q ;
  wire \DFF_781.CK ;
  wire \DFF_781.D ;
  wire \DFF_781.Q ;
  wire \DFF_782.CK ;
  wire \DFF_782.D ;
  wire \DFF_782.Q ;
  wire \DFF_783.CK ;
  wire \DFF_783.D ;
  wire \DFF_783.Q ;
  wire \DFF_784.CK ;
  wire \DFF_784.D ;
  wire \DFF_784.Q ;
  wire \DFF_785.CK ;
  wire \DFF_785.D ;
  wire \DFF_785.Q ;
  wire \DFF_786.CK ;
  wire \DFF_786.D ;
  wire \DFF_786.Q ;
  wire \DFF_787.CK ;
  wire \DFF_787.D ;
  wire \DFF_787.Q ;
  wire \DFF_788.CK ;
  wire \DFF_788.D ;
  wire \DFF_788.Q ;
  wire \DFF_789.CK ;
  wire \DFF_789.D ;
  wire \DFF_789.Q ;
  wire \DFF_79.CK ;
  wire \DFF_79.D ;
  wire \DFF_79.Q ;
  wire \DFF_790.CK ;
  wire \DFF_790.D ;
  wire \DFF_790.Q ;
  wire \DFF_791.CK ;
  wire \DFF_791.D ;
  wire \DFF_791.Q ;
  wire \DFF_792.CK ;
  wire \DFF_792.D ;
  wire \DFF_792.Q ;
  wire \DFF_793.CK ;
  wire \DFF_793.D ;
  wire \DFF_793.Q ;
  wire \DFF_794.CK ;
  wire \DFF_794.D ;
  wire \DFF_794.Q ;
  wire \DFF_795.CK ;
  wire \DFF_795.D ;
  wire \DFF_795.Q ;
  wire \DFF_796.CK ;
  wire \DFF_796.D ;
  wire \DFF_796.Q ;
  wire \DFF_797.CK ;
  wire \DFF_797.D ;
  wire \DFF_797.Q ;
  wire \DFF_798.CK ;
  wire \DFF_798.D ;
  wire \DFF_798.Q ;
  wire \DFF_799.CK ;
  wire \DFF_799.D ;
  wire \DFF_799.Q ;
  wire \DFF_8.CK ;
  wire \DFF_8.D ;
  wire \DFF_8.Q ;
  wire \DFF_80.CK ;
  wire \DFF_80.D ;
  wire \DFF_80.Q ;
  wire \DFF_800.CK ;
  wire \DFF_800.D ;
  wire \DFF_800.Q ;
  wire \DFF_801.CK ;
  wire \DFF_801.D ;
  wire \DFF_801.Q ;
  wire \DFF_802.CK ;
  wire \DFF_802.D ;
  wire \DFF_802.Q ;
  wire \DFF_803.CK ;
  wire \DFF_803.D ;
  wire \DFF_803.Q ;
  wire \DFF_804.CK ;
  wire \DFF_804.D ;
  wire \DFF_804.Q ;
  wire \DFF_805.CK ;
  wire \DFF_805.D ;
  wire \DFF_805.Q ;
  wire \DFF_806.CK ;
  wire \DFF_806.D ;
  wire \DFF_806.Q ;
  wire \DFF_807.CK ;
  wire \DFF_807.D ;
  wire \DFF_807.Q ;
  wire \DFF_808.CK ;
  wire \DFF_808.D ;
  wire \DFF_808.Q ;
  wire \DFF_809.CK ;
  wire \DFF_809.D ;
  wire \DFF_809.Q ;
  wire \DFF_81.CK ;
  wire \DFF_81.D ;
  wire \DFF_81.Q ;
  wire \DFF_810.CK ;
  wire \DFF_810.D ;
  wire \DFF_810.Q ;
  wire \DFF_811.CK ;
  wire \DFF_811.D ;
  wire \DFF_811.Q ;
  wire \DFF_812.CK ;
  wire \DFF_812.D ;
  wire \DFF_812.Q ;
  wire \DFF_813.CK ;
  wire \DFF_813.D ;
  wire \DFF_813.Q ;
  wire \DFF_814.CK ;
  wire \DFF_814.D ;
  wire \DFF_814.Q ;
  wire \DFF_815.CK ;
  wire \DFF_815.D ;
  wire \DFF_815.Q ;
  wire \DFF_816.CK ;
  wire \DFF_816.D ;
  wire \DFF_816.Q ;
  wire \DFF_817.CK ;
  wire \DFF_817.D ;
  wire \DFF_817.Q ;
  wire \DFF_818.CK ;
  wire \DFF_818.D ;
  wire \DFF_818.Q ;
  wire \DFF_819.CK ;
  wire \DFF_819.D ;
  wire \DFF_819.Q ;
  wire \DFF_82.CK ;
  wire \DFF_82.D ;
  wire \DFF_82.Q ;
  wire \DFF_820.CK ;
  wire \DFF_820.D ;
  wire \DFF_820.Q ;
  wire \DFF_821.CK ;
  wire \DFF_821.D ;
  wire \DFF_821.Q ;
  wire \DFF_822.CK ;
  wire \DFF_822.D ;
  wire \DFF_822.Q ;
  wire \DFF_823.CK ;
  wire \DFF_823.D ;
  wire \DFF_823.Q ;
  wire \DFF_824.CK ;
  wire \DFF_824.D ;
  wire \DFF_824.Q ;
  wire \DFF_825.CK ;
  wire \DFF_825.D ;
  wire \DFF_825.Q ;
  wire \DFF_826.CK ;
  wire \DFF_826.D ;
  wire \DFF_826.Q ;
  wire \DFF_827.CK ;
  wire \DFF_827.D ;
  wire \DFF_827.Q ;
  wire \DFF_828.CK ;
  wire \DFF_828.D ;
  wire \DFF_828.Q ;
  wire \DFF_829.CK ;
  wire \DFF_829.D ;
  wire \DFF_829.Q ;
  wire \DFF_83.CK ;
  wire \DFF_83.D ;
  wire \DFF_83.Q ;
  wire \DFF_830.CK ;
  wire \DFF_830.D ;
  wire \DFF_830.Q ;
  wire \DFF_831.CK ;
  wire \DFF_831.D ;
  wire \DFF_831.Q ;
  wire \DFF_832.CK ;
  wire \DFF_832.D ;
  wire \DFF_832.Q ;
  wire \DFF_833.CK ;
  wire \DFF_833.D ;
  wire \DFF_833.Q ;
  wire \DFF_834.CK ;
  wire \DFF_834.D ;
  wire \DFF_834.Q ;
  wire \DFF_835.CK ;
  wire \DFF_835.D ;
  wire \DFF_835.Q ;
  wire \DFF_836.CK ;
  wire \DFF_836.D ;
  wire \DFF_836.Q ;
  wire \DFF_837.CK ;
  wire \DFF_837.D ;
  wire \DFF_837.Q ;
  wire \DFF_838.CK ;
  wire \DFF_838.D ;
  wire \DFF_838.Q ;
  wire \DFF_839.CK ;
  wire \DFF_839.D ;
  wire \DFF_839.Q ;
  wire \DFF_84.CK ;
  wire \DFF_84.D ;
  wire \DFF_84.Q ;
  wire \DFF_840.CK ;
  wire \DFF_840.D ;
  wire \DFF_840.Q ;
  wire \DFF_841.CK ;
  wire \DFF_841.D ;
  wire \DFF_841.Q ;
  wire \DFF_842.CK ;
  wire \DFF_842.D ;
  wire \DFF_842.Q ;
  wire \DFF_843.CK ;
  wire \DFF_843.D ;
  wire \DFF_843.Q ;
  wire \DFF_844.CK ;
  wire \DFF_844.D ;
  wire \DFF_844.Q ;
  wire \DFF_845.CK ;
  wire \DFF_845.D ;
  wire \DFF_845.Q ;
  wire \DFF_846.CK ;
  wire \DFF_846.D ;
  wire \DFF_846.Q ;
  wire \DFF_847.CK ;
  wire \DFF_847.D ;
  wire \DFF_847.Q ;
  wire \DFF_848.CK ;
  wire \DFF_848.D ;
  wire \DFF_848.Q ;
  wire \DFF_849.CK ;
  wire \DFF_849.D ;
  wire \DFF_849.Q ;
  wire \DFF_85.CK ;
  wire \DFF_85.D ;
  wire \DFF_85.Q ;
  wire \DFF_850.CK ;
  wire \DFF_850.D ;
  wire \DFF_850.Q ;
  wire \DFF_851.CK ;
  wire \DFF_851.D ;
  wire \DFF_851.Q ;
  wire \DFF_852.CK ;
  wire \DFF_852.D ;
  wire \DFF_852.Q ;
  wire \DFF_853.CK ;
  wire \DFF_853.D ;
  wire \DFF_853.Q ;
  wire \DFF_854.CK ;
  wire \DFF_854.D ;
  wire \DFF_854.Q ;
  wire \DFF_855.CK ;
  wire \DFF_855.D ;
  wire \DFF_855.Q ;
  wire \DFF_856.CK ;
  wire \DFF_856.D ;
  wire \DFF_856.Q ;
  wire \DFF_857.CK ;
  wire \DFF_857.D ;
  wire \DFF_857.Q ;
  wire \DFF_858.CK ;
  wire \DFF_858.D ;
  wire \DFF_858.Q ;
  wire \DFF_859.CK ;
  wire \DFF_859.D ;
  wire \DFF_859.Q ;
  wire \DFF_86.CK ;
  wire \DFF_86.D ;
  wire \DFF_86.Q ;
  wire \DFF_860.CK ;
  wire \DFF_860.D ;
  wire \DFF_860.Q ;
  wire \DFF_861.CK ;
  wire \DFF_861.D ;
  wire \DFF_861.Q ;
  wire \DFF_862.CK ;
  wire \DFF_862.D ;
  wire \DFF_862.Q ;
  wire \DFF_863.CK ;
  wire \DFF_863.D ;
  wire \DFF_863.Q ;
  wire \DFF_864.CK ;
  wire \DFF_864.D ;
  wire \DFF_864.Q ;
  wire \DFF_865.CK ;
  wire \DFF_865.D ;
  wire \DFF_865.Q ;
  wire \DFF_866.CK ;
  wire \DFF_866.D ;
  wire \DFF_866.Q ;
  wire \DFF_867.CK ;
  wire \DFF_867.D ;
  wire \DFF_867.Q ;
  wire \DFF_868.CK ;
  wire \DFF_868.D ;
  wire \DFF_868.Q ;
  wire \DFF_869.CK ;
  wire \DFF_869.D ;
  wire \DFF_869.Q ;
  wire \DFF_87.CK ;
  wire \DFF_87.D ;
  wire \DFF_87.Q ;
  wire \DFF_870.CK ;
  wire \DFF_870.D ;
  wire \DFF_870.Q ;
  wire \DFF_871.CK ;
  wire \DFF_871.D ;
  wire \DFF_871.Q ;
  wire \DFF_872.CK ;
  wire \DFF_872.D ;
  wire \DFF_872.Q ;
  wire \DFF_873.CK ;
  wire \DFF_873.D ;
  wire \DFF_873.Q ;
  wire \DFF_874.CK ;
  wire \DFF_874.D ;
  wire \DFF_874.Q ;
  wire \DFF_875.CK ;
  wire \DFF_875.D ;
  wire \DFF_875.Q ;
  wire \DFF_876.CK ;
  wire \DFF_876.D ;
  wire \DFF_876.Q ;
  wire \DFF_877.CK ;
  wire \DFF_877.D ;
  wire \DFF_877.Q ;
  wire \DFF_878.CK ;
  wire \DFF_878.D ;
  wire \DFF_878.Q ;
  wire \DFF_879.CK ;
  wire \DFF_879.D ;
  wire \DFF_879.Q ;
  wire \DFF_88.CK ;
  wire \DFF_88.D ;
  wire \DFF_88.Q ;
  wire \DFF_880.CK ;
  wire \DFF_880.D ;
  wire \DFF_880.Q ;
  wire \DFF_881.CK ;
  wire \DFF_881.D ;
  wire \DFF_881.Q ;
  wire \DFF_882.CK ;
  wire \DFF_882.D ;
  wire \DFF_882.Q ;
  wire \DFF_883.CK ;
  wire \DFF_883.D ;
  wire \DFF_883.Q ;
  wire \DFF_884.CK ;
  wire \DFF_884.D ;
  wire \DFF_884.Q ;
  wire \DFF_885.CK ;
  wire \DFF_885.D ;
  wire \DFF_885.Q ;
  wire \DFF_886.CK ;
  wire \DFF_886.D ;
  wire \DFF_886.Q ;
  wire \DFF_887.CK ;
  wire \DFF_887.D ;
  wire \DFF_887.Q ;
  wire \DFF_888.CK ;
  wire \DFF_888.D ;
  wire \DFF_888.Q ;
  wire \DFF_889.CK ;
  wire \DFF_889.D ;
  wire \DFF_889.Q ;
  wire \DFF_89.CK ;
  wire \DFF_89.D ;
  wire \DFF_89.Q ;
  wire \DFF_890.CK ;
  wire \DFF_890.D ;
  wire \DFF_890.Q ;
  wire \DFF_891.CK ;
  wire \DFF_891.D ;
  wire \DFF_891.Q ;
  wire \DFF_892.CK ;
  wire \DFF_892.D ;
  wire \DFF_892.Q ;
  wire \DFF_893.CK ;
  wire \DFF_893.D ;
  wire \DFF_893.Q ;
  wire \DFF_894.CK ;
  wire \DFF_894.D ;
  wire \DFF_894.Q ;
  wire \DFF_895.CK ;
  wire \DFF_895.D ;
  wire \DFF_895.Q ;
  wire \DFF_896.CK ;
  wire \DFF_896.D ;
  wire \DFF_896.Q ;
  wire \DFF_897.CK ;
  wire \DFF_897.D ;
  wire \DFF_897.Q ;
  wire \DFF_898.CK ;
  wire \DFF_898.D ;
  wire \DFF_898.Q ;
  wire \DFF_899.CK ;
  wire \DFF_899.D ;
  wire \DFF_899.Q ;
  wire \DFF_9.CK ;
  wire \DFF_9.D ;
  wire \DFF_9.Q ;
  wire \DFF_90.CK ;
  wire \DFF_90.D ;
  wire \DFF_90.Q ;
  wire \DFF_900.CK ;
  wire \DFF_900.D ;
  wire \DFF_900.Q ;
  wire \DFF_901.CK ;
  wire \DFF_901.D ;
  wire \DFF_901.Q ;
  wire \DFF_902.CK ;
  wire \DFF_902.D ;
  wire \DFF_902.Q ;
  wire \DFF_903.CK ;
  wire \DFF_903.D ;
  wire \DFF_903.Q ;
  wire \DFF_904.CK ;
  wire \DFF_904.D ;
  wire \DFF_904.Q ;
  wire \DFF_905.CK ;
  wire \DFF_905.D ;
  wire \DFF_905.Q ;
  wire \DFF_906.CK ;
  wire \DFF_906.D ;
  wire \DFF_906.Q ;
  wire \DFF_907.CK ;
  wire \DFF_907.D ;
  wire \DFF_907.Q ;
  wire \DFF_908.CK ;
  wire \DFF_908.D ;
  wire \DFF_908.Q ;
  wire \DFF_909.CK ;
  wire \DFF_909.D ;
  wire \DFF_909.Q ;
  wire \DFF_91.CK ;
  wire \DFF_91.D ;
  wire \DFF_91.Q ;
  wire \DFF_910.CK ;
  wire \DFF_910.D ;
  wire \DFF_910.Q ;
  wire \DFF_911.CK ;
  wire \DFF_911.D ;
  wire \DFF_911.Q ;
  wire \DFF_912.CK ;
  wire \DFF_912.D ;
  wire \DFF_912.Q ;
  wire \DFF_913.CK ;
  wire \DFF_913.D ;
  wire \DFF_913.Q ;
  wire \DFF_914.CK ;
  wire \DFF_914.D ;
  wire \DFF_914.Q ;
  wire \DFF_915.CK ;
  wire \DFF_915.D ;
  wire \DFF_915.Q ;
  wire \DFF_916.CK ;
  wire \DFF_916.D ;
  wire \DFF_916.Q ;
  wire \DFF_917.CK ;
  wire \DFF_917.D ;
  wire \DFF_917.Q ;
  wire \DFF_918.CK ;
  wire \DFF_918.D ;
  wire \DFF_918.Q ;
  wire \DFF_919.CK ;
  wire \DFF_919.D ;
  wire \DFF_919.Q ;
  wire \DFF_92.CK ;
  wire \DFF_92.D ;
  wire \DFF_92.Q ;
  wire \DFF_920.CK ;
  wire \DFF_920.D ;
  wire \DFF_920.Q ;
  wire \DFF_921.CK ;
  wire \DFF_921.D ;
  wire \DFF_921.Q ;
  wire \DFF_922.CK ;
  wire \DFF_922.D ;
  wire \DFF_922.Q ;
  wire \DFF_923.CK ;
  wire \DFF_923.D ;
  wire \DFF_923.Q ;
  wire \DFF_924.CK ;
  wire \DFF_924.D ;
  wire \DFF_924.Q ;
  wire \DFF_925.CK ;
  wire \DFF_925.D ;
  wire \DFF_925.Q ;
  wire \DFF_926.CK ;
  wire \DFF_926.D ;
  wire \DFF_926.Q ;
  wire \DFF_927.CK ;
  wire \DFF_927.D ;
  wire \DFF_927.Q ;
  wire \DFF_928.CK ;
  wire \DFF_928.D ;
  wire \DFF_928.Q ;
  wire \DFF_929.CK ;
  wire \DFF_929.D ;
  wire \DFF_929.Q ;
  wire \DFF_93.CK ;
  wire \DFF_93.D ;
  wire \DFF_93.Q ;
  wire \DFF_930.CK ;
  wire \DFF_930.D ;
  wire \DFF_930.Q ;
  wire \DFF_931.CK ;
  wire \DFF_931.D ;
  wire \DFF_931.Q ;
  wire \DFF_932.CK ;
  wire \DFF_932.D ;
  wire \DFF_932.Q ;
  wire \DFF_933.CK ;
  wire \DFF_933.D ;
  wire \DFF_933.Q ;
  wire \DFF_934.CK ;
  wire \DFF_934.D ;
  wire \DFF_934.Q ;
  wire \DFF_935.CK ;
  wire \DFF_935.D ;
  wire \DFF_935.Q ;
  wire \DFF_936.CK ;
  wire \DFF_936.D ;
  wire \DFF_936.Q ;
  wire \DFF_937.CK ;
  wire \DFF_937.D ;
  wire \DFF_937.Q ;
  wire \DFF_938.CK ;
  wire \DFF_938.D ;
  wire \DFF_938.Q ;
  wire \DFF_939.CK ;
  wire \DFF_939.D ;
  wire \DFF_939.Q ;
  wire \DFF_94.CK ;
  wire \DFF_94.D ;
  wire \DFF_94.Q ;
  wire \DFF_940.CK ;
  wire \DFF_940.D ;
  wire \DFF_940.Q ;
  wire \DFF_941.CK ;
  wire \DFF_941.D ;
  wire \DFF_941.Q ;
  wire \DFF_942.CK ;
  wire \DFF_942.D ;
  wire \DFF_942.Q ;
  wire \DFF_943.CK ;
  wire \DFF_943.D ;
  wire \DFF_943.Q ;
  wire \DFF_944.CK ;
  wire \DFF_944.D ;
  wire \DFF_944.Q ;
  wire \DFF_945.CK ;
  wire \DFF_945.D ;
  wire \DFF_945.Q ;
  wire \DFF_946.CK ;
  wire \DFF_946.D ;
  wire \DFF_946.Q ;
  wire \DFF_947.CK ;
  wire \DFF_947.D ;
  wire \DFF_947.Q ;
  wire \DFF_948.CK ;
  wire \DFF_948.D ;
  wire \DFF_948.Q ;
  wire \DFF_949.CK ;
  wire \DFF_949.D ;
  wire \DFF_949.Q ;
  wire \DFF_95.CK ;
  wire \DFF_95.D ;
  wire \DFF_95.Q ;
  wire \DFF_950.CK ;
  wire \DFF_950.D ;
  wire \DFF_950.Q ;
  wire \DFF_951.CK ;
  wire \DFF_951.D ;
  wire \DFF_951.Q ;
  wire \DFF_952.CK ;
  wire \DFF_952.D ;
  wire \DFF_952.Q ;
  wire \DFF_953.CK ;
  wire \DFF_953.D ;
  wire \DFF_953.Q ;
  wire \DFF_954.CK ;
  wire \DFF_954.D ;
  wire \DFF_954.Q ;
  wire \DFF_955.CK ;
  wire \DFF_955.D ;
  wire \DFF_955.Q ;
  wire \DFF_956.CK ;
  wire \DFF_956.D ;
  wire \DFF_956.Q ;
  wire \DFF_957.CK ;
  wire \DFF_957.D ;
  wire \DFF_957.Q ;
  wire \DFF_958.CK ;
  wire \DFF_958.D ;
  wire \DFF_958.Q ;
  wire \DFF_959.CK ;
  wire \DFF_959.D ;
  wire \DFF_959.Q ;
  wire \DFF_96.CK ;
  wire \DFF_96.D ;
  wire \DFF_96.Q ;
  wire \DFF_960.CK ;
  wire \DFF_960.D ;
  wire \DFF_960.Q ;
  wire \DFF_961.CK ;
  wire \DFF_961.D ;
  wire \DFF_961.Q ;
  wire \DFF_962.CK ;
  wire \DFF_962.D ;
  wire \DFF_962.Q ;
  wire \DFF_963.CK ;
  wire \DFF_963.D ;
  wire \DFF_963.Q ;
  wire \DFF_964.CK ;
  wire \DFF_964.D ;
  wire \DFF_964.Q ;
  wire \DFF_965.CK ;
  wire \DFF_965.D ;
  wire \DFF_965.Q ;
  wire \DFF_966.CK ;
  wire \DFF_966.D ;
  wire \DFF_966.Q ;
  wire \DFF_967.CK ;
  wire \DFF_967.D ;
  wire \DFF_967.Q ;
  wire \DFF_968.CK ;
  wire \DFF_968.D ;
  wire \DFF_968.Q ;
  wire \DFF_969.CK ;
  wire \DFF_969.D ;
  wire \DFF_969.Q ;
  wire \DFF_97.CK ;
  wire \DFF_97.D ;
  wire \DFF_97.Q ;
  wire \DFF_970.CK ;
  wire \DFF_970.D ;
  wire \DFF_970.Q ;
  wire \DFF_971.CK ;
  wire \DFF_971.D ;
  wire \DFF_971.Q ;
  wire \DFF_972.CK ;
  wire \DFF_972.D ;
  wire \DFF_972.Q ;
  wire \DFF_973.CK ;
  wire \DFF_973.D ;
  wire \DFF_973.Q ;
  wire \DFF_974.CK ;
  wire \DFF_974.D ;
  wire \DFF_974.Q ;
  wire \DFF_975.CK ;
  wire \DFF_975.D ;
  wire \DFF_975.Q ;
  wire \DFF_976.CK ;
  wire \DFF_976.D ;
  wire \DFF_976.Q ;
  wire \DFF_977.CK ;
  wire \DFF_977.D ;
  wire \DFF_977.Q ;
  wire \DFF_978.CK ;
  wire \DFF_978.D ;
  wire \DFF_978.Q ;
  wire \DFF_979.CK ;
  wire \DFF_979.D ;
  wire \DFF_979.Q ;
  wire \DFF_98.CK ;
  wire \DFF_98.D ;
  wire \DFF_98.Q ;
  wire \DFF_980.CK ;
  wire \DFF_980.D ;
  wire \DFF_980.Q ;
  wire \DFF_981.CK ;
  wire \DFF_981.D ;
  wire \DFF_981.Q ;
  wire \DFF_982.CK ;
  wire \DFF_982.D ;
  wire \DFF_982.Q ;
  wire \DFF_983.CK ;
  wire \DFF_983.D ;
  wire \DFF_983.Q ;
  wire \DFF_984.CK ;
  wire \DFF_984.D ;
  wire \DFF_984.Q ;
  wire \DFF_985.CK ;
  wire \DFF_985.D ;
  wire \DFF_985.Q ;
  wire \DFF_986.CK ;
  wire \DFF_986.D ;
  wire \DFF_986.Q ;
  wire \DFF_987.CK ;
  wire \DFF_987.D ;
  wire \DFF_987.Q ;
  wire \DFF_988.CK ;
  wire \DFF_988.D ;
  wire \DFF_988.Q ;
  wire \DFF_989.CK ;
  wire \DFF_989.D ;
  wire \DFF_989.Q ;
  wire \DFF_99.CK ;
  wire \DFF_99.D ;
  wire \DFF_99.Q ;
  wire \DFF_990.CK ;
  wire \DFF_990.D ;
  wire \DFF_990.Q ;
  wire \DFF_991.CK ;
  wire \DFF_991.D ;
  wire \DFF_991.Q ;
  wire \DFF_992.CK ;
  wire \DFF_992.D ;
  wire \DFF_992.Q ;
  wire \DFF_993.CK ;
  wire \DFF_993.D ;
  wire \DFF_993.Q ;
  wire \DFF_994.CK ;
  wire \DFF_994.D ;
  wire \DFF_994.Q ;
  wire \DFF_995.CK ;
  wire \DFF_995.D ;
  wire \DFF_995.Q ;
  wire \DFF_996.CK ;
  wire \DFF_996.D ;
  wire \DFF_996.Q ;
  wire \DFF_997.CK ;
  wire \DFF_997.D ;
  wire \DFF_997.Q ;
  wire \DFF_998.CK ;
  wire \DFF_998.D ;
  wire \DFF_998.Q ;
  wire \DFF_999.CK ;
  wire \DFF_999.D ;
  wire \DFF_999.Q ;
  input GND;
  wire I13708;
  wire I13847;
  wire I13968;
  wire I13979;
  wire I13990;
  wire I13995;
  wire I14033;
  wire I14046;
  wire I14050;
  wire I14054;
  wire I14079;
  wire I14119;
  wire I14222;
  wire I14241;
  wire I14267;
  wire I14271;
  wire I14301;
  wire I14326;
  wire I14381;
  wire I14409;
  wire I14455;
  wire I14475;
  wire I14505;
  wire I14537;
  wire I14550;
  wire I14567;
  wire I14584;
  wire I14593;
  wire I14679;
  wire I14742;
  wire I14773;
  wire I14797;
  wire I14823;
  wire I14827;
  wire I14836;
  wire I14839;
  wire I14862;
  wire I14866;
  wire I14893;
  wire I14896;
  wire I14902;
  wire I14905;
  wire I14932;
  wire I14935;
  wire I14967;
  wire I14970;
  wire I14999;
  wire I15030;
  wire I15033;
  wire I15070;
  wire I15073;
  wire I15162;
  wire I15205;
  wire I15223;
  wire I15250;
  wire I15382;
  wire I15448;
  wire I15474;
  wire I15533;
  wire I15550;
  wire I15556;
  wire I15564;
  wire I15569;
  wire I15577;
  wire I15587;
  wire I15590;
  wire I15593;
  wire I15600;
  wire I15609;
  wire I15617;
  wire I15620;
  wire I15623;
  wire I15626;
  wire I15633;
  wire I15636;
  wire I15647;
  wire I15650;
  wire I15667;
  wire I15682;
  wire I15702;
  wire I15705;
  wire I15727;
  wire I15736;
  wire I15773;
  wire I15782;
  wire I15788;
  wire I15811;
  wire I15814;
  wire I15821;
  wire I15831;
  wire I15834;
  wire I15843;
  wire I15846;
  wire I15862;
  wire I15869;
  wire I15878;
  wire I15893;
  wire I15906;
  wire I15915;
  wire I15918;
  wire I15921;
  wire I15929;
  wire I15932;
  wire I15942;
  wire I15954;
  wire I15981;
  wire I15987;
  wire I16028;
  wire I16040;
  wire I16057;
  wire I16077;
  wire I16090;
  wire I16102;
  wire I16117;
  wire I16120;
  wire I16135;
  wire I16150;
  wire I16163;
  wire I16289;
  wire I16438;
  wire I16452;
  wire I16460;
  wire I16468;
  wire I16471;
  wire I16476;
  wire I16479;
  wire I16486;
  wire I16489;
  wire I16492;
  wire I16498;
  wire I16502;
  wire I16512;
  wire I16521;
  wire I16526;
  wire I16535;
  wire I16538;
  wire I16555;
  wire I16564;
  wire I16579;
  wire I16593;
  wire I16596;
  wire I16610;
  wire I16613;
  wire I16651;
  wire I16660;
  wire I16663;
  wire I16688;
  wire I16709;
  wire I16775;
  wire I17008;
  wire I17094;
  wire I17098;
  wire I17101;
  wire I17104;
  wire I17108;
  wire I17111;
  wire I17114;
  wire I17118;
  wire I17121;
  wire I17125;
  wire I17128;
  wire I17131;
  wire I17136;
  wire I17140;
  wire I17143;
  wire I17148;
  wire I17154;
  wire I17159;
  wire I17166;
  wire I17173;
  wire I17181;
  wire I17188;
  wire I17198;
  wire I17207;
  wire I17228;
  wire I17249;
  wire I17276;
  wire I17355;
  wire I17374;
  wire I17392;
  wire I17401;
  wire I17420;
  wire I17425;
  wire I17436;
  wire I17442;
  wire I17456;
  wire I17471;
  wire I17488;
  wire I17491;
  wire I17507;
  wire I17590;
  wire I17609;
  wire I17612;
  wire I17615;
  wire I17633;
  wire I17636;
  wire I17639;
  wire I17650;
  wire I17653;
  wire I17658;
  wire I17661;
  wire I17668;
  wire I17671;
  wire I17675;
  wire I17679;
  wire I17695;
  wire I17699;
  wire I17704;
  wire I17723;
  wire I17747;
  wire I17750;
  wire I17763;
  wire I17780;
  wire I17808;
  wire I17976;
  wire I18003;
  wire I18006;
  wire I18009;
  wire I18028;
  wire I18031;
  wire I18034;
  wire I18048;
  wire I18051;
  wire I18071;
  wire I18078;
  wire I18083;
  wire I18089;
  wire I18101;
  wire I18104;
  wire I18120;
  wire I18125;
  wire I18131;
  wire I18135;
  wire I18143;
  wire I18151;
  wire I18154;
  wire I18165;
  wire I18168;
  wire I18177;
  wire I18180;
  wire I18214;
  wire I18221;
  wire I18224;
  wire I18238;
  wire I18245;
  wire I18248;
  wire I18252;
  wire I18259;
  wire I18262;
  wire I18265;
  wire I18270;
  wire I18280;
  wire I18285;
  wire I18301;
  wire I18307;
  wire I18310;
  wire I18313;
  wire I18320;
  wire I18323;
  wire I18341;
  wire I18344;
  wire I18350;
  wire I18364;
  wire I18367;
  wire I18373;
  wire I18376;
  wire I18379;
  wire I18382;
  wire I18398;
  wire I18408;
  wire I18411;
  wire I18434;
  wire I18443;
  wire I18446;
  wire I18469;
  wire I18476;
  wire I18479;
  wire I18482;
  wire I18518;
  wire I18523;
  wire I18526;
  wire I18571;
  wire I18574;
  wire I18674;
  wire I18810;
  wire I18822;
  wire I18829;
  wire I18832;
  wire I18839;
  wire I18842;
  wire I18849;
  wire I18852;
  wire I18855;
  wire I18858;
  wire I18861;
  wire I18865;
  wire I18868;
  wire I18872;
  wire I18875;
  wire I18879;
  wire I19384;
  wire I19661;
  wire I19707;
  wire I19719;
  wire I19756;
  wire I19772;
  wire I19786;
  wire I19796;
  wire I19813;
  wire I19927;
  wire I20216;
  wire I20529;
  wire I20542;
  wire I20562;
  wire I20584;
  wire I20690;
  wire I20846;
  wire I20895;
  wire I20913;
  wire I20937;
  wire I21006;
  wire I21033;
  wire I21036;
  wire I21067;
  wire I21100;
  wire I21115;
  wire I21181;
  wire I21189;
  wire I21199;
  wire I21210;
  wire I21222;
  wire I21810;
  wire I21922;
  wire I21934;
  wire I22031;
  wire I22177;
  wire I22180;
  wire I22745;
  wire I22748;
  wire I22785;
  wire I22788;
  wire I22886;
  wire I22889;
  wire I24920;
  wire I26195;
  wire I26479;
  wire I26503;
  wire I26508;
  wire I26516;
  wire I26705;
  wire I26880;
  wire I26925;
  wire I27232;
  wire I27253;
  wire I27314;
  wire I27579;
  wire I27730;
  wire I27735;
  wire I27749;
  wire I28349;
  wire I28576;
  wire I28582;
  wire I28588;
  wire I28591;
  wire I28594;
  wire I29371;
  input VDD;
  wire g1;
  input g100;
  wire g10003;
  wire g1002;
  wire g10029;
  wire g10031;
  wire g10061;
  wire g1008;
  wire g10087;
  wire g101;
  wire g10107;
  output g10122;
  wire g10139;
  wire g10141;
  wire g10142;
  wire g1018;
  wire g10198;
  wire g102;
  wire g10216;
  wire g10230;
  wire g10233;
  wire g1024;
  wire g10272;
  wire g10273;
  wire g10287;
  wire g10288;
  wire g10295;
  wire g1030;
  output g10306;
  wire g10318;
  wire g10319;
  wire g10323;
  wire g10347;
  wire g10348;
  wire g10349;
  wire g10350;
  wire g10351;
  wire g10352;
  wire g10353;
  wire g10354;
  wire g10355;
  wire g10356;
  wire g10357;
  wire g10358;
  wire g10359;
  wire g1036;
  wire g10360;
  wire g10361;
  wire g10362;
  wire g10363;
  wire g10366;
  wire g10367;
  wire g10368;
  wire g10369;
  wire g10370;
  wire g10371;
  wire g10372;
  wire g10373;
  wire g10374;
  wire g10375;
  wire g10376;
  wire g10377;
  wire g10378;
  wire g10379;
  wire g10380;
  wire g10381;
  wire g10382;
  wire g10383;
  wire g10384;
  wire g10385;
  wire g10386;
  wire g10387;
  wire g10388;
  wire g10389;
  wire g10390;
  wire g10391;
  wire g10392;
  wire g10393;
  wire g10394;
  wire g10395;
  wire g10396;
  wire g10397;
  wire g10398;
  wire g10399;
  wire g10400;
  wire g10401;
  wire g10402;
  wire g10403;
  wire g10404;
  wire g10405;
  wire g10406;
  wire g10407;
  wire g10408;
  wire g10409;
  wire g1041;
  wire g10410;
  wire g10411;
  wire g10412;
  wire g10413;
  wire g10414;
  wire g10415;
  wire g10420;
  wire g10427;
  wire g10428;
  wire g1046;
  wire g10473;
  wire g10489;
  wire g10490;
  wire g10497;
  wire g10499;
  output g10500;
  wire g10518;
  wire g10519;
  wire g1052;
  output g10527;
  wire g10540;
  wire g10541;
  wire g1056;
  wire g10564;
  wire g10581;
  wire g10582;
  wire g10588;
  wire g106;
  wire g1061;
  wire g10615;
  wire g10664;
  wire g1070;
  wire g1075;
  wire g1079;
  wire g10795;
  wire g10823;
  wire g1083;
  wire g1087;
  wire g10877;
  wire g1094;
  wire g10960;
  wire g10980;
  wire g1099;
  wire g110;
  wire g11011;
  wire g11017;
  wire g1105;
  wire g111;
  wire g1111;
  wire g11136;
  wire g1116;
  wire g112;
  wire g11237;
  wire g1124;
  wire g1129;
  wire g11290;
  input g113;
  wire g11317;
  output g11349;
  wire g1135;
  output g11388;
  input g114;
  wire g1141;
  output g11418;
  output g11447;
  wire g1146;
  input g115;
  wire g1152;
  wire g1157;
  input g116;
  output g11678;
  wire g117;
  wire g11705;
  wire g11706;
  wire g1171;
  wire g11714;
  wire g11720;
  wire g11721;
  wire g11735;
  wire g11736;
  wire g11741;
  wire g11744;
  wire g11753;
  wire g11754;
  wire g11762;
  wire g11769;
  output g11770;
  wire g11772;
  wire g1178;
  wire g11790;
  wire g11793;
  wire g11796;
  wire g11820;
  wire g11823;
  wire g11826;
  wire g11829;
  wire g1183;
  wire g11832;
  wire g11833;
  wire g11842;
  wire g11845;
  wire g11852;
  wire g11855;
  wire g11861;
  wire g11872;
  wire g11875;
  wire g11878;
  wire g11884;
  wire g1189;
  wire g11894;
  wire g11897;
  wire g11900;
  wire g11917;
  wire g11920;
  wire g11929;
  wire g1193;
  wire g11931;
  wire g11941;
  wire g11966;
  wire g11986;
  wire g11987;
  wire g1199;
  input g120;
  wire g12039;
  wire g1205;
  wire g12077;
  wire g121;
  wire g12108;
  wire g1211;
  wire g1216;
  wire g12183;
  output g12184;
  wire g1221;
  output g12238;
  wire g1227;
  output g12300;
  wire g1233;
  output g12350;
  wire g1236;
  wire g12367;
  output g12368;
  wire g1239;
  wire g12399;
  input g124;
  wire g1242;
  output g12422;
  wire g12430;
  wire g12440;
  wire g1246;
  output g12470;
  wire g12477;
  wire g1249;
  wire g12490;
  input g125;
  wire g1252;
  wire g1256;
  wire g1259;
  input g126;
  wire g1263;
  wire g12640;
  wire g1266;
  input g127;
  wire g1270;
  wire g12729;
  wire g12738;
  wire g1274;
  wire g1277;
  wire g12778;
  wire g12779;
  wire g128;
  wire g1280;
  wire g12804;
  wire g12805;
  wire g12823;
  wire g1283;
  wire g12830;
  wire g12831;
  output g12832;
  output g12833;
  wire g1287;
  wire g12875;
  wire g1291;
  output g12919;
  output g12923;
  wire g12952;
  wire g1296;
  wire g1300;
  wire g13036;
  wire g13037;
  output g13039;
  output g13049;
  wire g13051;
  wire g1306;
  wire g13061;
  wire g13062;
  output g13068;
  wire g13070;
  wire g13082;
  output g13085;
  wire g13087;
  output g13099;
  wire g13106;
  wire g1311;
  wire g13117;
  wire g1312;
  wire g13138;
  wire g13174;
  wire g13189;
  wire g1319;
  wire g1322;
  output g13259;
  output g13272;
  wire g13302;
  wire g1333;
  wire g1339;
  input g134;
  wire g13412;
  wire g1345;
  wire g13484;
  wire g13494;
  input g135;
  wire g13505;
  wire g1351;
  wire g13510;
  wire g13522;
  wire g136;
  wire g1361;
  wire g1367;
  wire g1373;
  wire g1379;
  wire g1384;
  wire g13856;
  output g13865;
  output g13881;
  wire g1389;
  output g13895;
  output g13906;
  output g13926;
  wire g1395;
  output g13966;
  wire g1399;
  wire g1404;
  output g14096;
  output g14125;
  wire g1413;
  output g14147;
  wire g14149;
  wire g14150;
  output g14167;
  wire g14169;
  wire g14173;
  wire g1418;
  wire g14183;
  wire g14184;
  output g14189;
  wire g14191;
  wire g14198;
  wire g142;
  output g14201;
  wire g14203;
  wire g14205;
  output g14217;
  wire g14219;
  wire g1422;
  wire g14255;
  wire g1426;
  wire g14277;
  wire g1430;
  wire g14308;
  wire g14332;
  wire g14357;
  wire g14359;
  wire g1437;
  wire g14385;
  wire g14386;
  wire g1442;
  output g14421;
  wire g14441;
  wire g14443;
  output g14451;
  wire g1448;
  wire g14509;
  wire g14510;
  output g14518;
  wire g1454;
  wire g14562;
  wire g14563;
  wire g14564;
  wire g14582;
  wire g1459;
  output g14597;
  wire g146;
  wire g14609;
  output g14635;
  wire g14639;
  output g14662;
  wire g1467;
  output g14673;
  wire g14676;
  output g14694;
  output g14705;
  wire g1472;
  output g14738;
  output g14749;
  output g14779;
  wire g1478;
  wire g14790;
  output g14828;
  wire g1484;
  wire g14873;
  wire g1489;
  wire g14912;
  wire g1495;
  wire g150;
  wire g1500;
  wire g15078;
  wire g15079;
  wire g15083;
  wire g15084;
  wire g1514;
  wire g1521;
  wire g1526;
  wire g153;
  wire g1532;
  wire g1536;
  wire g1542;
  wire g1548;
  wire g1554;
  wire g1559;
  wire g1564;
  wire g157;
  wire g1570;
  wire g1576;
  wire g1579;
  wire g1582;
  wire g1585;
  wire g1589;
  wire g1592;
  wire g15932;
  wire g16;
  wire g160;
  wire g1600;
  wire g1604;
  wire g1608;
  wire g1612;
  wire g1616;
  wire g1620;
  wire g16216;
  wire g16228;
  wire g1624;
  wire g16284;
  wire g16300;
  wire g1632;
  wire g16320;
  wire g1636;
  wire g164;
  wire g1644;
  wire g1648;
  wire g16530;
  wire g16540;
  wire g1657;
  wire g16579;
  wire g16580;
  output g16603;
  wire g16609;
  output g16624;
  output g16627;
  wire g16631;
  wire g16632;
  wire g1664;
  wire g16643;
  wire g16644;
  output g16656;
  output g16659;
  wire g16661;
  wire g16676;
  wire g16677;
  wire g1668;
  output g16686;
  output g16693;
  wire g16695;
  wire g16708;
  wire g16709;
  output g16718;
  output g16722;
  wire g16726;
  wire g16727;
  wire g16738;
  output g16744;
  output g16748;
  wire g16750;
  wire g16767;
  wire g1677;
  output g16775;
  wire g168;
  wire g1682;
  wire g1687;
  wire g16872;
  wire g16873;
  output g16874;
  wire g1691;
  wire g16920;
  output g16924;
  output g16955;
  wire g16958;
  wire g1696;
  wire g16960;
  wire g16963;
  wire g16968;
  wire g1700;
  wire g17010;
  wire g1706;
  wire g17085;
  wire g17088;
  wire g1710;
  wire g1714;
  wire g17141;
  wire g17155;
  wire g17157;
  wire g17197;
  wire g1720;
  wire g17216;
  wire g17221;
  wire g1724;
  wire g17242;
  wire g1728;
  output g17291;
  wire g17292;
  wire g17301;
  output g17316;
  output g17320;
  wire g17325;
  wire g1736;
  wire g17366;
  wire g174;
  wire g1740;
  output g17400;
  output g17404;
  wire g17408;
  wire g17410;
  wire g17411;
  output g17423;
  wire g17429;
  wire g17431;
  wire g1744;
  wire g17465;
  wire g17466;
  wire g17470;
  wire g17471;
  wire g1748;
  wire g17487;
  wire g17489;
  wire g17491;
  wire g17512;
  output g17519;
  wire g1752;
  wire g1756;
  output g17577;
  output g17580;
  wire g17590;
  wire g1760;
  output g17604;
  output g17607;
  output g17639;
  output g17646;
  output g17649;
  output g17674;
  output g17678;
  wire g1768;
  output g17685;
  output g17688;
  output g17711;
  output g17715;
  wire g1772;
  output g17722;
  wire g17733;
  output g17739;
  output g17743;
  output g17760;
  output g17764;
  output g17778;
  wire g17782;
  output g17787;
  wire g1779;
  wire g17794;
  output g17813;
  output g17819;
  wire g1783;
  output g17845;
  output g17871;
  wire g1792;
  wire g1798;
  wire g1802;
  wire g18088;
  output g18092;
  wire g18093;
  output g18094;
  output g18095;
  output g18096;
  output g18097;
  output g18098;
  output g18099;
  output g18100;
  output g18101;
  wire g1811;
  wire g1816;
  wire g182;
  wire g1821;
  wire g18215;
  wire g18216;
  wire g1825;
  wire g18273;
  wire g18274;
  wire g1830;
  wire g1834;
  wire g1840;
  wire g18421;
  wire g18422;
  wire g1844;
  wire g1848;
  wire g18527;
  wire g18528;
  wire g1854;
  wire g1858;
  wire g18597;
  wire g18598;
  wire g1862;
  wire g18695;
  wire g18696;
  wire g1870;
  wire g18726;
  wire g18727;
  wire g1874;
  wire g1878;
  wire g1882;
  wire g18827;
  wire g18828;
  wire g18829;
  wire g18830;
  wire g18831;
  wire g18832;
  wire g1886;
  wire g18874;
  wire g18875;
  wire g18876;
  wire g18877;
  wire g18878;
  wire g18880;
  output g18881;
  wire g18882;
  wire g18883;
  wire g18884;
  wire g18885;
  wire g18886;
  wire g18887;
  wire g18888;
  wire g18889;
  wire g18891;
  wire g18892;
  wire g18894;
  wire g18895;
  wire g18896;
  wire g18897;
  wire g18898;
  wire g1890;
  wire g18903;
  wire g18904;
  wire g18905;
  wire g18907;
  wire g18908;
  wire g18911;
  wire g18916;
  wire g18917;
  wire g18926;
  wire g18929;
  wire g18931;
  wire g18932;
  wire g18938;
  wire g18939;
  wire g1894;
  wire g18940;
  wire g18944;
  wire g18945;
  wire g18946;
  wire g18947;
  wire g18952;
  wire g18953;
  wire g18954;
  wire g18975;
  wire g18976;
  wire g18977;
  wire g18978;
  wire g18979;
  wire g18980;
  wire g18983;
  wire g18984;
  wire g18988;
  wire g18989;
  wire g18990;
  wire g18991;
  wire g19;
  wire g1902;
  wire g1906;
  wire g19067;
  wire g19068;
  wire g191;
  wire g1913;
  wire g19144;
  wire g1917;
  wire g19208;
  wire g1926;
  wire g19273;
  wire g19276;
  wire g1932;
  wire g19330;
  output g19334;
  wire g19343;
  wire g19345;
  wire g19351;
  wire g19352;
  output g19357;
  wire g1936;
  wire g19360;
  wire g19365;
  wire g19366;
  wire g19368;
  wire g19370;
  wire g19373;
  wire g19376;
  wire g19379;
  wire g19385;
  wire g19386;
  wire g19387;
  wire g19389;
  wire g19394;
  wire g19395;
  wire g19396;
  wire g19397;
  wire g19398;
  wire g19399;
  wire g194;
  wire g19409;
  wire g19410;
  wire g19411;
  wire g19412;
  wire g19414;
  wire g19415;
  wire g19416;
  wire g19417;
  wire g19421;
  wire g19429;
  wire g19431;
  wire g19432;
  wire g19433;
  wire g19434;
  wire g19435;
  wire g19437;
  wire g19438;
  wire g19439;
  wire g19440;
  wire g19443;
  wire g19445;
  wire g19446;
  wire g1945;
  wire g19451;
  wire g19452;
  wire g19454;
  wire g19458;
  wire g19468;
  wire g19469;
  wire g19470;
  wire g19471;
  wire g19472;
  wire g19473;
  wire g19476;
  wire g19477;
  wire g19478;
  wire g19479;
  wire g19480;
  wire g19481;
  wire g19482;
  wire g19489;
  wire g19490;
  wire g19491;
  wire g19492;
  wire g19493;
  wire g19494;
  wire g19498;
  wire g19499;
  wire g1950;
  wire g19503;
  wire g19504;
  wire g19505;
  wire g19517;
  wire g19519;
  wire g19520;
  wire g19523;
  wire g19526;
  wire g19527;
  wire g19528;
  wire g19529;
  wire g19531;
  wire g19532;
  wire g19537;
  wire g19538;
  wire g19539;
  wire g19541;
  wire g19542;
  wire g19543;
  wire g19544;
  wire g1955;
  wire g19552;
  wire g19553;
  wire g19554;
  wire g19558;
  wire g19559;
  wire g19565;
  wire g19566;
  wire g19567;
  wire g19569;
  wire g19570;
  wire g19573;
  wire g19574;
  wire g19577;
  wire g19579;
  wire g19580;
  wire g19586;
  wire g1959;
  wire g19600;
  wire g19602;
  wire g19603;
  wire g19606;
  wire g19612;
  wire g19617;
  wire g19618;
  wire g19620;
  wire g19626;
  wire g19629;
  wire g19630;
  wire g19633;
  wire g19634;
  wire g19635;
  wire g19636;
  wire g19638;
  wire g1964;
  wire g19644;
  wire g19649;
  wire g19650;
  wire g19652;
  wire g19653;
  wire g19654;
  wire g19657;
  wire g19658;
  wire g19659;
  wire g19662;
  wire g19666;
  wire g19670;
  wire g19672;
  wire g19673;
  wire g19675;
  wire g19676;
  wire g19677;
  wire g19678;
  wire g19679;
  wire g1968;
  wire g19682;
  wire g19683;
  wire g19685;
  wire g19686;
  wire g19687;
  wire g19688;
  wire g19689;
  wire g19690;
  wire g19694;
  wire g19695;
  wire g19696;
  wire g19697;
  wire g19698;
  wire g19709;
  wire g19710;
  wire g19711;
  wire g19712;
  wire g19713;
  wire g19714;
  wire g19718;
  wire g19719;
  wire g19730;
  wire g19731;
  wire g19732;
  wire g19733;
  wire g19734;
  wire g19737;
  wire g19739;
  wire g1974;
  wire g19741;
  wire g19742;
  wire g19743;
  wire g19744;
  wire g19745;
  wire g19747;
  wire g19748;
  wire g19750;
  wire g19753;
  wire g19754;
  wire g19755;
  wire g19757;
  wire g19760;
  wire g19761;
  wire g19762;
  wire g19763;
  wire g19765;
  wire g19766;
  wire g19769;
  wire g19770;
  wire g19771;
  wire g19772;
  wire g19773;
  wire g19776;
  wire g19777;
  wire g19779;
  wire g1978;
  wire g19780;
  wire g19781;
  wire g19783;
  wire g19785;
  wire g19786;
  wire g19787;
  wire g19789;
  wire g19790;
  wire g19794;
  wire g19798;
  wire g19799;
  wire g19800;
  wire g1982;
  wire g19852;
  wire g19860;
  wire g19861;
  wire g19862;
  wire g19865;
  wire g19872;
  wire g19878;
  wire g1988;
  wire g19881;
  wire g19885;
  wire g199;
  wire g19902;
  wire g19905;
  wire g19912;
  wire g19915;
  wire g1992;
  wire g19930;
  wire g19931;
  wire g19947;
  wire g19950;
  wire g19952;
  wire g1996;
  wire g19960;
  wire g19961;
  wire g19963;
  wire g19964;
  wire g19979;
  wire g19980;
  wire g19996;
  wire g19998;
  wire g20004;
  wire g20005;
  wire g20006;
  wire g20008;
  wire g20009;
  wire g20010;
  wire g20025;
  wire g20026;
  wire g20028;
  wire g20036;
  wire g20037;
  wire g20038;
  wire g2004;
  wire g20040;
  wire g20041;
  output g20049;
  wire g20050;
  wire g20052;
  wire g20053;
  wire g20054;
  wire g20057;
  wire g20058;
  wire g20059;
  wire g20064;
  wire g20066;
  wire g20067;
  wire g20071;
  wire g20072;
  wire g20079;
  wire g2008;
  wire g20080;
  wire g20087;
  wire g20088;
  wire g20089;
  wire g20090;
  wire g20091;
  wire g20096;
  wire g20097;
  wire g20101;
  wire g20102;
  wire g20103;
  wire g20104;
  wire g20105;
  wire g20106;
  wire g20110;
  wire g20113;
  wire g2012;
  wire g20128;
  wire g20129;
  wire g20130;
  wire g20132;
  wire g20144;
  wire g20145;
  wire g20146;
  wire g20147;
  wire g20153;
  wire g20157;
  wire g20158;
  wire g20159;
  wire g2016;
  wire g20164;
  wire g20166;
  wire g20167;
  wire g20168;
  wire g20178;
  wire g20179;
  wire g20180;
  wire g20182;
  wire g20190;
  wire g20191;
  wire g20194;
  wire g20195;
  wire g20197;
  wire g2020;
  wire g20204;
  wire g20207;
  wire g20208;
  wire g20209;
  wire g20210;
  wire g20211;
  wire g20213;
  wire g20229;
  wire g20231;
  wire g20232;
  wire g20233;
  wire g20235;
  wire g20238;
  wire g20239;
  wire g2024;
  wire g20240;
  wire g20242;
  wire g20247;
  wire g20265;
  wire g20266;
  wire g20267;
  wire g20268;
  wire g20270;
  wire g20273;
  wire g20274;
  wire g20275;
  wire g20277;
  wire g2028;
  wire g203;
  wire g20320;
  wire g20321;
  wire g20322;
  wire g20323;
  wire g20324;
  wire g20325;
  wire g20326;
  wire g20327;
  wire g20329;
  wire g2036;
  wire g20372;
  wire g20373;
  wire g20374;
  wire g20379;
  wire g20380;
  wire g20381;
  wire g20382;
  wire g20383;
  wire g20384;
  wire g20385;
  wire g20386;
  wire g20387;
  wire g20389;
  wire g2040;
  wire g20432;
  wire g20433;
  wire g20434;
  wire g20435;
  wire g20441;
  wire g20442;
  wire g20443;
  wire g20444;
  wire g20445;
  wire g20446;
  wire g20447;
  wire g20448;
  wire g20449;
  wire g20450;
  wire g20451;
  wire g20452;
  wire g2047;
  wire g20494;
  wire g20495;
  wire g20496;
  wire g20497;
  wire g20498;
  wire g20499;
  wire g20500;
  wire g20501;
  wire g20502;
  wire g20503;
  wire g20504;
  wire g20505;
  wire g20506;
  wire g20507;
  wire g20508;
  wire g20509;
  wire g2051;
  wire g20510;
  wire g20511;
  wire g20512;
  wire g20513;
  wire g20514;
  wire g20515;
  wire g20523;
  wire g20524;
  wire g20525;
  wire g20526;
  wire g20527;
  wire g20528;
  wire g20529;
  wire g20530;
  wire g20532;
  wire g20533;
  wire g20534;
  wire g20535;
  wire g20536;
  wire g20537;
  wire g20538;
  wire g20539;
  wire g20541;
  wire g20542;
  wire g20543;
  wire g20544;
  wire g20545;
  wire g20546;
  wire g20547;
  wire g20548;
  wire g20549;
  wire g20551;
  wire g20552;
  wire g20553;
  wire g20554;
  wire g20555;
  wire g20556;
  output g20557;
  wire g20558;
  wire g20560;
  wire g20561;
  wire g20562;
  wire g20563;
  wire g20564;
  wire g20565;
  wire g20566;
  wire g20567;
  wire g20568;
  wire g20569;
  wire g20570;
  wire g20571;
  wire g20573;
  wire g20574;
  wire g20575;
  wire g20576;
  wire g20577;
  wire g20578;
  wire g20579;
  wire g20580;
  wire g20582;
  wire g20583;
  wire g20584;
  wire g20585;
  wire g20586;
  wire g20587;
  wire g20588;
  wire g20589;
  wire g20590;
  wire g20591;
  wire g20592;
  wire g20593;
  wire g20594;
  wire g20597;
  wire g20598;
  wire g20599;
  wire g2060;
  wire g20600;
  wire g20601;
  wire g20603;
  wire g20604;
  wire g20605;
  wire g20606;
  wire g20607;
  wire g20608;
  wire g20609;
  wire g20610;
  wire g20611;
  wire g20612;
  wire g20613;
  wire g20614;
  wire g20615;
  wire g20616;
  wire g20617;
  wire g20618;
  wire g20622;
  wire g20623;
  wire g20624;
  wire g20625;
  wire g20626;
  wire g20627;
  wire g20629;
  wire g20630;
  wire g20631;
  wire g20632;
  wire g20633;
  wire g20634;
  wire g20635;
  wire g20636;
  wire g20637;
  wire g20638;
  wire g20639;
  wire g20640;
  wire g20641;
  wire g20642;
  wire g20648;
  wire g20649;
  wire g20650;
  wire g20651;
  output g20652;
  wire g20653;
  output g20654;
  wire g20655;
  wire g20656;
  wire g20657;
  wire g20659;
  wire g2066;
  wire g20660;
  wire g20661;
  wire g20662;
  wire g20663;
  wire g20664;
  wire g20665;
  wire g20666;
  wire g20667;
  wire g20668;
  wire g20669;
  wire g20670;
  wire g20671;
  wire g20672;
  wire g20673;
  wire g20674;
  wire g20679;
  wire g20680;
  wire g20681;
  wire g20682;
  wire g20695;
  wire g20696;
  wire g20697;
  wire g20698;
  wire g20699;
  wire g2070;
  wire g20700;
  wire g20701;
  wire g20702;
  wire g20703;
  wire g20704;
  wire g20706;
  wire g20707;
  wire g20708;
  wire g20709;
  wire g20710;
  wire g20711;
  wire g20712;
  wire g20713;
  wire g20714;
  wire g20715;
  wire g20716;
  wire g20732;
  wire g20737;
  wire g20738;
  output g20763;
  wire g20764;
  wire g20766;
  wire g20767;
  wire g20768;
  wire g20769;
  wire g20770;
  wire g20771;
  wire g20772;
  wire g20774;
  wire g20775;
  wire g20776;
  wire g20777;
  wire g20778;
  wire g20779;
  wire g20780;
  wire g2079;
  wire g2084;
  wire g20852;
  wire g20853;
  wire g20869;
  wire g20874;
  wire g2089;
  output g20899;
  wire g209;
  wire g20900;
  output g20901;
  wire g20902;
  wire g20903;
  wire g20904;
  wire g20909;
  wire g20910;
  wire g20911;
  wire g20912;
  wire g20913;
  wire g20914;
  wire g20916;
  wire g20917;
  wire g20918;
  wire g20919;
  wire g20920;
  wire g20921;
  wire g20923;
  wire g2093;
  wire g20978;
  wire g2098;
  wire g20993;
  wire g20994;
  wire g21010;
  wire g2102;
  wire g21036;
  wire g21048;
  wire g21049;
  wire g21050;
  wire g21051;
  wire g21052;
  wire g21053;
  wire g21054;
  wire g21055;
  wire g21056;
  wire g21057;
  wire g21058;
  wire g21059;
  wire g21060;
  wire g21068;
  wire g21069;
  wire g2108;
  wire g2112;
  wire g21123;
  wire g21138;
  wire g21139;
  wire g21155;
  wire g21156;
  wire g2116;
  wire g21160;
  wire g21175;
  output g21176;
  wire g21177;
  wire g21178;
  wire g21179;
  wire g21180;
  wire g21181;
  wire g21182;
  wire g21183;
  wire g21184;
  wire g21185;
  wire g21189;
  wire g21204;
  wire g21205;
  wire g2122;
  wire g21221;
  wire g21222;
  wire g21225;
  wire g21228;
  output g21245;
  wire g21246;
  wire g21247;
  wire g21248;
  wire g21249;
  wire g21252;
  wire g2126;
  wire g21267;
  wire g21268;
  wire g21269;
  output g21270;
  wire g21271;
  wire g21274;
  wire g21275;
  wire g21279;
  wire g21281;
  wire g21282;
  wire g21286;
  wire g21291;
  output g21292;
  wire g21293;
  wire g21295;
  wire g21299;
  wire g2130;
  wire g21300;
  wire g21304;
  wire g21305;
  wire g21308;
  wire g21329;
  wire g21336;
  wire g21337;
  wire g21343;
  wire g21346;
  wire g21349;
  wire g21352;
  wire g21355;
  wire g21358;
  wire g21362;
  wire g21366;
  wire g21369;
  wire g21370;
  wire g21379;
  wire g2138;
  wire g21380;
  wire g21381;
  wire g21383;
  wire g21395;
  wire g21396;
  wire g21397;
  wire g21398;
  wire g21399;
  wire g21400;
  wire g21406;
  wire g21407;
  wire g21408;
  wire g21409;
  wire g21410;
  wire g21411;
  wire g21412;
  wire g21414;
  wire g21418;
  wire g21421;
  wire g21422;
  wire g21423;
  wire g21424;
  wire g21425;
  wire g21426;
  wire g21427;
  wire g21428;
  wire g21431;
  wire g21434;
  wire g2145;
  wire g21451;
  wire g21454;
  wire g21455;
  wire g21456;
  wire g21457;
  wire g21458;
  wire g21461;
  wire g21463;
  wire g21466;
  wire g21467;
  wire g215;
  wire g2151;
  wire g21511;
  wire g2152;
  wire g2153;
  wire g21560;
  wire g21561;
  wire g21604;
  wire g21607;
  wire g21608;
  wire g21609;
  wire g2161;
  wire g21610;
  wire g2165;
  wire g21665;
  wire g21669;
  wire g21673;
  wire g21677;
  wire g21681;
  wire g21685;
  wire g21689;
  wire g2169;
  wire g21693;
  wire g21697;
  output g21698;
  wire g21722;
  wire g21723;
  wire g21724;
  wire g21725;
  wire g21726;
  output g21727;
  wire g2173;
  wire g2177;
  wire g218;
  wire g2181;
  wire g2185;
  wire g21891;
  wire g21892;
  wire g21893;
  wire g21894;
  wire g21895;
  wire g21896;
  wire g21897;
  wire g21898;
  wire g21899;
  wire g21900;
  wire g21901;
  wire g21902;
  wire g21903;
  wire g21904;
  wire g21905;
  wire g2193;
  wire g2197;
  wire g22;
  wire g2204;
  wire g2208;
  wire g22144;
  wire g22146;
  wire g22147;
  wire g22148;
  wire g22153;
  wire g22154;
  wire g22155;
  wire g22156;
  wire g22166;
  wire g22167;
  wire g22168;
  wire g22169;
  wire g2217;
  wire g22170;
  wire g22173;
  wire g22176;
  wire g22177;
  wire g22178;
  wire g22179;
  wire g22180;
  wire g22181;
  wire g22182;
  wire g22192;
  wire g22194;
  wire g22197;
  wire g22198;
  wire g22199;
  wire g222;
  wire g22200;
  wire g22201;
  wire g22202;
  wire g22210;
  wire g22213;
  wire g22214;
  wire g22215;
  wire g22220;
  wire g22223;
  wire g22224;
  wire g22227;
  wire g2223;
  wire g2227;
  wire g22300;
  wire g22303;
  wire g22305;
  wire g22317;
  wire g22330;
  wire g22338;
  wire g22339;
  wire g22341;
  wire g22358;
  wire g2236;
  wire g22360;
  wire g22409;
  wire g2241;
  wire g22455;
  wire g22456;
  wire g2246;
  wire g22493;
  wire g22494;
  wire g22495;
  wire g225;
  wire g2250;
  wire g22519;
  wire g22520;
  wire g22526;
  wire g22528;
  wire g22542;
  wire g22543;
  wire g2255;
  wire g2259;
  wire g22593;
  wire g22635;
  wire g22647;
  wire g2265;
  wire g22658;
  wire g22683;
  wire g2269;
  wire g22698;
  wire g22721;
  wire g2273;
  wire g22758;
  wire g22763;
  wire g2279;
  wire g2283;
  wire g22830;
  wire g22840;
  wire g22841;
  wire g22847;
  wire g22854;
  wire g22855;
  wire g22856;
  wire g22865;
  wire g22866;
  wire g22867;
  wire g22868;
  wire g2287;
  wire g22882;
  wire g22883;
  wire g22884;
  wire g22898;
  wire g22903;
  wire g22906;
  wire g22907;
  wire g22922;
  wire g22923;
  wire g22926;
  wire g22935;
  wire g22936;
  wire g2295;
  wire g22973;
  wire g22974;
  wire g22975;
  wire g22976;
  wire g22979;
  wire g22981;
  wire g22985;
  wire g22986;
  wire g22987;
  wire g22988;
  wire g22989;
  wire g2299;
  wire g22995;
  wire g22996;
  wire g22997;
  wire g22998;
  wire g22999;
  wire g23000;
  wire g23001;
  output g23002;
  wire g23003;
  wire g23004;
  wire g23005;
  wire g23011;
  wire g23012;
  wire g23013;
  wire g23014;
  wire g23015;
  wire g23016;
  wire g23017;
  wire g23018;
  wire g23019;
  wire g23020;
  wire g23021;
  wire g23022;
  wire g23026;
  wire g23027;
  wire g23028;
  wire g23029;
  wire g2303;
  wire g23030;
  wire g23031;
  wire g23032;
  wire g23041;
  wire g23046;
  wire g23057;
  wire g23058;
  wire g23059;
  wire g23060;
  wire g23061;
  wire g23066;
  wire g2307;
  wire g23084;
  wire g23085;
  wire g23086;
  wire g2311;
  wire g23111;
  wire g23128;
  wire g23138;
  wire g2315;
  wire g23152;
  wire g23170;
  wire g23189;
  wire g2319;
  output g23190;
  wire g23191;
  wire g23196;
  wire g232;
  wire g23203;
  wire g23214;
  wire g23215;
  wire g23216;
  wire g23221;
  wire g23222;
  wire g23226;
  wire g23227;
  wire g23228;
  wire g23232;
  wire g23233;
  wire g23235;
  wire g23236;
  wire g23237;
  wire g23238;
  wire g23242;
  wire g23243;
  wire g23245;
  wire g23246;
  wire g23247;
  wire g23248;
  wire g23249;
  wire g23250;
  wire g23253;
  wire g23256;
  wire g23257;
  wire g23258;
  wire g23259;
  wire g23260;
  wire g23263;
  wire g23264;
  wire g2327;
  wire g23270;
  wire g23271;
  wire g23272;
  wire g23273;
  wire g23274;
  wire g23277;
  wire g23278;
  wire g23279;
  wire g23282;
  wire g23283;
  wire g23284;
  wire g23289;
  wire g23290;
  wire g23291;
  wire g23299;
  wire g23300;
  wire g23301;
  wire g23302;
  wire g23303;
  wire g23304;
  wire g23305;
  wire g23306;
  wire g23307;
  wire g2331;
  wire g23312;
  wire g23313;
  wire g23320;
  wire g23321;
  wire g23322;
  wire g23323;
  wire g23332;
  wire g23333;
  wire g23334;
  wire g23335;
  wire g23336;
  wire g23337;
  wire g23338;
  wire g23339;
  wire g23340;
  wire g23347;
  wire g23350;
  wire g23351;
  wire g23352;
  wire g23353;
  wire g23354;
  wire g23355;
  wire g23356;
  wire g23359;
  wire g23360;
  wire g23361;
  wire g23362;
  wire g23375;
  wire g23376;
  wire g23377;
  wire g23378;
  wire g2338;
  wire g23384;
  wire g23385;
  wire g23388;
  wire g23390;
  wire g23394;
  wire g23395;
  wire g23398;
  wire g23399;
  wire g23403;
  wire g23406;
  wire g23408;
  wire g23409;
  wire g23410;
  wire g23414;
  wire g23417;
  wire g23418;
  wire g23419;
  wire g2342;
  wire g23420;
  wire g23421;
  wire g23422;
  wire g23426;
  wire g23427;
  wire g23429;
  wire g23431;
  wire g23432;
  wire g23433;
  wire g23434;
  wire g23435;
  wire g23440;
  wire g23443;
  wire g23446;
  wire g23447;
  wire g23448;
  wire g23449;
  wire g23450;
  wire g23452;
  wire g23453;
  wire g23456;
  wire g23459;
  wire g23460;
  wire g23461;
  wire g23473;
  wire g23476;
  wire g23477;
  wire g23478;
  wire g23479;
  wire g23482;
  wire g23483;
  wire g23485;
  wire g23486;
  wire g23487;
  wire g23488;
  wire g23489;
  wire g23490;
  wire g23491;
  wire g23492;
  wire g23493;
  wire g23499;
  wire g23500;
  wire g23501;
  wire g23502;
  wire g23503;
  wire g23504;
  wire g23505;
  wire g23506;
  wire g23507;
  wire g23508;
  wire g23509;
  wire g2351;
  wire g23510;
  wire g23515;
  wire g23516;
  wire g23517;
  wire g23518;
  wire g23519;
  wire g23520;
  wire g23521;
  wire g23522;
  wire g23523;
  wire g23524;
  wire g23525;
  wire g23526;
  wire g23527;
  wire g23528;
  wire g23534;
  wire g23537;
  wire g23538;
  wire g23539;
  wire g23541;
  wire g23542;
  wire g23543;
  wire g23544;
  wire g23545;
  wire g23546;
  wire g23547;
  wire g23548;
  wire g23549;
  wire g23555;
  wire g23558;
  wire g23559;
  wire g23565;
  wire g23566;
  wire g23567;
  wire g23568;
  wire g23569;
  wire g2357;
  wire g23570;
  wire g23571;
  wire g23582;
  wire g23585;
  wire g23589;
  wire g23607;
  wire g23608;
  wire g23609;
  wire g2361;
  wire g23610;
  wire g23611;
  output g23612;
  wire g23613;
  wire g23629;
  wire g23647;
  wire g23648;
  wire g23649;
  output g23652;
  wire g23653;
  wire g23665;
  output g23683;
  wire g23684;
  wire g23698;
  wire g2370;
  wire g23732;
  wire g23749;
  wire g2375;
  output g23759;
  wire g23760;
  wire g23767;
  wire g23768;
  wire g23769;
  wire g23777;
  wire g23787;
  wire g23788;
  wire g23792;
  wire g23793;
  wire g23794;
  wire g2380;
  wire g23812;
  wire g23813;
  wire g23814;
  wire g23815;
  wire g23819;
  wire g23820;
  wire g23821;
  wire g23823;
  wire g23838;
  wire g23839;
  wire g2384;
  wire g23840;
  wire g23841;
  wire g23842;
  wire g23843;
  wire g23847;
  wire g23848;
  wire g23849;
  wire g23858;
  wire g23859;
  wire g23860;
  wire g23861;
  wire g23862;
  wire g23863;
  wire g23864;
  wire g23868;
  wire g23869;
  wire g23870;
  wire g23874;
  wire g23875;
  wire g23876;
  wire g23877;
  wire g23878;
  wire g23879;
  wire g23880;
  wire g23881;
  wire g23882;
  wire g23886;
  wire g23887;
  wire g23888;
  wire g2389;
  wire g23893;
  wire g23894;
  wire g23895;
  wire g23896;
  wire g23897;
  wire g23898;
  wire g23899;
  wire g239;
  wire g23902;
  wire g23903;
  wire g23904;
  wire g23905;
  wire g23906;
  wire g23907;
  wire g23912;
  wire g23913;
  wire g23914;
  wire g23915;
  wire g23916;
  wire g23922;
  wire g23923;
  wire g23924;
  wire g23925;
  wire g23926;
  wire g23927;
  wire g23928;
  wire g23929;
  wire g2393;
  wire g23930;
  wire g23935;
  wire g23936;
  wire g23937;
  wire g23938;
  wire g23939;
  wire g23940;
  wire g23941;
  wire g23942;
  wire g23943;
  wire g23944;
  wire g23945;
  wire g23946;
  wire g23947;
  wire g23952;
  wire g23953;
  wire g23954;
  wire g23961;
  wire g23962;
  wire g23963;
  wire g23964;
  wire g23965;
  wire g23966;
  wire g23967;
  wire g23968;
  wire g23969;
  wire g23970;
  wire g23982;
  wire g23983;
  wire g23984;
  wire g23985;
  wire g23986;
  wire g23987;
  wire g23988;
  wire g2399;
  wire g23992;
  wire g23993;
  wire g23994;
  wire g23995;
  wire g23999;
  wire g24000;
  wire g24003;
  wire g24010;
  wire g24013;
  wire g24017;
  wire g2403;
  wire g2407;
  wire g2413;
  output g24151;
  wire g24152;
  wire g24153;
  wire g24154;
  wire g24155;
  wire g24156;
  wire g24157;
  wire g24158;
  wire g24159;
  wire g24160;
  output g24161;
  output g24162;
  output g24163;
  output g24164;
  output g24165;
  output g24166;
  output g24167;
  output g24168;
  output g24169;
  wire g2417;
  output g24170;
  output g24171;
  output g24172;
  output g24173;
  output g24174;
  output g24175;
  output g24176;
  output g24177;
  output g24178;
  output g24179;
  output g24180;
  output g24181;
  output g24182;
  output g24183;
  output g24184;
  output g24185;
  wire g24200;
  wire g24201;
  wire g24202;
  wire g24203;
  wire g24204;
  wire g24205;
  wire g24206;
  wire g24207;
  wire g24208;
  wire g24209;
  wire g2421;
  wire g24210;
  wire g24211;
  wire g24212;
  wire g24213;
  wire g24214;
  wire g24215;
  wire g24216;
  wire g24229;
  wire g24231;
  wire g24232;
  wire g24233;
  wire g24234;
  wire g24235;
  wire g24236;
  wire g24237;
  wire g24238;
  wire g24239;
  wire g24240;
  wire g24241;
  wire g24242;
  wire g24243;
  wire g24244;
  wire g24245;
  wire g24246;
  wire g24247;
  wire g24248;
  wire g24249;
  wire g24250;
  wire g24251;
  wire g24252;
  wire g24253;
  wire g24254;
  wire g24255;
  wire g24256;
  wire g24257;
  wire g24258;
  wire g24259;
  wire g24260;
  wire g24261;
  wire g24262;
  wire g24263;
  wire g24264;
  wire g24265;
  wire g24266;
  wire g24267;
  wire g24268;
  wire g24269;
  wire g24270;
  wire g24271;
  wire g24272;
  wire g24273;
  wire g24274;
  wire g24275;
  wire g24276;
  wire g24277;
  wire g24278;
  wire g24279;
  wire g24280;
  wire g24281;
  wire g24282;
  wire g2429;
  wire g24298;
  wire g2433;
  wire g24334;
  wire g24335;
  wire g24336;
  wire g24337;
  wire g24338;
  wire g24339;
  wire g24340;
  wire g24341;
  wire g24342;
  wire g24343;
  wire g24344;
  wire g24345;
  wire g24346;
  wire g24347;
  wire g24348;
  wire g24349;
  wire g24350;
  wire g24351;
  wire g24352;
  wire g24353;
  wire g24354;
  wire g24355;
  wire g24356;
  wire g24358;
  wire g24359;
  wire g24360;
  wire g24364;
  wire g24365;
  wire g24366;
  wire g24367;
  wire g24368;
  wire g2437;
  wire g24375;
  wire g24376;
  wire g24377;
  wire g24379;
  wire g24386;
  wire g24394;
  wire g24405;
  wire g24407;
  wire g2441;
  wire g24417;
  wire g24418;
  wire g24419;
  wire g24424;
  wire g24425;
  wire g24426;
  wire g24428;
  wire g24429;
  wire g24431;
  wire g24438;
  wire g2445;
  wire g24452;
  wire g2449;
  wire g24490;
  wire g2453;
  wire g24575;
  wire g246;
  wire g2461;
  wire g24619;
  wire g2465;
  wire g2472;
  wire g24759;
  wire g2476;
  wire g24819;
  wire g24836;
  wire g2485;
  wire g24850;
  wire g24866;
  wire g24869;
  wire g24891;
  wire g24893;
  wire g2491;
  wire g24911;
  wire g24920;
  wire g2495;
  wire g25027;
  wire g2504;
  wire g25051;
  wire g25064;
  wire g25067;
  wire g25073;
  wire g25084;
  wire g25085;
  wire g2509;
  wire g25102;
  wire g25103;
  output g25114;
  wire g25115;
  wire g25123;
  wire g25124;
  wire g2514;
  wire g25140;
  wire g25142;
  wire g25143;
  wire g25158;
  wire g25159;
  output g25167;
  wire g25168;
  wire g25171;
  wire g2518;
  wire g25180;
  wire g25185;
  wire g25198;
  wire g25206;
  wire g25214;
  output g25219;
  wire g25220;
  wire g25221;
  wire g25222;
  wire g2523;
  wire g25231;
  wire g25232;
  wire g25240;
  wire g25241;
  wire g25248;
  wire g25249;
  wire g25250;
  output g25259;
  wire g25260;
  wire g25266;
  wire g25267;
  wire g2527;
  wire g25272;
  wire g25286;
  wire g25287;
  wire g25288;
  wire g25289;
  wire g25296;
  wire g25297;
  wire g25298;
  wire g25324;
  wire g25325;
  wire g25326;
  wire g2533;
  wire g25369;
  wire g2537;
  wire g25370;
  wire g25380;
  wire g25409;
  wire g2541;
  wire g25410;
  wire g25423;
  wire g25424;
  wire g25448;
  wire g25451;
  wire g25452;
  wire g25465;
  wire g2547;
  wire g25480;
  wire g25481;
  wire g255;
  wire g25505;
  wire g25506;
  wire g2551;
  wire g25513;
  wire g25517;
  wire g25523;
  wire g25524;
  wire g25525;
  wire g25528;
  wire g25531;
  wire g25533;
  wire g25537;
  wire g25538;
  wire g25544;
  wire g25546;
  wire g25547;
  wire g25548;
  wire g2555;
  wire g25552;
  wire g25553;
  wire g25554;
  wire g25555;
  wire g25558;
  wire g25560;
  wire g25561;
  wire g25563;
  wire g25566;
  output g25582;
  output g25583;
  output g25584;
  output g25585;
  output g25586;
  output g25587;
  output g25588;
  output g25589;
  output g25590;
  wire g25591;
  wire g25592;
  wire g25593;
  wire g25594;
  wire g25595;
  wire g25596;
  wire g25597;
  wire g25598;
  wire g25599;
  wire g25600;
  wire g25601;
  wire g25602;
  wire g25603;
  wire g25604;
  wire g25605;
  wire g25606;
  wire g25607;
  wire g25608;
  wire g25609;
  wire g25610;
  wire g25611;
  wire g25612;
  wire g25613;
  wire g25614;
  wire g25615;
  wire g25616;
  wire g25617;
  wire g25618;
  wire g25619;
  wire g25620;
  wire g25621;
  wire g25622;
  wire g25623;
  wire g25624;
  wire g25625;
  wire g25626;
  wire g25627;
  wire g25628;
  wire g25629;
  wire g2563;
  wire g25630;
  wire g25631;
  wire g25632;
  wire g25633;
  wire g25634;
  wire g25635;
  wire g25636;
  wire g25637;
  wire g25638;
  wire g25639;
  wire g25640;
  wire g25641;
  wire g25642;
  wire g25643;
  wire g25644;
  wire g25645;
  wire g25646;
  wire g25647;
  wire g25648;
  wire g25649;
  wire g25650;
  wire g25651;
  wire g25652;
  wire g25653;
  wire g25654;
  wire g25655;
  wire g25656;
  wire g25657;
  wire g25658;
  wire g25659;
  wire g25660;
  wire g25661;
  wire g25662;
  wire g25663;
  wire g25664;
  wire g25665;
  wire g25666;
  wire g25667;
  wire g25668;
  wire g25669;
  wire g2567;
  wire g25670;
  wire g25671;
  wire g25672;
  wire g25673;
  wire g25674;
  wire g25675;
  wire g25676;
  wire g25677;
  wire g25678;
  wire g25679;
  wire g25680;
  wire g25681;
  wire g25682;
  wire g25683;
  wire g25684;
  wire g25685;
  wire g25686;
  wire g25687;
  wire g25688;
  wire g25689;
  wire g25690;
  wire g25691;
  wire g25692;
  wire g25693;
  wire g25694;
  wire g25695;
  wire g25696;
  wire g25697;
  wire g25698;
  wire g25699;
  wire g25700;
  wire g25701;
  wire g25702;
  wire g25703;
  wire g25704;
  wire g25705;
  wire g25706;
  wire g25707;
  wire g25708;
  wire g25709;
  wire g2571;
  wire g25710;
  wire g25711;
  wire g25712;
  wire g25713;
  wire g25714;
  wire g25715;
  wire g25716;
  wire g25717;
  wire g25718;
  wire g25719;
  wire g25720;
  wire g25721;
  wire g25722;
  wire g25723;
  wire g25724;
  wire g25725;
  wire g25726;
  wire g25727;
  wire g25728;
  wire g25729;
  wire g25730;
  wire g25731;
  wire g25732;
  wire g25733;
  wire g25734;
  wire g25735;
  wire g25736;
  wire g25737;
  wire g25738;
  wire g25739;
  wire g25740;
  wire g25741;
  wire g25742;
  wire g25743;
  wire g25744;
  wire g25745;
  wire g25746;
  wire g25747;
  wire g25748;
  wire g25749;
  wire g2575;
  wire g25750;
  wire g25751;
  wire g25752;
  wire g25753;
  wire g25754;
  wire g25755;
  wire g25756;
  wire g25757;
  wire g25758;
  wire g25759;
  wire g25760;
  wire g25761;
  wire g25762;
  wire g25763;
  wire g25764;
  wire g25768;
  wire g25771;
  wire g25775;
  wire g25782;
  wire g2579;
  wire g2583;
  wire g25831;
  wire g25850;
  wire g25866;
  wire g2587;
  wire g25903;
  wire g2595;
  wire g25986;
  wire g2599;
  wire g26019;
  wire g26048;
  wire g2606;
  wire g26079;
  wire g26088;
  wire g2610;
  wire g26105;
  wire g26131;
  wire g26187;
  wire g2619;
  wire g262;
  wire g2625;
  wire g26257;
  wire g26260;
  wire g26274;
  wire g26279;
  wire g26287;
  wire g2629;
  wire g26292;
  wire g26294;
  wire g26301;
  wire g26304;
  wire g26312;
  wire g26337;
  wire g2638;
  wire g2643;
  wire g2648;
  wire g26510;
  wire g2652;
  wire g2657;
  wire g2661;
  wire g2667;
  wire g2671;
  wire g2675;
  output g26801;
  wire g26802;
  wire g2681;
  wire g26811;
  wire g26814;
  wire g26817;
  wire g26818;
  wire g26820;
  wire g26824;
  wire g26825;
  wire g26829;
  wire g26833;
  wire g26834;
  wire g26835;
  wire g26838;
  wire g26839;
  wire g26840;
  wire g26842;
  wire g26843;
  wire g26846;
  wire g26847;
  wire g26848;
  wire g26849;
  wire g2685;
  wire g26850;
  wire g26851;
  wire g26853;
  wire g26854;
  wire g26855;
  wire g26856;
  wire g26858;
  wire g26859;
  wire g26860;
  wire g26862;
  wire g26864;
  wire g26869;
  wire g26870;
  output g26875;
  output g26876;
  output g26877;
  wire g26880;
  wire g26881;
  wire g26882;
  wire g26883;
  wire g26884;
  wire g26885;
  wire g26886;
  wire g26887;
  wire g26888;
  wire g26889;
  wire g2689;
  wire g26890;
  wire g26891;
  wire g26892;
  wire g26893;
  wire g26894;
  wire g26895;
  wire g26896;
  wire g26897;
  wire g26898;
  wire g26899;
  wire g269;
  wire g26900;
  wire g26901;
  wire g26902;
  wire g26903;
  wire g26904;
  wire g26905;
  wire g26906;
  wire g26907;
  wire g26908;
  wire g26909;
  wire g26910;
  wire g26911;
  wire g26912;
  wire g26913;
  wire g26914;
  wire g26915;
  wire g26916;
  wire g26917;
  wire g26918;
  wire g26919;
  wire g26920;
  wire g26921;
  wire g26922;
  wire g26923;
  wire g26924;
  wire g26925;
  wire g26926;
  wire g26927;
  wire g26928;
  wire g26929;
  wire g26930;
  wire g26931;
  wire g26932;
  wire g26933;
  wire g26934;
  wire g26935;
  wire g26936;
  wire g26937;
  wire g26938;
  wire g26939;
  wire g26940;
  wire g26941;
  wire g26942;
  wire g26943;
  wire g26944;
  wire g26945;
  wire g26946;
  wire g26947;
  wire g26948;
  wire g26949;
  wire g26950;
  wire g26951;
  wire g26952;
  wire g26953;
  wire g26954;
  wire g26955;
  wire g26956;
  wire g26957;
  wire g26958;
  wire g26959;
  wire g26960;
  wire g26961;
  wire g26962;
  wire g26963;
  wire g26964;
  wire g26965;
  wire g26966;
  wire g26967;
  wire g26968;
  wire g26969;
  wire g2697;
  wire g26970;
  wire g26971;
  wire g27013;
  wire g2704;
  wire g2710;
  wire g2711;
  wire g2712;
  wire g27121;
  wire g2715;
  wire g2719;
  wire g2724;
  wire g2729;
  wire g27320;
  wire g2735;
  wire g2741;
  wire g27438;
  wire g2748;
  wire g27511;
  wire g27527;
  wire g2756;
  wire g27576;
  wire g27585;
  wire g2759;
  wire g2763;
  wire g27662;
  wire g2767;
  wire g27675;
  wire g27678;
  wire g27686;
  wire g27698;
  wire g27708;
  wire g27709;
  wire g2771;
  wire g27736;
  wire g27737;
  wire g2775;
  wire g27765;
  wire g27773;
  wire g27774;
  wire g2779;
  wire g278;
  wire g27822;
  wire g2783;
  output g27831;
  wire g27832;
  wire g2787;
  wire g27880;
  wire g27881;
  wire g2791;
  wire g27928;
  wire g27929;
  wire g27930;
  wire g2795;
  wire g27956;
  wire g27961;
  wire g27967;
  wire g2799;
  wire g27993;
  wire g27996;
  wire g27998;
  wire g28;
  wire g28009;
  wire g2803;
  output g28030;
  output g28041;
  output g28042;
  wire g28043;
  wire g28044;
  wire g28045;
  wire g28046;
  wire g28047;
  wire g28048;
  wire g28049;
  wire g28050;
  wire g28051;
  wire g28052;
  wire g28053;
  wire g28054;
  wire g28055;
  wire g28056;
  wire g28057;
  wire g28058;
  wire g28059;
  wire g28060;
  wire g28061;
  wire g28062;
  wire g28063;
  wire g28064;
  wire g28065;
  wire g28066;
  wire g28067;
  wire g28068;
  wire g28069;
  wire g2807;
  wire g28070;
  wire g28071;
  wire g28072;
  wire g28073;
  wire g28074;
  wire g28075;
  wire g28076;
  wire g28077;
  wire g28078;
  wire g28079;
  wire g28080;
  wire g28081;
  wire g28082;
  wire g28083;
  wire g28084;
  wire g28085;
  wire g28086;
  wire g28087;
  wire g28088;
  wire g28089;
  wire g28090;
  wire g28091;
  wire g28092;
  wire g28093;
  wire g28094;
  wire g28095;
  wire g28096;
  wire g28097;
  wire g28098;
  wire g28099;
  wire g28100;
  wire g28101;
  wire g28102;
  wire g28103;
  wire g28104;
  wire g28105;
  wire g2811;
  wire g28142;
  wire g28147;
  wire g2815;
  wire g28155;
  wire g28156;
  wire g28157;
  wire g28161;
  wire g28162;
  wire g28163;
  wire g28166;
  wire g28173;
  wire g28181;
  wire g28184;
  wire g28187;
  wire g2819;
  wire g2823;
  wire g28262;
  wire g2827;
  wire g283;
  wire g2831;
  wire g2834;
  wire g28367;
  wire g2837;
  wire g2841;
  wire g2844;
  wire g2848;
  wire g2852;
  wire g2856;
  wire g2860;
  wire g2864;
  wire g28652;
  wire g2868;
  wire g287;
  wire g28709;
  wire g2873;
  wire g28752;
  output g28753;
  wire g28754;
  wire g28779;
  wire g2878;
  wire g28819;
  wire g2882;
  wire g2886;
  wire g2890;
  wire g28917;
  wire g2894;
  wire g28954;
  wire g2898;
  wire g29013;
  wire g2902;
  wire g29041;
  wire g29042;
  wire g29043;
  wire g2907;
  wire g291;
  wire g2912;
  wire g29147;
  wire g2917;
  wire g29185;
  wire g29194;
  wire g29195;
  wire g29209;
  output g29210;
  output g29211;
  output g29212;
  output g29213;
  output g29214;
  output g29215;
  output g29216;
  output g29217;
  output g29218;
  output g29219;
  wire g2922;
  output g29220;
  output g29221;
  wire g29222;
  wire g29223;
  wire g29224;
  wire g29225;
  wire g29226;
  wire g29227;
  wire g29228;
  wire g29229;
  wire g29230;
  wire g29231;
  wire g29232;
  wire g29233;
  wire g29234;
  wire g29235;
  wire g29236;
  wire g29237;
  wire g29238;
  wire g29239;
  wire g29240;
  wire g29241;
  wire g29242;
  wire g29243;
  wire g29244;
  wire g29245;
  wire g29246;
  wire g29247;
  wire g29248;
  wire g29249;
  wire g29250;
  wire g29251;
  wire g29252;
  wire g29253;
  wire g29254;
  wire g29255;
  wire g29256;
  wire g29257;
  wire g29258;
  wire g29259;
  wire g29260;
  wire g29261;
  wire g29262;
  wire g29263;
  wire g29264;
  wire g29265;
  wire g29266;
  wire g29267;
  wire g29268;
  wire g29269;
  wire g2927;
  wire g29270;
  wire g29271;
  wire g29272;
  wire g29273;
  wire g29274;
  wire g29275;
  wire g29276;
  wire g29277;
  wire g29278;
  wire g29279;
  wire g29280;
  wire g29281;
  wire g29282;
  wire g29283;
  wire g29284;
  wire g29285;
  wire g29286;
  wire g29287;
  wire g29288;
  wire g29289;
  wire g29290;
  wire g29291;
  wire g29292;
  wire g29293;
  wire g29294;
  wire g29295;
  wire g29296;
  wire g29297;
  wire g29298;
  wire g29299;
  wire g29300;
  wire g29301;
  wire g29302;
  wire g29303;
  wire g29304;
  wire g29305;
  wire g29306;
  wire g29307;
  wire g29308;
  wire g29309;
  wire g29317;
  wire g2932;
  wire g2936;
  wire g29368;
  wire g29371;
  wire g29374;
  wire g29379;
  wire g294;
  wire g2941;
  wire g2946;
  wire g29491;
  wire g29498;
  wire g2950;
  wire g2955;
  wire g2960;
  wire g2965;
  wire g2970;
  wire g29744;
  wire g2975;
  wire g298;
  wire g2980;
  wire g29814;
  wire g2984;
  wire g2988;
  wire g2994;
  wire g2999;
  wire g30012;
  wire g3003;
  wire g3004;
  wire g30072;
  wire g301;
  wire g3010;
  wire g30105;
  wire g30116;
  wire g30155;
  wire g3017;
  wire g30182;
  wire g3021;
  wire g30218;
  wire g30237;
  wire g3025;
  wire g3029;
  wire g30295;
  wire g30301;
  wire g30322;
  output g30327;
  output g30329;
  output g30330;
  output g30331;
  output g30332;
  wire g30333;
  wire g30334;
  wire g30335;
  wire g30336;
  wire g30337;
  wire g30338;
  wire g30339;
  wire g3034;
  wire g30340;
  wire g30341;
  wire g30342;
  wire g30343;
  wire g30344;
  wire g30345;
  wire g30346;
  wire g30347;
  wire g30348;
  wire g30349;
  wire g30350;
  wire g30351;
  wire g30352;
  wire g30353;
  wire g30354;
  wire g30355;
  wire g30356;
  wire g30357;
  wire g30358;
  wire g30359;
  wire g30360;
  wire g30361;
  wire g30362;
  wire g30363;
  wire g30364;
  wire g30365;
  wire g30366;
  wire g30367;
  wire g30368;
  wire g30369;
  wire g30370;
  wire g30371;
  wire g30372;
  wire g30373;
  wire g30374;
  wire g30375;
  wire g30376;
  wire g30377;
  wire g30378;
  wire g30379;
  wire g30380;
  wire g30381;
  wire g30382;
  wire g30383;
  wire g30384;
  wire g30385;
  wire g30386;
  wire g30387;
  wire g30388;
  wire g30389;
  wire g30390;
  wire g30391;
  wire g30392;
  wire g30393;
  wire g30394;
  wire g30395;
  wire g30396;
  wire g30397;
  wire g30398;
  wire g30399;
  wire g3040;
  wire g30400;
  wire g30401;
  wire g30402;
  wire g30403;
  wire g30404;
  wire g30405;
  wire g30406;
  wire g30407;
  wire g30408;
  wire g30409;
  wire g30410;
  wire g30411;
  wire g30412;
  wire g30413;
  wire g30414;
  wire g30415;
  wire g30416;
  wire g30417;
  wire g30418;
  wire g30419;
  wire g30420;
  wire g30421;
  wire g30422;
  wire g30423;
  wire g30424;
  wire g30425;
  wire g30426;
  wire g30427;
  wire g30428;
  wire g30429;
  wire g30430;
  wire g30431;
  wire g30432;
  wire g30433;
  wire g30434;
  wire g30435;
  wire g30436;
  wire g30437;
  wire g30438;
  wire g30439;
  wire g30440;
  wire g30441;
  wire g30442;
  wire g30443;
  wire g30444;
  wire g30445;
  wire g30446;
  wire g30447;
  wire g30448;
  wire g30449;
  wire g3045;
  wire g30450;
  wire g30451;
  wire g30452;
  wire g30453;
  wire g30454;
  wire g30455;
  wire g30456;
  wire g30457;
  wire g30458;
  wire g30459;
  wire g30460;
  wire g30461;
  wire g30462;
  wire g30463;
  wire g30464;
  wire g30465;
  wire g30466;
  wire g30467;
  wire g30468;
  wire g30469;
  wire g30470;
  wire g30471;
  wire g30472;
  wire g30473;
  wire g30474;
  wire g30475;
  wire g30476;
  wire g30477;
  wire g30478;
  wire g30479;
  wire g30480;
  wire g30481;
  wire g30482;
  wire g30483;
  wire g30484;
  wire g30485;
  wire g30486;
  wire g30487;
  wire g30488;
  wire g30489;
  wire g30490;
  wire g30491;
  wire g30492;
  wire g30493;
  wire g30494;
  wire g30495;
  wire g30496;
  wire g30497;
  wire g30498;
  wire g30499;
  wire g305;
  wire g3050;
  wire g30500;
  wire g30501;
  wire g30502;
  wire g30503;
  wire g30504;
  wire g30505;
  wire g30506;
  wire g30507;
  wire g30508;
  wire g30509;
  wire g30510;
  wire g30511;
  wire g30512;
  wire g30513;
  wire g30514;
  wire g30515;
  wire g30516;
  wire g30517;
  wire g30518;
  wire g30519;
  wire g30520;
  wire g30521;
  wire g30522;
  wire g30523;
  wire g30524;
  wire g30525;
  wire g30526;
  wire g30527;
  wire g30528;
  wire g30529;
  wire g30530;
  wire g30531;
  wire g30532;
  wire g30533;
  wire g30534;
  wire g30535;
  wire g30536;
  wire g30537;
  wire g30538;
  wire g30539;
  wire g30540;
  wire g30541;
  wire g30542;
  wire g30543;
  wire g30544;
  wire g30545;
  wire g30546;
  wire g30547;
  wire g30548;
  wire g30549;
  wire g30550;
  wire g30551;
  wire g30552;
  wire g30553;
  wire g30554;
  wire g30555;
  wire g30556;
  wire g30557;
  wire g30558;
  wire g30559;
  wire g30560;
  wire g30561;
  wire g30562;
  wire g30563;
  wire g30565;
  wire g3057;
  wire g30591;
  wire g3061;
  wire g30610;
  wire g3065;
  wire g3068;
  wire g3072;
  wire g30729;
  wire g3080;
  wire g3085;
  wire g3089;
  wire g30917;
  wire g3092;
  wire g30928;
  wire g30931;
  wire g3096;
  wire g31;
  wire g3100;
  wire g3103;
  wire g3106;
  wire g311;
  wire g3111;
  wire g3115;
  wire g3119;
  wire g3125;
  wire g3129;
  wire g3133;
  wire g3139;
  wire g3143;
  wire g3147;
  wire g3151;
  output g31521;
  wire g31522;
  wire g3155;
  wire g31578;
  wire g316;
  wire g3161;
  wire g31655;
  output g31656;
  wire g31657;
  output g31665;
  wire g31666;
  wire g31667;
  wire g3167;
  wire g3171;
  wire g3179;
  wire g31791;
  output g31793;
  output g31860;
  output g31861;
  output g31862;
  output g31863;
  wire g31864;
  wire g31865;
  wire g31866;
  wire g31867;
  wire g31868;
  wire g31869;
  wire g3187;
  wire g31870;
  wire g31871;
  wire g31872;
  wire g31873;
  wire g31874;
  wire g31875;
  wire g31876;
  wire g31877;
  wire g31878;
  wire g31879;
  wire g31880;
  wire g31881;
  wire g31882;
  wire g31883;
  wire g31884;
  wire g31885;
  wire g31886;
  wire g31887;
  wire g31888;
  wire g31889;
  wire g31890;
  wire g31891;
  wire g31892;
  wire g31893;
  wire g31894;
  wire g31895;
  wire g31896;
  wire g31897;
  wire g31898;
  wire g31899;
  wire g319;
  wire g31900;
  wire g31901;
  wire g31902;
  wire g31903;
  wire g31904;
  wire g31905;
  wire g31906;
  wire g31907;
  wire g31908;
  wire g31909;
  wire g3191;
  wire g31910;
  wire g31911;
  wire g31912;
  wire g31913;
  wire g31914;
  wire g31915;
  wire g31916;
  wire g31917;
  wire g31918;
  wire g31919;
  wire g31920;
  wire g31921;
  wire g31922;
  wire g31923;
  wire g31924;
  wire g31925;
  wire g31926;
  wire g31927;
  wire g31928;
  wire g31929;
  wire g31930;
  wire g31931;
  wire g31932;
  wire g3195;
  wire g3199;
  wire g32021;
  wire g32024;
  wire g32027;
  wire g3203;
  wire g3207;
  wire g3211;
  wire g3215;
  output g32185;
  wire g32186;
  wire g3219;
  wire g3223;
  wire g3227;
  wire g3231;
  wire g3235;
  wire g32363;
  wire g32381;
  wire g3239;
  wire g324;
  wire g32407;
  output g32429;
  wire g3243;
  output g32454;
  wire g3247;
  wire g3251;
  wire g3255;
  wire g3259;
  wire g3263;
  wire g3267;
  wire g3274;
  wire g3281;
  wire g3288;
  wire g329;
  output g32975;
  wire g32976;
  wire g32977;
  wire g32978;
  wire g32979;
  wire g3298;
  wire g32980;
  wire g32981;
  wire g32982;
  wire g32983;
  wire g32984;
  wire g32985;
  wire g32986;
  wire g32987;
  wire g32988;
  wire g32989;
  wire g32990;
  wire g32991;
  wire g32992;
  wire g32993;
  wire g32994;
  wire g32995;
  wire g32996;
  wire g32997;
  wire g32998;
  wire g32999;
  wire g33000;
  wire g33001;
  wire g33002;
  wire g33003;
  wire g33004;
  wire g33005;
  wire g33006;
  wire g33007;
  wire g33008;
  wire g33009;
  wire g33010;
  wire g33011;
  wire g33012;
  wire g33013;
  wire g33014;
  wire g33015;
  wire g33016;
  wire g33017;
  wire g33018;
  wire g33019;
  wire g33020;
  wire g33021;
  wire g33022;
  wire g33023;
  wire g33024;
  wire g33025;
  wire g33026;
  wire g33027;
  wire g33028;
  wire g33029;
  wire g3303;
  wire g33030;
  wire g33031;
  wire g33032;
  wire g33033;
  wire g33034;
  wire g33035;
  wire g33036;
  wire g33037;
  wire g33038;
  wire g33039;
  wire g33040;
  wire g33041;
  wire g33042;
  wire g33043;
  wire g33044;
  wire g33045;
  wire g33046;
  wire g33047;
  wire g33048;
  wire g33049;
  wire g33050;
  wire g33051;
  wire g33052;
  wire g33053;
  wire g33054;
  wire g33055;
  wire g33056;
  wire g33057;
  wire g33058;
  wire g33059;
  wire g33060;
  wire g33061;
  wire g33062;
  wire g33063;
  wire g33064;
  wire g33065;
  wire g33066;
  wire g33067;
  wire g33068;
  wire g33069;
  wire g33070;
  wire g33076;
  output g33079;
  wire g33080;
  wire g3310;
  wire g33120;
  wire g33149;
  wire g33164;
  wire g3317;
  wire g33176;
  wire g33187;
  wire g33197;
  wire g33204;
  wire g3321;
  wire g33212;
  wire g33219;
  wire g33228;
  wire g3325;
  wire g33283;
  wire g3329;
  wire g333;
  wire g33318;
  wire g33323;
  wire g3333;
  wire g33354;
  wire g33377;
  wire g3338;
  wire g33388;
  wire g33391;
  wire g3343;
  output g33435;
  wire g33436;
  wire g3347;
  wire g3352;
  output g33533;
  wire g33534;
  wire g33535;
  wire g33536;
  wire g33537;
  wire g33538;
  wire g33539;
  wire g33540;
  wire g33541;
  wire g33542;
  wire g33543;
  wire g33544;
  wire g33545;
  wire g33546;
  wire g33547;
  wire g33548;
  wire g33549;
  wire g3355;
  wire g33550;
  wire g33551;
  wire g33552;
  wire g33553;
  wire g33554;
  wire g33555;
  wire g33556;
  wire g33557;
  wire g33558;
  wire g33559;
  wire g33560;
  wire g33561;
  wire g33562;
  wire g33563;
  wire g33564;
  wire g33565;
  wire g33566;
  wire g33567;
  wire g33568;
  wire g33569;
  wire g33570;
  wire g33571;
  wire g33572;
  wire g33573;
  wire g33574;
  wire g33575;
  wire g33576;
  wire g33577;
  wire g33578;
  wire g33579;
  wire g33580;
  wire g33581;
  wire g33582;
  wire g33583;
  wire g33584;
  wire g33585;
  wire g33586;
  wire g33587;
  wire g33588;
  wire g33589;
  wire g33590;
  wire g33591;
  wire g33592;
  wire g33593;
  wire g33594;
  wire g33595;
  wire g33596;
  wire g33597;
  wire g33598;
  wire g33599;
  wire g336;
  wire g33600;
  wire g33601;
  wire g33602;
  wire g33603;
  wire g33604;
  wire g33605;
  wire g33606;
  wire g33607;
  wire g33608;
  wire g33609;
  wire g3361;
  wire g33610;
  wire g33611;
  wire g33612;
  wire g33613;
  wire g33614;
  wire g33615;
  wire g33616;
  wire g33617;
  wire g33618;
  wire g33619;
  wire g33620;
  wire g33621;
  wire g33622;
  wire g33623;
  wire g33624;
  wire g33625;
  wire g33626;
  wire g33627;
  wire g33628;
  wire g33631;
  output g33636;
  wire g33637;
  wire g33638;
  wire g33641;
  wire g33645;
  wire g33648;
  wire g33653;
  output g33659;
  wire g33660;
  wire g33661;
  wire g33665;
  wire g33670;
  wire g3368;
  wire g33682;
  wire g33688;
  wire g33691;
  wire g33696;
  wire g33698;
  wire g33702;
  wire g33705;
  wire g33708;
  wire g33712;
  wire g33713;
  wire g33716;
  wire g3372;
  wire g33726;
  wire g33729;
  wire g33736;
  wire g33744;
  wire g33750;
  wire g33755;
  wire g3376;
  wire g33761;
  wire g33766;
  wire g33772;
  wire g33778;
  wire g33791;
  wire g3380;
  wire g33800;
  wire g33804;
  wire g33806;
  wire g33813;
  wire g33827;
  wire g33839;
  wire g33845;
  wire g3385;
  wire g33850;
  output g33874;
  wire g33875;
  output g33894;
  wire g33895;
  wire g3391;
  wire g33912;
  wire g33916;
  wire g33917;
  wire g33918;
  wire g33920;
  wire g33923;
  wire g33926;
  wire g33928;
  wire g33929;
  wire g33931;
  wire g33932;
  wire g33934;
  output g33935;
  wire g33936;
  wire g33937;
  output g33945;
  output g33946;
  output g33947;
  output g33948;
  output g33949;
  output g33950;
  output g33959;
  wire g3396;
  wire g33960;
  wire g33961;
  wire g33962;
  wire g33963;
  wire g33964;
  wire g33965;
  wire g33966;
  wire g33967;
  wire g33968;
  wire g33969;
  wire g33970;
  wire g33971;
  wire g33972;
  wire g33973;
  wire g33974;
  wire g33975;
  wire g33976;
  wire g33977;
  wire g33978;
  wire g33979;
  wire g33980;
  wire g33981;
  wire g33982;
  wire g33983;
  wire g33984;
  wire g33985;
  wire g33986;
  wire g33987;
  wire g33988;
  wire g33989;
  wire g33990;
  wire g33991;
  wire g33992;
  wire g33993;
  wire g33994;
  wire g33995;
  wire g33996;
  wire g33997;
  wire g33998;
  wire g33999;
  wire g34;
  wire g34000;
  wire g34001;
  wire g34002;
  wire g34003;
  wire g34004;
  wire g34005;
  wire g34006;
  wire g34007;
  wire g34008;
  wire g34009;
  wire g3401;
  wire g34010;
  wire g34011;
  wire g34012;
  wire g34013;
  wire g34014;
  wire g34015;
  wire g34016;
  wire g34017;
  wire g34018;
  wire g34019;
  wire g34020;
  wire g34021;
  wire g34022;
  wire g34023;
  wire g34024;
  wire g34025;
  wire g34026;
  wire g34027;
  wire g34028;
  wire g34029;
  wire g34030;
  wire g34031;
  wire g34032;
  wire g34033;
  wire g34034;
  wire g34035;
  wire g34036;
  wire g34037;
  wire g34038;
  wire g34039;
  wire g34040;
  wire g34041;
  wire g34052;
  wire g34059;
  wire g3408;
  wire g341;
  wire g34118;
  wire g3412;
  wire g34121;
  wire g34122;
  wire g34123;
  wire g34126;
  wire g34127;
  wire g34130;
  wire g34131;
  wire g34134;
  wire g34142;
  wire g34144;
  wire g34145;
  wire g34150;
  wire g34151;
  wire g34152;
  wire g34153;
  wire g34159;
  wire g3416;
  wire g34160;
  wire g3419;
  wire g34195;
  output g34201;
  wire g34202;
  wire g34208;
  wire g34209;
  wire g34210;
  output g34221;
  wire g34222;
  wire g3423;
  output g34232;
  output g34233;
  output g34234;
  output g34235;
  output g34236;
  output g34237;
  output g34238;
  output g34239;
  output g34240;
  wire g34241;
  wire g34242;
  wire g34243;
  wire g34244;
  wire g34245;
  wire g34246;
  wire g34247;
  wire g34248;
  wire g34249;
  wire g34250;
  wire g34251;
  wire g34252;
  wire g34253;
  wire g34254;
  wire g34255;
  wire g34256;
  wire g34257;
  wire g34258;
  wire g34259;
  wire g34260;
  wire g34261;
  wire g34262;
  wire g34263;
  wire g34264;
  wire g34265;
  wire g34266;
  wire g34267;
  wire g34268;
  wire g34269;
  wire g34272;
  wire g34273;
  wire g34274;
  wire g34275;
  wire g34276;
  wire g34277;
  wire g34278;
  wire g34280;
  wire g34282;
  wire g34283;
  wire g34285;
  wire g34286;
  wire g34288;
  wire g34289;
  wire g34290;
  wire g34292;
  wire g34293;
  wire g34294;
  wire g34296;
  wire g34297;
  wire g34300;
  wire g34302;
  wire g34303;
  wire g34304;
  wire g34305;
  wire g34306;
  wire g3431;
  wire g34314;
  wire g34318;
  wire g34321;
  wire g34331;
  wire g34347;
  wire g34349;
  wire g34350;
  wire g34352;
  wire g34353;
  wire g34358;
  wire g3436;
  wire g34366;
  wire g34368;
  wire g34369;
  wire g34372;
  wire g34373;
  wire g34374;
  wire g34376;
  wire g34377;
  wire g34379;
  output g34383;
  wire g34384;
  wire g34387;
  wire g34391;
  wire g34399;
  wire g344;
  wire g3440;
  wire g34402;
  wire g34403;
  wire g34404;
  wire g34405;
  wire g34406;
  wire g34407;
  wire g34411;
  wire g34412;
  wire g34416;
  wire g34417;
  wire g34421;
  output g34425;
  wire g34426;
  wire g34427;
  wire g34428;
  wire g34429;
  wire g3443;
  wire g34430;
  wire g34431;
  wire g34432;
  wire g34433;
  wire g34434;
  output g34435;
  output g34436;
  output g34437;
  wire g34438;
  wire g34439;
  wire g34440;
  wire g34441;
  wire g34442;
  wire g34443;
  wire g34444;
  wire g34445;
  wire g34446;
  wire g34447;
  wire g34448;
  wire g34449;
  wire g34450;
  wire g34451;
  wire g34452;
  wire g34453;
  wire g34454;
  wire g34455;
  wire g34456;
  wire g34457;
  wire g34458;
  wire g34459;
  wire g34460;
  wire g34461;
  wire g34462;
  wire g34463;
  wire g34464;
  wire g34465;
  wire g34466;
  wire g34467;
  wire g34468;
  wire g3447;
  wire g34471;
  wire g34472;
  wire g34480;
  wire g34494;
  wire g34501;
  wire g34504;
  wire g34505;
  wire g3451;
  wire g34510;
  wire g34511;
  wire g34512;
  wire g34521;
  wire g34522;
  wire g3454;
  wire g34540;
  wire g3457;
  wire g34570;
  wire g34579;
  wire g34589;
  wire g34590;
  wire g34591;
  wire g34592;
  wire g34593;
  wire g34594;
  wire g34595;
  wire g34596;
  output g34597;
  wire g34598;
  wire g34599;
  wire g34600;
  wire g34601;
  wire g34602;
  wire g34603;
  wire g34604;
  wire g34605;
  wire g34606;
  wire g34607;
  wire g34608;
  wire g34609;
  wire g34610;
  wire g34611;
  wire g34612;
  wire g34613;
  wire g34614;
  wire g34615;
  wire g34616;
  wire g34617;
  wire g34618;
  wire g34619;
  wire g3462;
  wire g34620;
  wire g34621;
  wire g34622;
  wire g34623;
  wire g34624;
  wire g34625;
  wire g34626;
  wire g34627;
  wire g34628;
  wire g34629;
  wire g34630;
  wire g34631;
  wire g34632;
  wire g34633;
  wire g34634;
  wire g34635;
  wire g34636;
  wire g34637;
  wire g34638;
  wire g34639;
  wire g34640;
  wire g34641;
  wire g34642;
  wire g34643;
  wire g34644;
  wire g34645;
  wire g34646;
  wire g34647;
  wire g34648;
  wire g34649;
  wire g34650;
  wire g34653;
  wire g34654;
  wire g34656;
  wire g34657;
  wire g34659;
  wire g3466;
  wire g34660;
  wire g34663;
  wire g34688;
  wire g34690;
  wire g34699;
  wire g347;
  wire g3470;
  wire g34708;
  wire g34711;
  wire g34712;
  wire g34713;
  wire g34714;
  wire g34716;
  wire g34717;
  wire g34718;
  wire g34719;
  wire g34720;
  wire g34721;
  wire g34722;
  wire g34723;
  wire g34724;
  wire g34725;
  wire g34726;
  wire g34727;
  wire g34728;
  wire g34729;
  wire g34730;
  wire g34731;
  wire g34732;
  wire g34733;
  wire g34734;
  wire g34735;
  wire g34736;
  wire g34739;
  wire g34749;
  wire g34755;
  wire g34759;
  wire g3476;
  wire g34760;
  wire g34767;
  wire g34768;
  wire g34769;
  wire g34770;
  wire g34772;
  wire g34773;
  wire g34775;
  wire g34776;
  wire g34777;
  wire g34778;
  wire g34781;
  wire g34783;
  wire g34784;
  wire g34785;
  wire g34786;
  wire g34787;
  output g34788;
  wire g34789;
  wire g34790;
  wire g34791;
  wire g34792;
  wire g34793;
  wire g34794;
  wire g34795;
  wire g34796;
  wire g34797;
  wire g34798;
  wire g34799;
  wire g3480;
  wire g34800;
  wire g34801;
  wire g34802;
  wire g34803;
  wire g34804;
  wire g34805;
  wire g34806;
  wire g34807;
  wire g34808;
  wire g34809;
  wire g34810;
  wire g34812;
  wire g34813;
  wire g34816;
  wire g34820;
  wire g34823;
  wire g34827;
  wire g34830;
  wire g34833;
  wire g34836;
  output g34839;
  wire g3484;
  wire g34840;
  wire g34843;
  wire g34846;
  wire g34847;
  wire g34848;
  wire g34849;
  wire g34850;
  wire g34851;
  wire g34852;
  wire g34855;
  wire g34877;
  wire g34878;
  wire g34879;
  wire g34880;
  wire g34881;
  wire g34882;
  wire g34884;
  wire g34887;
  wire g34890;
  wire g34893;
  wire g34894;
  wire g34897;
  wire g3490;
  wire g34900;
  wire g34903;
  wire g34906;
  wire g34910;
  wire g34911;
  output g34913;
  wire g34914;
  output g34915;
  wire g34916;
  output g34917;
  wire g34918;
  output g34919;
  wire g34920;
  output g34921;
  wire g34922;
  output g34923;
  wire g34924;
  output g34925;
  wire g34926;
  output g34927;
  wire g34928;
  wire g34929;
  wire g34930;
  wire g34935;
  wire g3494;
  wire g34943;
  wire g34944;
  wire g34945;
  wire g34946;
  wire g34947;
  wire g34949;
  wire g34950;
  wire g34951;
  wire g34952;
  wire g34954;
  output g34956;
  wire g34957;
  wire g34970;
  wire g34971;
  output g34972;
  wire g34973;
  wire g34974;
  wire g34975;
  wire g34976;
  wire g34977;
  wire g34978;
  wire g34979;
  wire g3498;
  wire g34980;
  wire g34982;
  wire g34983;
  wire g34984;
  wire g34985;
  wire g34986;
  wire g34987;
  wire g34988;
  wire g34989;
  wire g34990;
  wire g34991;
  wire g34992;
  wire g34993;
  wire g34994;
  wire g34995;
  wire g34996;
  wire g34997;
  wire g34998;
  input g35;
  wire g35000;
  wire g35001;
  wire g35002;
  wire g3502;
  wire g3506;
  wire g351;
  wire g3512;
  wire g3518;
  wire g3522;
  wire g3530;
  wire g3538;
  wire g3542;
  wire g3546;
  wire g355;
  wire g3550;
  wire g3554;
  wire g3558;
  wire g3562;
  wire g3566;
  wire g3570;
  wire g3574;
  wire g3578;
  wire g358;
  wire g3582;
  wire g3586;
  wire g3590;
  wire g3594;
  wire g3598;
  input g36;
  wire g3602;
  wire g3606;
  wire g3610;
  wire g3614;
  wire g3618;
  wire g3625;
  wire g3632;
  wire g3639;
  wire g3649;
  wire g365;
  wire g3654;
  wire g3661;
  wire g3668;
  wire g3672;
  wire g3676;
  wire g3680;
  wire g3684;
  wire g3689;
  wire g3694;
  wire g3698;
  wire g37;
  wire g370;
  wire g3703;
  wire g3706;
  wire g3712;
  wire g3719;
  wire g3723;
  wire g3727;
  wire g3731;
  wire g3736;
  wire g3742;
  wire g3747;
  wire g3752;
  wire g3759;
  wire g376;
  wire g3763;
  wire g3767;
  wire g3770;
  wire g3774;
  wire g3782;
  wire g3787;
  wire g3791;
  wire g3794;
  wire g3798;
  wire g3802;
  wire g3805;
  wire g3808;
  wire g3813;
  wire g3817;
  wire g3821;
  wire g3827;
  wire g3831;
  wire g3835;
  wire g3841;
  wire g3845;
  wire g3849;
  wire g385;
  wire g3853;
  wire g3857;
  wire g3863;
  wire g3869;
  wire g3873;
  wire g3881;
  wire g3889;
  wire g3893;
  wire g3897;
  wire g3901;
  wire g3905;
  wire g3909;
  wire g391;
  wire g3913;
  wire g3917;
  wire g392;
  wire g3921;
  wire g3925;
  wire g3929;
  wire g3933;
  wire g3937;
  wire g3941;
  wire g3945;
  wire g3949;
  wire g3953;
  wire g3957;
  wire g3961;
  wire g3965;
  wire g3969;
  wire g3976;
  wire g3983;
  wire g3990;
  wire g4000;
  wire g4005;
  wire g401;
  wire g4012;
  wire g4019;
  wire g4023;
  wire g4027;
  wire g4031;
  wire g4035;
  wire g4040;
  wire g4045;
  wire g4049;
  wire g405;
  wire g4054;
  wire g4057;
  wire g4064;
  wire g4072;
  wire g4076;
  wire g4082;
  wire g4087;
  wire g4093;
  wire g4098;
  wire g4104;
  wire g4108;
  wire g411;
  wire g4112;
  wire g4116;
  wire g4119;
  wire g4122;
  wire g4125;
  wire g4129;
  wire g4132;
  wire g4135;
  wire g4138;
  wire g4141;
  wire g4145;
  wire g4146;
  wire g4153;
  wire g4157;
  wire g4164;
  wire g4165;
  wire g4169;
  wire g417;
  wire g4172;
  wire g4176;
  wire g4180;
  wire g4185;
  wire g4188;
  wire g4191;
  wire g4194;
  wire g4197;
  wire g4200;
  wire g4204;
  wire g4207;
  wire g4210;
  wire g4213;
  wire g4216;
  wire g4219;
  wire g4222;
  wire g4226;
  wire g4229;
  wire g4232;
  wire g4235;
  wire g4239;
  wire g424;
  wire g4242;
  wire g4245;
  wire g4249;
  wire g4253;
  wire g4258;
  wire g4264;
  wire g4269;
  wire g4273;
  wire g4277;
  wire g4281;
  wire g4284;
  wire g4287;
  wire g429;
  wire g4291;
  wire g4294;
  wire g4297;
  wire g43;
  wire g4300;
  wire g4304;
  wire g4308;
  wire g4311;
  wire g4322;
  wire g433;
  wire g4332;
  wire g4340;
  wire g4349;
  wire g4358;
  wire g4366;
  wire g4369;
  wire g437;
  wire g4372;
  wire g4375;
  wire g4382;
  wire g4388;
  wire g4392;
  input g44;
  wire g4401;
  wire g4405;
  wire g4408;
  wire g441;
  wire g4411;
  wire g4414;
  wire g4417;
  wire g4420;
  wire g4423;
  wire g4427;
  wire g4430;
  wire g4434;
  wire g4438;
  wire g4443;
  wire g4446;
  wire g4449;
  wire g4452;
  wire g4455;
  wire g4456;
  wire g4459;
  wire g446;
  wire g4462;
  wire g4467;
  wire g4473;
  wire g4474;
  wire g4477;
  wire g4480;
  wire g4483;
  wire g4486;
  wire g4489;
  wire g4492;
  wire g4495;
  wire g4498;
  wire g45;
  wire g4501;
  wire g4504;
  wire g4507;
  wire g4512;
  wire g4515;
  wire g4519;
  wire g452;
  wire g4520;
  wire g4521;
  wire g4527;
  wire g4531;
  wire g4534;
  wire g4537;
  wire g4540;
  wire g4543;
  wire g4546;
  wire g4549;
  wire g4552;
  wire g4555;
  wire g4558;
  wire g4561;
  wire g4564;
  wire g4567;
  wire g457;
  wire g4570;
  wire g4571;
  wire g4572;
  wire g4575;
  wire g4578;
  wire g4581;
  wire g4584;
  wire g4593;
  wire g46;
  wire g460;
  wire g4601;
  wire g4608;
  wire g4616;
  wire g4621;
  wire g4628;
  wire g4633;
  wire g4639;
  wire g464;
  wire g4643;
  wire g4646;
  wire g4653;
  wire g4659;
  wire g4664;
  wire g4669;
  wire g4674;
  wire g468;
  wire g4681;
  wire g4688;
  wire g4698;
  wire g47;
  wire g4704;
  wire g4709;
  wire g471;
  wire g4717;
  wire g4722;
  wire g4727;
  wire g4732;
  wire g4737;
  wire g4741;
  wire g4742;
  wire g4743;
  wire g4749;
  wire g475;
  wire g4754;
  wire g4760;
  wire g4765;
  wire g4771;
  wire g4776;
  wire g4785;
  wire g479;
  wire g4793;
  wire g48;
  wire g4801;
  wire g4809;
  wire g4812;
  wire g4815;
  wire g4818;
  wire g482;
  wire g4821;
  wire g4826;
  wire g4831;
  wire g4836;
  wire g4843;
  wire g4849;
  wire g4854;
  wire g4859;
  wire g4864;
  wire g4871;
  wire g4878;
  wire g4888;
  wire g4894;
  wire g4899;
  wire g49;
  wire g490;
  wire g4907;
  wire g4912;
  wire g4917;
  wire g4922;
  wire g4927;
  wire g4931;
  wire g4932;
  wire g4933;
  wire g4939;
  wire g4944;
  wire g4950;
  wire g4955;
  wire g496;
  wire g4961;
  wire g4966;
  wire g4975;
  wire g4983;
  wire g499;
  wire g4991;
  wire g4999;
  input g5;
  wire g50;
  wire g5002;
  wire g5005;
  wire g5008;
  wire g5011;
  wire g5016;
  wire g5022;
  wire g5029;
  wire g5033;
  wire g5037;
  wire g504;
  wire g5041;
  wire g5046;
  wire g5052;
  wire g5057;
  wire g5062;
  wire g5069;
  wire g5073;
  wire g5077;
  wire g5080;
  wire g5084;
  wire g5092;
  wire g5097;
  wire g51;
  wire g5101;
  wire g5105;
  wire g5109;
  wire g5112;
  wire g5115;
  wire g5120;
  wire g5124;
  wire g5128;
  wire g513;
  wire g5134;
  wire g5138;
  wire g5142;
  wire g5148;
  wire g5152;
  wire g5156;
  wire g5160;
  wire g5164;
  wire g5170;
  wire g5176;
  wire g518;
  wire g5180;
  wire g5188;
  wire g5196;
  wire g52;
  wire g5200;
  wire g5204;
  wire g5208;
  wire g5212;
  wire g5216;
  wire g5220;
  wire g5224;
  wire g5228;
  wire g5232;
  wire g5236;
  wire g5240;
  wire g5244;
  wire g5248;
  wire g5252;
  wire g5256;
  wire g5260;
  wire g5264;
  wire g5268;
  wire g5272;
  wire g5276;
  wire g528;
  wire g5283;
  wire g5290;
  wire g5297;
  input g53;
  wire g5308;
  wire g5313;
  wire g5320;
  wire g5327;
  wire g5331;
  wire g5335;
  wire g5339;
  wire g534;
  wire g5343;
  wire g5348;
  wire g5352;
  wire g5357;
  wire g5360;
  wire g5366;
  wire g5373;
  wire g5377;
  wire g538;
  wire g5381;
  wire g5385;
  wire g5390;
  wire g5396;
  input g54;
  wire g5401;
  wire g5406;
  wire g5413;
  wire g5417;
  wire g542;
  wire g5421;
  wire g5424;
  wire g5428;
  wire g5436;
  wire g5441;
  wire g5445;
  wire g5448;
  wire g5452;
  wire g5456;
  wire g5459;
  wire g546;
  wire g5462;
  wire g5467;
  wire g5471;
  wire g5475;
  wire g5481;
  wire g5485;
  wire g5489;
  wire g5495;
  wire g5499;
  wire g55;
  wire g550;
  wire g5503;
  wire g5507;
  wire g5511;
  wire g5517;
  wire g5523;
  wire g5527;
  wire g5535;
  wire g554;
  wire g5543;
  wire g5547;
  wire g5551;
  wire g5555;
  wire g5559;
  wire g5563;
  wire g5567;
  wire g5571;
  wire g5575;
  wire g5579;
  wire g5583;
  wire g5587;
  wire g559;
  wire g5591;
  wire g5595;
  wire g5599;
  input g56;
  wire g5603;
  wire g5607;
  wire g5611;
  wire g5615;
  wire g5619;
  wire g562;
  wire g5623;
  wire g5630;
  wire g5637;
  wire g5644;
  wire g5654;
  wire g5659;
  wire g5666;
  wire g5673;
  wire g5677;
  wire g568;
  wire g5681;
  wire g5685;
  wire g5689;
  wire g5694;
  wire g5698;
  input g57;
  wire g5703;
  wire g5706;
  wire g5712;
  wire g5719;
  wire g572;
  wire g5723;
  wire g5727;
  wire g5731;
  wire g5736;
  wire g5742;
  wire g5747;
  wire g5752;
  wire g5759;
  wire g5763;
  wire g5767;
  wire g577;
  wire g5770;
  wire g5774;
  wire g5782;
  wire g5787;
  wire g5791;
  wire g5794;
  wire g5798;
  wire g5802;
  wire g5805;
  wire g5808;
  wire g5813;
  wire g5817;
  wire g582;
  wire g5821;
  wire g5827;
  wire g5831;
  wire g5835;
  wire g5841;
  wire g5845;
  wire g5849;
  wire g5853;
  wire g5857;
  wire g586;
  wire g5863;
  wire g5869;
  wire g5873;
  wire g5881;
  wire g5889;
  wire g5893;
  wire g5897;
  wire g59;
  wire g590;
  wire g5901;
  wire g5905;
  wire g5909;
  wire g5913;
  wire g5917;
  wire g5921;
  wire g5925;
  wire g5929;
  wire g5933;
  wire g5937;
  wire g5941;
  wire g5945;
  wire g5949;
  wire g595;
  wire g5953;
  wire g5957;
  wire g5961;
  wire g5965;
  wire g5969;
  wire g5976;
  wire g5983;
  wire g599;
  wire g5990;
  wire g6;
  wire g6000;
  wire g6005;
  wire g6012;
  wire g6019;
  wire g6023;
  wire g6027;
  wire g6031;
  wire g6035;
  wire g604;
  wire g6040;
  wire g6044;
  wire g6049;
  wire g6052;
  wire g6058;
  wire g6065;
  wire g6069;
  wire g6073;
  wire g6077;
  wire g608;
  wire g6082;
  wire g6088;
  wire g6093;
  wire g6098;
  wire g6105;
  wire g6109;
  wire g6113;
  wire g6116;
  wire g6120;
  wire g6128;
  wire g613;
  wire g6133;
  wire g6137;
  wire g6140;
  wire g6144;
  wire g6148;
  wire g6151;
  wire g6154;
  wire g6159;
  wire g6163;
  wire g6167;
  wire g617;
  wire g6173;
  wire g6177;
  wire g6181;
  wire g6187;
  wire g6191;
  wire g6195;
  wire g6199;
  wire g6203;
  wire g6209;
  wire g6215;
  wire g6219;
  wire g622;
  wire g6227;
  wire g6235;
  wire g6239;
  wire g6243;
  wire g6247;
  wire g6251;
  wire g6255;
  wire g6259;
  wire g626;
  wire g6263;
  wire g6267;
  wire g6271;
  wire g6275;
  wire g6279;
  wire g6283;
  wire g6287;
  wire g6291;
  wire g6295;
  wire g6299;
  wire g63;
  wire g6303;
  wire g6307;
  wire g6311;
  wire g6315;
  wire g632;
  wire g6322;
  wire g6329;
  wire g6336;
  wire g6346;
  wire g6351;
  wire g6358;
  wire g6365;
  wire g6369;
  wire g637;
  wire g6373;
  wire g6377;
  wire g6381;
  wire g6386;
  wire g6390;
  wire g6395;
  wire g6398;
  input g64;
  wire g640;
  wire g6404;
  wire g6411;
  wire g6415;
  wire g6419;
  wire g6423;
  wire g6428;
  wire g6434;
  wire g6439;
  wire g6444;
  wire g645;
  wire g6451;
  wire g6455;
  wire g6459;
  wire g6462;
  wire g6466;
  wire g6474;
  wire g6479;
  wire g6483;
  wire g6486;
  wire g6490;
  wire g6494;
  wire g6497;
  wire g65;
  wire g650;
  wire g6500;
  wire g6505;
  wire g6509;
  wire g6513;
  wire g6519;
  wire g6523;
  wire g6527;
  wire g6533;
  wire g6537;
  wire g6541;
  wire g6545;
  wire g6549;
  wire g655;
  wire g6555;
  wire g6561;
  wire g6565;
  wire g6573;
  wire g6581;
  wire g6585;
  wire g6589;
  wire g6593;
  wire g6597;
  wire g66;
  wire g6601;
  wire g6605;
  wire g6609;
  wire g661;
  wire g6613;
  wire g6617;
  wire g6621;
  wire g6625;
  wire g6629;
  wire g6633;
  wire g6637;
  wire g6641;
  wire g6645;
  wire g6649;
  wire g6653;
  wire g6657;
  wire g6661;
  wire g6668;
  wire g667;
  wire g6675;
  wire g6682;
  wire g6692;
  wire g6697;
  wire g6704;
  wire g671;
  wire g6711;
  wire g6715;
  wire g6719;
  wire g6723;
  wire g6727;
  wire g6732;
  wire g6736;
  wire g6741;
  input g6744;
  input g6745;
  input g6746;
  input g6747;
  input g6748;
  input g6749;
  input g6750;
  input g6751;
  input g6752;
  input g6753;
  wire g6754;
  wire g6755;
  wire g6756;
  wire g676;
  wire g6767;
  wire g6772;
  wire g6782;
  wire g6789;
  wire g681;
  wire g6821;
  wire g6832;
  wire g6856;
  wire g686;
  wire g6867;
  wire g6868;
  wire g6869;
  wire g6875;
  wire g6888;
  wire g6905;
  wire g691;
  wire g6928;
  wire g6946;
  wire g6955;
  wire g6961;
  wire g6971;
  wire g6972;
  wire g6973;
  wire g6974;
  wire g6976;
  wire g6977;
  wire g699;
  wire g7;
  wire g70;
  wire g7004;
  wire g7028;
  wire g703;
  wire g7051;
  wire g7074;
  wire g7097;
  wire g71;
  wire g7117;
  wire g7121;
  wire g714;
  wire g7148;
  wire g7161;
  wire g718;
  wire g7196;
  input g72;
  wire g723;
  wire g7231;
  output g7243;
  output g7245;
  output g7257;
  output g7260;
  wire g728;
  input g73;
  wire g732;
  wire g736;
  wire g739;
  wire g74;
  wire g744;
  wire g7474;
  wire g749;
  wire g7502;
  wire g7515;
  wire g7516;
  wire g7526;
  wire g7527;
  wire g753;
  output g7540;
  wire g7542;
  wire g7543;
  wire g7558;
  wire g7565;
  wire g7566;
  wire g758;
  wire g7586;
  wire g7593;
  wire g7594;
  wire g7595;
  wire g7596;
  wire g7615;
  wire g7616;
  wire g7617;
  wire g7618;
  wire g7623;
  wire g7624;
  wire g7625;
  wire g7626;
  wire g763;
  wire g7632;
  wire g7633;
  wire g7634;
  wire g7640;
  wire g7647;
  wire g7648;
  wire g7659;
  wire g7660;
  wire g767;
  wire g7674;
  wire g7689;
  wire g7704;
  wire g7717;
  wire g772;
  wire g7738;
  wire g7753;
  wire g776;
  wire g7766;
  wire g7791;
  wire g781;
  wire g7812;
  wire g7831;
  wire g785;
  wire g79;
  wire g790;
  output g7916;
  wire g794;
  output g7946;
  wire g799;
  wire g7993;
  wire g7994;
  wire g8;
  wire g802;
  wire g8032;
  wire g8038;
  wire g807;
  wire g8085;
  wire g812;
  output g8132;
  wire g8134;
  wire g8135;
  wire g817;
  output g8178;
  output g8215;
  wire g822;
  output g8235;
  wire g827;
  output g8277;
  output g8279;
  output g8283;
  wire g8285;
  output g8291;
  wire g832;
  output g8342;
  output g8344;
  output g8353;
  wire g8355;
  output g8358;
  wire g837;
  output g8398;
  input g84;
  output g8403;
  wire g8405;
  wire g8411;
  output g8416;
  wire g843;
  wire g847;
  wire g8470;
  output g8475;
  wire g8481;
  wire g85;
  wire g8515;
  wire g854;
  wire g8542;
  wire g8572;
  wire g859;
  wire g8595;
  wire g86;
  wire g8607;
  wire g862;
  wire g869;
  wire g8703;
  wire g8712;
  output g8719;
  wire g872;
  wire g8740;
  wire g875;
  wire g8757;
  wire g8763;
  wire g8778;
  wire g878;
  output g8783;
  output g8784;
  output g8785;
  output g8786;
  output g8787;
  output g8788;
  output g8789;
  wire g8791;
  wire g8792;
  wire g8795;
  wire g8805;
  wire g881;
  wire g8812;
  wire g8818;
  wire g8821;
  output g8839;
  wire g884;
  wire g8841;
  wire g8844;
  wire g887;
  output g8870;
  wire g8876;
  wire g8879;
  wire g8880;
  wire g890;
  output g8915;
  output g8916;
  output g8917;
  output g8918;
  output g8919;
  output g8920;
  wire g8922;
  wire g8925;
  wire g896;
  wire g8971;
  wire g8974;
  wire g8989;
  wire g9;
  input g90;
  wire g901;
  output g9019;
  wire g9021;
  wire g904;
  output g9048;
  wire g907;
  wire g9071;
  input g91;
  wire g911;
  wire g914;
  wire g9152;
  wire g9153;
  wire g9154;
  wire g9155;
  wire g918;
  wire g9185;
  wire g9186;
  input g92;
  wire g921;
  wire g9213;
  wire g9245;
  wire g925;
  output g9251;
  wire g9280;
  wire g9281;
  wire g929;
  wire g93;
  wire g930;
  wire g933;
  wire g9340;
  wire g936;
  wire g939;
  wire g94;
  wire g9417;
  wire g943;
  wire g947;
  wire g9477;
  wire g9478;
  output g9497;
  wire g952;
  output g9553;
  output g9555;
  wire g956;
  output g9615;
  output g9617;
  wire g962;
  wire g9637;
  wire g967;
  wire g968;
  output g9680;
  output g9682;
  wire g9687;
  wire g969;
  output g9741;
  output g9743;
  wire g9746;
  wire g9747;
  wire g976;
  wire g9772;
  wire g9780;
  wire g979;
  output g9817;
  wire g9864;
  input g99;
  wire g990;
  wire g9917;
  wire g9935;
  wire g996;
  al_oa21ftt _04563_ (
    .a(\DFF_746.Q ),
    .b(\DFF_233.Q ),
    .c(\DFF_845.Q ),
    .y(_00000_)
  );
  al_oai21 _04564_ (
    .a(\DFF_302.Q ),
    .b(\DFF_746.Q ),
    .c(_00000_),
    .y(_00001_)
  );
  al_nand3fft _04565_ (
    .a(\DFF_845.Q ),
    .b(\DFF_746.Q ),
    .c(\DFF_1112.Q ),
    .y(_00002_)
  );
  al_nand3ftt _04566_ (
    .a(\DFF_845.Q ),
    .b(\DFF_284.Q ),
    .c(\DFF_746.Q ),
    .y(_00003_)
  );
  al_and3 _04567_ (
    .a(_00002_),
    .b(_00003_),
    .c(_00001_),
    .y(\DFF_1220.D )
  );
  al_inv _04568_ (
    .a(\DFF_576.Q ),
    .y(g23652)
  );
  al_and3 _04569_ (
    .a(\DFF_598.Q ),
    .b(\DFF_68.Q ),
    .c(\DFF_1098.Q ),
    .y(g26801)
  );
  al_nand2 _04570_ (
    .a(g113),
    .b(\DFF_1035.Q ),
    .y(g31665)
  );
  al_and3fft _04571_ (
    .a(\DFF_1074.Q ),
    .b(g57),
    .c(g54),
    .y(_00004_)
  );
  al_nand3fft _04572_ (
    .a(g56),
    .b(g53),
    .c(_00004_),
    .y(_00005_)
  );
  al_inv _04573_ (
    .a(_00005_),
    .y(\DFF_748.D )
  );
  al_inv _04574_ (
    .a(\DFF_865.Q ),
    .y(g23759)
  );
  al_inv _04575_ (
    .a(\DFF_748.Q ),
    .y(g23190)
  );
  al_inv _04576_ (
    .a(g5),
    .y(g12833)
  );
  al_and3fft _04577_ (
    .a(\DFF_894.Q ),
    .b(\DFF_849.Q ),
    .c(\DFF_1311.Q ),
    .y(_00006_)
  );
  al_and3fft _04578_ (
    .a(\DFF_412.Q ),
    .b(\DFF_452.Q ),
    .c(\DFF_62.Q ),
    .y(_00007_)
  );
  al_nand3 _04579_ (
    .a(\DFF_270.Q ),
    .b(\DFF_604.Q ),
    .c(\DFF_1373.Q ),
    .y(_00008_)
  );
  al_nand3ftt _04580_ (
    .a(_00008_),
    .b(_00006_),
    .c(_00007_),
    .y(_00009_)
  );
  al_and2 _04581_ (
    .a(\DFF_792.Q ),
    .b(_00009_),
    .y(g28753)
  );
  al_nand2 _04582_ (
    .a(\DFF_1289.Q ),
    .b(\DFF_852.Q ),
    .y(_00010_)
  );
  al_aoi21ttf _04583_ (
    .a(\DFF_1336.Q ),
    .b(\DFF_899.Q ),
    .c(_00010_),
    .y(_00011_)
  );
  al_aoi21ttf _04584_ (
    .a(\DFF_155.Q ),
    .b(\DFF_1282.Q ),
    .c(_00011_),
    .y(_00012_)
  );
  al_nand2 _04585_ (
    .a(\DFF_15.Q ),
    .b(\DFF_531.Q ),
    .y(_00013_)
  );
  al_aoi21ttf _04586_ (
    .a(\DFF_95.Q ),
    .b(\DFF_1151.Q ),
    .c(_00013_),
    .y(_00014_)
  );
  al_nand2 _04587_ (
    .a(\DFF_311.Q ),
    .b(\DFF_733.Q ),
    .y(_00015_)
  );
  al_aoi21ttf _04588_ (
    .a(\DFF_1403.Q ),
    .b(\DFF_399.Q ),
    .c(_00015_),
    .y(_00016_)
  );
  al_and3 _04589_ (
    .a(_00014_),
    .b(_00016_),
    .c(_00012_),
    .y(g32185)
  );
  al_and2ft _04590_ (
    .a(\DFF_1127.Q ),
    .b(\DFF_646.Q ),
    .y(g25259)
  );
  al_inv _04591_ (
    .a(\DFF_994.Q ),
    .y(g23002)
  );
  al_and2ft _04592_ (
    .a(\DFF_794.Q ),
    .b(\DFF_1344.Q ),
    .y(g25167)
  );
  al_nand2 _04593_ (
    .a(g113),
    .b(\DFF_881.Q ),
    .y(g31656)
  );
  al_oa21ftt _04594_ (
    .a(\DFF_746.Q ),
    .b(\DFF_931.Q ),
    .c(\DFF_845.Q ),
    .y(_00017_)
  );
  al_oai21 _04595_ (
    .a(\DFF_319.Q ),
    .b(\DFF_746.Q ),
    .c(_00017_),
    .y(_00018_)
  );
  al_and3fft _04596_ (
    .a(\DFF_845.Q ),
    .b(\DFF_746.Q ),
    .c(\DFF_1.Q ),
    .y(_00019_)
  );
  al_nand3ftt _04597_ (
    .a(\DFF_845.Q ),
    .b(\DFF_1288.Q ),
    .c(\DFF_746.Q ),
    .y(_00020_)
  );
  al_and3ftt _04598_ (
    .a(_00019_),
    .b(_00020_),
    .c(_00018_),
    .y(\DFF_1111.D )
  );
  al_inv _04599_ (
    .a(\DFF_489.Q ),
    .y(g23612)
  );
  al_or3 _04600_ (
    .a(\DFF_619.Q ),
    .b(\DFF_761.Q ),
    .c(\DFF_1222.Q ),
    .y(_00021_)
  );
  al_and3fft _04601_ (
    .a(\DFF_512.Q ),
    .b(_00021_),
    .c(\DFF_790.Q ),
    .y(_00022_)
  );
  al_and3fft _04602_ (
    .a(\DFF_355.Q ),
    .b(\DFF_1229.Q ),
    .c(\DFF_547.Q ),
    .y(_00023_)
  );
  al_and3fft _04603_ (
    .a(\DFF_547.Q ),
    .b(\DFF_1229.Q ),
    .c(\DFF_355.Q ),
    .y(_00024_)
  );
  al_nor3fft _04604_ (
    .a(\DFF_512.Q ),
    .b(\DFF_790.Q ),
    .c(_00021_),
    .y(_00025_)
  );
  al_nand2 _04605_ (
    .a(_00024_),
    .b(_00025_),
    .y(_00026_)
  );
  al_aoi21ttf _04606_ (
    .a(_00022_),
    .b(_00023_),
    .c(_00026_),
    .y(_00027_)
  );
  al_inv _04607_ (
    .a(\DFF_790.Q ),
    .y(_00028_)
  );
  al_nor2 _04608_ (
    .a(\DFF_619.Q ),
    .b(\DFF_1222.Q ),
    .y(_00029_)
  );
  al_nand3fft _04609_ (
    .a(\DFF_761.Q ),
    .b(\DFF_512.Q ),
    .c(_00029_),
    .y(_00030_)
  );
  al_and3fft _04610_ (
    .a(_00028_),
    .b(_00030_),
    .c(_00024_),
    .y(_00031_)
  );
  al_and3ftt _04611_ (
    .a(\DFF_355.Q ),
    .b(\DFF_547.Q ),
    .c(\DFF_1229.Q ),
    .y(_00032_)
  );
  al_nand2ft _04612_ (
    .a(\DFF_512.Q ),
    .b(\DFF_619.Q ),
    .y(_00033_)
  );
  al_nor3fft _04613_ (
    .a(\DFF_761.Q ),
    .b(\DFF_1222.Q ),
    .c(_00033_),
    .y(_00034_)
  );
  al_and3 _04614_ (
    .a(\DFF_790.Q ),
    .b(_00032_),
    .c(_00034_),
    .y(_00035_)
  );
  al_and2ft _04615_ (
    .a(\DFF_1229.Q ),
    .b(\DFF_547.Q ),
    .y(_00036_)
  );
  al_nand3ftt _04616_ (
    .a(\DFF_790.Q ),
    .b(\DFF_355.Q ),
    .c(_00036_),
    .y(_00037_)
  );
  al_ao21ftf _04617_ (
    .a(_00023_),
    .b(_00037_),
    .c(_00034_),
    .y(_00038_)
  );
  al_and3fft _04618_ (
    .a(_00031_),
    .b(_00035_),
    .c(_00038_),
    .y(_00039_)
  );
  al_ao21 _04619_ (
    .a(_00027_),
    .b(_00039_),
    .c(_00005_),
    .y(_00040_)
  );
  al_or3 _04620_ (
    .a(\DFF_512.Q ),
    .b(\DFF_790.Q ),
    .c(_00021_),
    .y(_00041_)
  );
  al_or3ftt _04621_ (
    .a(_00023_),
    .b(_00005_),
    .c(_00041_),
    .y(_00042_)
  );
  al_or3fft _04622_ (
    .a(\DFF_236.Q ),
    .b(_00023_),
    .c(_00041_),
    .y(_00043_)
  );
  al_inv _04623_ (
    .a(\DFF_899.Q ),
    .y(_00044_)
  );
  al_and3 _04624_ (
    .a(_00028_),
    .b(_00023_),
    .c(_00034_),
    .y(_00045_)
  );
  al_and2 _04625_ (
    .a(\DFF_761.Q ),
    .b(\DFF_1222.Q ),
    .y(_00046_)
  );
  al_and3ftt _04626_ (
    .a(_00033_),
    .b(_00023_),
    .c(_00046_),
    .y(_00047_)
  );
  al_nand3 _04627_ (
    .a(\DFF_790.Q ),
    .b(\DFF_1336.Q ),
    .c(_00047_),
    .y(_00048_)
  );
  al_ao21ftf _04628_ (
    .a(_00044_),
    .b(_00045_),
    .c(_00048_),
    .y(_00049_)
  );
  al_and3 _04629_ (
    .a(\DFF_1182.Q ),
    .b(_00023_),
    .c(_00022_),
    .y(_00050_)
  );
  al_ao21 _04630_ (
    .a(\DFF_1245.Q ),
    .b(_00031_),
    .c(_00050_),
    .y(_00051_)
  );
  al_nor3ftt _04631_ (
    .a(_00043_),
    .b(_00051_),
    .c(_00049_),
    .y(_00052_)
  );
  al_ao21 _04632_ (
    .a(_00042_),
    .b(_00040_),
    .c(_00052_),
    .y(_00053_)
  );
  al_or3 _04633_ (
    .a(\DFF_547.Q ),
    .b(\DFF_355.Q ),
    .c(\DFF_1229.Q ),
    .y(_00054_)
  );
  al_or3 _04634_ (
    .a(\DFF_512.Q ),
    .b(_00021_),
    .c(_00054_),
    .y(_00055_)
  );
  al_aoi21ftf _04635_ (
    .a(_00054_),
    .b(_00025_),
    .c(_00055_),
    .y(_00056_)
  );
  al_and3fft _04636_ (
    .a(\DFF_790.Q ),
    .b(_00021_),
    .c(\DFF_512.Q ),
    .y(_00057_)
  );
  al_and3fft _04637_ (
    .a(\DFF_547.Q ),
    .b(\DFF_355.Q ),
    .c(\DFF_1229.Q ),
    .y(_00058_)
  );
  al_oai21ftt _04638_ (
    .a(_00041_),
    .b(_00057_),
    .c(_00058_),
    .y(_00059_)
  );
  al_aoi21 _04639_ (
    .a(_00056_),
    .b(_00059_),
    .c(_00005_),
    .y(_00060_)
  );
  al_and3fft _04640_ (
    .a(\DFF_790.Q ),
    .b(_00030_),
    .c(_00058_),
    .y(_00061_)
  );
  al_aoi21ftf _04641_ (
    .a(\DFF_844.Q ),
    .b(g35),
    .c(_00061_),
    .y(_00062_)
  );
  al_and2ft _04642_ (
    .a(_00054_),
    .b(_00025_),
    .y(_00063_)
  );
  al_aoi21ftf _04643_ (
    .a(\DFF_50.Q ),
    .b(g35),
    .c(_00063_),
    .y(_00064_)
  );
  al_inv _04644_ (
    .a(\DFF_162.Q ),
    .y(_00065_)
  );
  al_inv _04645_ (
    .a(g35),
    .y(_00066_)
  );
  al_and2 _04646_ (
    .a(_00058_),
    .b(_00057_),
    .y(_00067_)
  );
  al_ao21ftf _04647_ (
    .a(_00066_),
    .b(_00065_),
    .c(_00067_),
    .y(_00068_)
  );
  al_nand3fft _04648_ (
    .a(_00062_),
    .b(_00064_),
    .c(_00068_),
    .y(_00069_)
  );
  al_nand2 _04649_ (
    .a(_00060_),
    .b(_00069_),
    .y(_00070_)
  );
  al_nand3ftt _04650_ (
    .a(\DFF_547.Q ),
    .b(\DFF_355.Q ),
    .c(\DFF_1229.Q ),
    .y(_00071_)
  );
  al_and3fft _04651_ (
    .a(_00071_),
    .b(_00005_),
    .c(_00022_),
    .y(_00072_)
  );
  al_nor2 _04652_ (
    .a(g56),
    .b(g53),
    .y(_00073_)
  );
  al_nand3ftt _04653_ (
    .a(\DFF_355.Q ),
    .b(\DFF_547.Q ),
    .c(\DFF_1229.Q ),
    .y(_00074_)
  );
  al_and3ftt _04654_ (
    .a(_00074_),
    .b(_00073_),
    .c(_00004_),
    .y(_00075_)
  );
  al_nand3 _04655_ (
    .a(\DFF_657.Q ),
    .b(_00057_),
    .c(_00075_),
    .y(_00076_)
  );
  al_inv _04656_ (
    .a(g53),
    .y(_00077_)
  );
  al_aoi21ftf _04657_ (
    .a(g56),
    .b(_00004_),
    .c(_00077_),
    .y(_00078_)
  );
  al_aoi21ttf _04658_ (
    .a(\DFF_477.Q ),
    .b(_00078_),
    .c(_00076_),
    .y(_00079_)
  );
  al_aoi21ttf _04659_ (
    .a(\DFF_721.Q ),
    .b(_00072_),
    .c(_00079_),
    .y(_00080_)
  );
  al_inv _04660_ (
    .a(\DFF_948.Q ),
    .y(_00081_)
  );
  al_or3ftt _04661_ (
    .a(_00024_),
    .b(_00005_),
    .c(_00041_),
    .y(_00082_)
  );
  al_or3fft _04662_ (
    .a(_00081_),
    .b(\DFF_595.Q ),
    .c(_00082_),
    .y(_00083_)
  );
  al_nor3fft _04663_ (
    .a(_00073_),
    .b(_00004_),
    .c(_00041_),
    .y(_00084_)
  );
  al_and2ft _04664_ (
    .a(_00071_),
    .b(_00084_),
    .y(_00085_)
  );
  al_aoi21ttf _04665_ (
    .a(\DFF_677.Q ),
    .b(_00085_),
    .c(_00083_),
    .y(_00086_)
  );
  al_nor3ftt _04666_ (
    .a(_00032_),
    .b(_00005_),
    .c(_00041_),
    .y(_00087_)
  );
  al_inv _04667_ (
    .a(\DFF_1046.Q ),
    .y(_00088_)
  );
  al_nor3fft _04668_ (
    .a(_00058_),
    .b(_00022_),
    .c(_00005_),
    .y(_00089_)
  );
  al_nand3fft _04669_ (
    .a(\DFF_1242.Q ),
    .b(_00088_),
    .c(_00089_),
    .y(_00090_)
  );
  al_ao21ttf _04670_ (
    .a(\DFF_75.Q ),
    .b(_00087_),
    .c(_00090_),
    .y(_00091_)
  );
  al_and3ftt _04671_ (
    .a(_00091_),
    .b(_00080_),
    .c(_00086_),
    .y(_00092_)
  );
  al_nand3 _04672_ (
    .a(_00070_),
    .b(_00092_),
    .c(_00053_),
    .y(\DFF_1222.D )
  );
  al_nand3 _04673_ (
    .a(\DFF_364.Q ),
    .b(_00023_),
    .c(_00022_),
    .y(_00093_)
  );
  al_or3fft _04674_ (
    .a(\DFF_69.Q ),
    .b(_00023_),
    .c(_00041_),
    .y(_00094_)
  );
  al_inv _04675_ (
    .a(\DFF_531.Q ),
    .y(_00095_)
  );
  al_nand3 _04676_ (
    .a(\DFF_790.Q ),
    .b(\DFF_15.Q ),
    .c(_00047_),
    .y(_00096_)
  );
  al_aoi21ftf _04677_ (
    .a(_00095_),
    .b(_00045_),
    .c(_00096_),
    .y(_00097_)
  );
  al_and3 _04678_ (
    .a(_00093_),
    .b(_00094_),
    .c(_00097_),
    .y(_00098_)
  );
  al_ao21 _04679_ (
    .a(_00042_),
    .b(_00040_),
    .c(_00098_),
    .y(_00099_)
  );
  al_inv _04680_ (
    .a(\DFF_1090.Q ),
    .y(_00100_)
  );
  al_ao21ftf _04681_ (
    .a(_00066_),
    .b(_00100_),
    .c(_00067_),
    .y(_00101_)
  );
  al_aoi21ftf _04682_ (
    .a(\DFF_789.Q ),
    .b(g35),
    .c(_00063_),
    .y(_00102_)
  );
  al_ao21ftf _04683_ (
    .a(\DFF_338.Q ),
    .b(g35),
    .c(_00061_),
    .y(_00103_)
  );
  al_or3fft _04684_ (
    .a(_00028_),
    .b(\DFF_593.Q ),
    .c(_00055_),
    .y(_00104_)
  );
  al_nor3fft _04685_ (
    .a(_00104_),
    .b(_00103_),
    .c(_00102_),
    .y(_00105_)
  );
  al_ao21ttf _04686_ (
    .a(_00101_),
    .b(_00105_),
    .c(_00060_),
    .y(_00106_)
  );
  al_or3fft _04687_ (
    .a(\DFF_1323.Q ),
    .b(_00081_),
    .c(_00082_),
    .y(_00107_)
  );
  al_nand3 _04688_ (
    .a(\DFF_144.Q ),
    .b(_00057_),
    .c(_00075_),
    .y(_00108_)
  );
  al_nand3 _04689_ (
    .a(\DFF_514.Q ),
    .b(_00077_),
    .c(_00005_),
    .y(_00109_)
  );
  al_and3 _04690_ (
    .a(_00108_),
    .b(_00109_),
    .c(_00107_),
    .y(_00110_)
  );
  al_nand3ftt _04691_ (
    .a(_00071_),
    .b(\DFF_1157.Q ),
    .c(_00084_),
    .y(_00111_)
  );
  al_ao21ttf _04692_ (
    .a(\DFF_276.Q ),
    .b(_00072_),
    .c(_00111_),
    .y(_00112_)
  );
  al_inv _04693_ (
    .a(\DFF_1136.Q ),
    .y(_00113_)
  );
  al_nand3fft _04694_ (
    .a(\DFF_1242.Q ),
    .b(_00113_),
    .c(_00089_),
    .y(_00114_)
  );
  al_aoi21ttf _04695_ (
    .a(\DFF_64.Q ),
    .b(_00087_),
    .c(_00114_),
    .y(_00115_)
  );
  al_and3ftt _04696_ (
    .a(_00112_),
    .b(_00110_),
    .c(_00115_),
    .y(_00116_)
  );
  al_and2 _04697_ (
    .a(_00116_),
    .b(_00106_),
    .y(_00117_)
  );
  al_ao21ttf _04698_ (
    .a(_00099_),
    .b(_00117_),
    .c(\DFF_1222.D ),
    .y(_00118_)
  );
  al_or3fft _04699_ (
    .a(_00099_),
    .b(_00117_),
    .c(\DFF_1222.D ),
    .y(_00119_)
  );
  al_nand2ft _04700_ (
    .a(\DFF_506.Q ),
    .b(g35),
    .y(_00120_)
  );
  al_or3 _04701_ (
    .a(\DFF_770.Q ),
    .b(_00054_),
    .c(_00041_),
    .y(_00121_)
  );
  al_ao21ttf _04702_ (
    .a(_00120_),
    .b(_00067_),
    .c(_00121_),
    .y(_00122_)
  );
  al_nand2ft _04703_ (
    .a(\DFF_89.Q ),
    .b(g35),
    .y(_00123_)
  );
  al_or3fft _04704_ (
    .a(_00058_),
    .b(_00123_),
    .c(_00041_),
    .y(_00124_)
  );
  al_nand2ft _04705_ (
    .a(\DFF_28.Q ),
    .b(g35),
    .y(_00125_)
  );
  al_and3ftt _04706_ (
    .a(_00054_),
    .b(_00125_),
    .c(_00025_),
    .y(_00126_)
  );
  al_nand2ft _04707_ (
    .a(\DFF_1200.Q ),
    .b(g35),
    .y(_00127_)
  );
  al_or3fft _04708_ (
    .a(\DFF_790.Q ),
    .b(_00127_),
    .c(_00055_),
    .y(_00128_)
  );
  al_and3ftt _04709_ (
    .a(_00126_),
    .b(_00124_),
    .c(_00128_),
    .y(_00129_)
  );
  al_aoi21ftf _04710_ (
    .a(_00122_),
    .b(_00129_),
    .c(_00060_),
    .y(_00130_)
  );
  al_nand3 _04711_ (
    .a(\DFF_1067.Q ),
    .b(_00057_),
    .c(_00075_),
    .y(_00131_)
  );
  al_nand3 _04712_ (
    .a(\DFF_1340.Q ),
    .b(_00022_),
    .c(_00075_),
    .y(_00132_)
  );
  al_nand3 _04713_ (
    .a(\DFF_1012.Q ),
    .b(_00077_),
    .c(_00005_),
    .y(_00133_)
  );
  al_nand3 _04714_ (
    .a(_00133_),
    .b(_00131_),
    .c(_00132_),
    .y(_00134_)
  );
  al_inv _04715_ (
    .a(\DFF_195.Q ),
    .y(_00135_)
  );
  al_inv _04716_ (
    .a(\DFF_1000.Q ),
    .y(_00136_)
  );
  al_and3fft _04717_ (
    .a(\DFF_790.Q ),
    .b(_00030_),
    .c(_00023_),
    .y(_00137_)
  );
  al_nand3fft _04718_ (
    .a(_00136_),
    .b(_00005_),
    .c(_00137_),
    .y(_00138_)
  );
  al_ao21ftf _04719_ (
    .a(_00082_),
    .b(_00135_),
    .c(_00138_),
    .y(_00139_)
  );
  al_nand3 _04720_ (
    .a(\DFF_507.Q ),
    .b(_00032_),
    .c(_00084_),
    .y(_00140_)
  );
  al_aoi21ftf _04721_ (
    .a(\DFF_453.Q ),
    .b(_00089_),
    .c(_00140_),
    .y(_00141_)
  );
  al_nand3fft _04722_ (
    .a(_00134_),
    .b(_00139_),
    .c(_00141_),
    .y(_00142_)
  );
  al_nor3fft _04723_ (
    .a(\DFF_790.Q ),
    .b(_00046_),
    .c(_00033_),
    .y(_00143_)
  );
  al_aoi21ftf _04724_ (
    .a(_00074_),
    .b(_00143_),
    .c(_00038_),
    .y(_00144_)
  );
  al_nand3ftt _04725_ (
    .a(_00031_),
    .b(_00027_),
    .c(_00144_),
    .y(_00145_)
  );
  al_and3 _04726_ (
    .a(\DFF_311.Q ),
    .b(_00023_),
    .c(_00143_),
    .y(_00146_)
  );
  al_and3 _04727_ (
    .a(\DFF_1301.Q ),
    .b(_00024_),
    .c(_00025_),
    .y(_00147_)
  );
  al_ao21 _04728_ (
    .a(\DFF_881.Q ),
    .b(_00031_),
    .c(_00147_),
    .y(_00148_)
  );
  al_and3 _04729_ (
    .a(\DFF_749.Q ),
    .b(_00023_),
    .c(_00022_),
    .y(_00149_)
  );
  al_aoi21 _04730_ (
    .a(\DFF_733.Q ),
    .b(_00045_),
    .c(_00149_),
    .y(_00150_)
  );
  al_nand3fft _04731_ (
    .a(_00146_),
    .b(_00148_),
    .c(_00150_),
    .y(_00151_)
  );
  al_nand3 _04732_ (
    .a(\DFF_748.D ),
    .b(_00145_),
    .c(_00151_),
    .y(_00152_)
  );
  al_nand3fft _04733_ (
    .a(_00130_),
    .b(_00142_),
    .c(_00152_),
    .y(\DFF_1229.D )
  );
  al_aoi21 _04734_ (
    .a(_00027_),
    .b(_00039_),
    .c(_00005_),
    .y(_00153_)
  );
  al_and3 _04735_ (
    .a(\DFF_790.Q ),
    .b(\DFF_1151.Q ),
    .c(_00047_),
    .y(_00154_)
  );
  al_ao21 _04736_ (
    .a(\DFF_95.Q ),
    .b(_00045_),
    .c(_00035_),
    .y(_00155_)
  );
  al_nand3 _04737_ (
    .a(\DFF_757.Q ),
    .b(_00023_),
    .c(_00022_),
    .y(_00156_)
  );
  al_nand3 _04738_ (
    .a(\DFF_994.Q ),
    .b(_00024_),
    .c(_00025_),
    .y(_00157_)
  );
  al_and3 _04739_ (
    .a(\DFF_1035.Q ),
    .b(_00024_),
    .c(_00022_),
    .y(_00158_)
  );
  al_and3ftt _04740_ (
    .a(_00158_),
    .b(_00156_),
    .c(_00157_),
    .y(_00159_)
  );
  al_nand3fft _04741_ (
    .a(_00154_),
    .b(_00155_),
    .c(_00159_),
    .y(_00160_)
  );
  al_nand3fft _04742_ (
    .a(\DFF_177.Q ),
    .b(_00071_),
    .c(_00084_),
    .y(_00161_)
  );
  al_aoi21ftf _04743_ (
    .a(_00082_),
    .b(\DFF_948.Q ),
    .c(_00161_),
    .y(_00162_)
  );
  al_ao21ftf _04744_ (
    .a(\DFF_231.Q ),
    .b(_00072_),
    .c(_00162_),
    .y(_00163_)
  );
  al_aoi21 _04745_ (
    .a(_00160_),
    .b(_00153_),
    .c(_00163_),
    .y(_00164_)
  );
  al_aoi21ftf _04746_ (
    .a(\DFF_328.Q ),
    .b(g35),
    .c(_00063_),
    .y(_00165_)
  );
  al_and3fft _04747_ (
    .a(_00054_),
    .b(_00041_),
    .c(\DFF_1391.Q ),
    .y(_00166_)
  );
  al_nand2ft _04748_ (
    .a(\DFF_560.Q ),
    .b(g35),
    .y(_00167_)
  );
  al_and3 _04749_ (
    .a(_00058_),
    .b(_00167_),
    .c(_00057_),
    .y(_00168_)
  );
  al_nand2ft _04750_ (
    .a(\DFF_812.Q ),
    .b(g35),
    .y(_00169_)
  );
  al_or3fft _04751_ (
    .a(_00058_),
    .b(_00169_),
    .c(_00041_),
    .y(_00170_)
  );
  al_nand2ft _04752_ (
    .a(\DFF_661.Q ),
    .b(g35),
    .y(_00171_)
  );
  al_or3fft _04753_ (
    .a(\DFF_790.Q ),
    .b(_00171_),
    .c(_00055_),
    .y(_00172_)
  );
  al_and3ftt _04754_ (
    .a(_00168_),
    .b(_00170_),
    .c(_00172_),
    .y(_00173_)
  );
  al_nand3fft _04755_ (
    .a(_00166_),
    .b(_00165_),
    .c(_00173_),
    .y(_00174_)
  );
  al_and3 _04756_ (
    .a(\DFF_1322.Q ),
    .b(_00077_),
    .c(_00005_),
    .y(_00175_)
  );
  al_and3 _04757_ (
    .a(\DFF_25.Q ),
    .b(_00023_),
    .c(_00084_),
    .y(_00176_)
  );
  al_and3 _04758_ (
    .a(\DFF_1417.Q ),
    .b(_00022_),
    .c(_00075_),
    .y(_00177_)
  );
  al_aoi21 _04759_ (
    .a(\DFF_1242.Q ),
    .b(_00089_),
    .c(_00177_),
    .y(_00178_)
  );
  al_nand3fft _04760_ (
    .a(_00175_),
    .b(_00176_),
    .c(_00178_),
    .y(_00179_)
  );
  al_aoi21 _04761_ (
    .a(_00060_),
    .b(_00174_),
    .c(_00179_),
    .y(_00180_)
  );
  al_ao21 _04762_ (
    .a(_00180_),
    .b(_00164_),
    .c(\DFF_1229.D ),
    .y(_00181_)
  );
  al_and3 _04763_ (
    .a(_00180_),
    .b(_00164_),
    .c(\DFF_1229.D ),
    .y(_00182_)
  );
  al_nand2ft _04764_ (
    .a(_00182_),
    .b(_00181_),
    .y(_00183_)
  );
  al_ao21 _04765_ (
    .a(_00118_),
    .b(_00119_),
    .c(_00183_),
    .y(_00184_)
  );
  al_and3 _04766_ (
    .a(_00118_),
    .b(_00119_),
    .c(_00183_),
    .y(_00185_)
  );
  al_nand2ft _04767_ (
    .a(_00185_),
    .b(_00184_),
    .y(_00186_)
  );
  al_aoi21ftf _04768_ (
    .a(\DFF_876.Q ),
    .b(g35),
    .c(_00063_),
    .y(_00187_)
  );
  al_or3 _04769_ (
    .a(\DFF_790.Q ),
    .b(_00054_),
    .c(_00030_),
    .y(_00188_)
  );
  al_inv _04770_ (
    .a(\DFF_874.Q ),
    .y(_00189_)
  );
  al_ao21ftf _04771_ (
    .a(_00066_),
    .b(_00189_),
    .c(_00061_),
    .y(_00190_)
  );
  al_ao21ftf _04772_ (
    .a(_00188_),
    .b(\DFF_715.Q ),
    .c(_00190_),
    .y(_00191_)
  );
  al_and3fft _04773_ (
    .a(_00054_),
    .b(_00030_),
    .c(\DFF_790.Q ),
    .y(_00192_)
  );
  al_and2ft _04774_ (
    .a(\DFF_896.Q ),
    .b(g35),
    .y(_00193_)
  );
  al_ao21ftf _04775_ (
    .a(\DFF_88.Q ),
    .b(g35),
    .c(_00067_),
    .y(_00194_)
  );
  al_aoi21ftf _04776_ (
    .a(_00193_),
    .b(_00192_),
    .c(_00194_),
    .y(_00195_)
  );
  al_nand3fft _04777_ (
    .a(_00187_),
    .b(_00191_),
    .c(_00195_),
    .y(_00196_)
  );
  al_nand2 _04778_ (
    .a(_00060_),
    .b(_00196_),
    .y(_00197_)
  );
  al_or3fft _04779_ (
    .a(\DFF_413.Q ),
    .b(_00034_),
    .c(_00037_),
    .y(_00198_)
  );
  al_oai21ftt _04780_ (
    .a(g100),
    .b(_00026_),
    .c(_00198_),
    .y(_00199_)
  );
  al_aoi21 _04781_ (
    .a(\DFF_1178.Q ),
    .b(_00031_),
    .c(_00035_),
    .y(_00200_)
  );
  al_ao21ftf _04782_ (
    .a(_00199_),
    .b(_00200_),
    .c(_00153_),
    .y(_00201_)
  );
  al_nor3fft _04783_ (
    .a(_00032_),
    .b(_00057_),
    .c(_00005_),
    .y(_00202_)
  );
  al_nand3 _04784_ (
    .a(\DFF_1041.Q ),
    .b(_00022_),
    .c(_00075_),
    .y(_00203_)
  );
  al_aoi21ttf _04785_ (
    .a(\DFF_206.Q ),
    .b(_00078_),
    .c(_00203_),
    .y(_00204_)
  );
  al_aoi21ttf _04786_ (
    .a(\DFF_1319.Q ),
    .b(_00202_),
    .c(_00204_),
    .y(_00205_)
  );
  al_nand3ftt _04787_ (
    .a(_00005_),
    .b(\DFF_767.Q ),
    .c(_00137_),
    .y(_00206_)
  );
  al_ao21ttf _04788_ (
    .a(\DFF_1314.Q ),
    .b(_00089_),
    .c(_00206_),
    .y(_00207_)
  );
  al_nand3 _04789_ (
    .a(\DFF_445.Q ),
    .b(_00032_),
    .c(_00084_),
    .y(_00208_)
  );
  al_aoi21ftf _04790_ (
    .a(_00082_),
    .b(\DFF_932.Q ),
    .c(_00208_),
    .y(_00209_)
  );
  al_and3ftt _04791_ (
    .a(_00207_),
    .b(_00209_),
    .c(_00205_),
    .y(_00210_)
  );
  al_nand3 _04792_ (
    .a(_00210_),
    .b(_00201_),
    .c(_00197_),
    .y(\DFF_512.D )
  );
  al_and3 _04793_ (
    .a(_00028_),
    .b(\DFF_399.Q ),
    .c(_00047_),
    .y(_00211_)
  );
  al_and3 _04794_ (
    .a(\DFF_790.Q ),
    .b(_00023_),
    .c(_00034_),
    .y(_00212_)
  );
  al_or3fft _04795_ (
    .a(\DFF_197.Q ),
    .b(_00034_),
    .c(_00037_),
    .y(_00213_)
  );
  al_ao21ttf _04796_ (
    .a(\DFF_1403.Q ),
    .b(_00212_),
    .c(_00213_),
    .y(_00214_)
  );
  al_and3fft _04797_ (
    .a(_00028_),
    .b(_00030_),
    .c(_00023_),
    .y(_00215_)
  );
  al_and3 _04798_ (
    .a(g127),
    .b(_00024_),
    .c(_00022_),
    .y(_00216_)
  );
  al_aoi21 _04799_ (
    .a(\DFF_242.Q ),
    .b(_00215_),
    .c(_00216_),
    .y(_00217_)
  );
  al_aoi21ftf _04800_ (
    .a(_00026_),
    .b(g92),
    .c(_00217_),
    .y(_00218_)
  );
  al_nand3fft _04801_ (
    .a(_00211_),
    .b(_00214_),
    .c(_00218_),
    .y(_00219_)
  );
  al_nand3 _04802_ (
    .a(\DFF_420.Q ),
    .b(_00077_),
    .c(_00005_),
    .y(_00220_)
  );
  al_aoi21ttf _04803_ (
    .a(\DFF_127.Q ),
    .b(_00089_),
    .c(_00220_),
    .y(_00221_)
  );
  al_ao21ttf _04804_ (
    .a(\DFF_1270.Q ),
    .b(_00202_),
    .c(_00221_),
    .y(_00222_)
  );
  al_aoi21 _04805_ (
    .a(_00153_),
    .b(_00219_),
    .c(_00222_),
    .y(_00223_)
  );
  al_aoi21ftf _04806_ (
    .a(\DFF_728.Q ),
    .b(g35),
    .c(_00067_),
    .y(_00224_)
  );
  al_aoi21ftf _04807_ (
    .a(\DFF_175.Q ),
    .b(g35),
    .c(_00063_),
    .y(_00225_)
  );
  al_inv _04808_ (
    .a(\DFF_966.Q ),
    .y(_00226_)
  );
  al_ao21ftf _04809_ (
    .a(_00066_),
    .b(_00226_),
    .c(_00061_),
    .y(_00227_)
  );
  al_or3 _04810_ (
    .a(g23612),
    .b(_00054_),
    .c(_00041_),
    .y(_00228_)
  );
  al_aoi21ftf _04811_ (
    .a(\DFF_953.Q ),
    .b(g35),
    .c(_00192_),
    .y(_00229_)
  );
  al_nor3fft _04812_ (
    .a(_00228_),
    .b(_00227_),
    .c(_00229_),
    .y(_00230_)
  );
  al_nand3fft _04813_ (
    .a(_00224_),
    .b(_00225_),
    .c(_00230_),
    .y(_00231_)
  );
  al_and3 _04814_ (
    .a(\DFF_974.Q ),
    .b(_00022_),
    .c(_00075_),
    .y(_00232_)
  );
  al_or3ftt _04815_ (
    .a(_00023_),
    .b(_00005_),
    .c(_00041_),
    .y(_00233_)
  );
  al_and3 _04816_ (
    .a(\DFF_323.Q ),
    .b(_00024_),
    .c(_00084_),
    .y(_00234_)
  );
  al_aoi21ftt _04817_ (
    .a(_00233_),
    .b(\DFF_673.Q ),
    .c(_00234_),
    .y(_00235_)
  );
  al_nand3ftt _04818_ (
    .a(_00041_),
    .b(\DFF_941.Q ),
    .c(_00075_),
    .y(_00236_)
  );
  al_nand3ftt _04819_ (
    .a(_00232_),
    .b(_00236_),
    .c(_00235_),
    .y(_00237_)
  );
  al_aoi21 _04820_ (
    .a(_00060_),
    .b(_00231_),
    .c(_00237_),
    .y(_00238_)
  );
  al_or3fft _04821_ (
    .a(_00238_),
    .b(_00223_),
    .c(\DFF_512.D ),
    .y(_00239_)
  );
  al_aoi21ttf _04822_ (
    .a(_00238_),
    .b(_00223_),
    .c(\DFF_512.D ),
    .y(_00240_)
  );
  al_nand2ft _04823_ (
    .a(_00240_),
    .b(_00239_),
    .y(_00241_)
  );
  al_nand2ft _04824_ (
    .a(\DFF_157.Q ),
    .b(g35),
    .y(_00242_)
  );
  al_and3fft _04825_ (
    .a(_00054_),
    .b(_00041_),
    .c(\DFF_597.Q ),
    .y(_00243_)
  );
  al_aoi21 _04826_ (
    .a(_00242_),
    .b(_00063_),
    .c(_00243_),
    .y(_00244_)
  );
  al_ao21ftf _04827_ (
    .a(\DFF_751.Q ),
    .b(g35),
    .c(_00061_),
    .y(_00245_)
  );
  al_aoi21ftf _04828_ (
    .a(\DFF_21.Q ),
    .b(g35),
    .c(_00192_),
    .y(_00246_)
  );
  al_ao21ftf _04829_ (
    .a(\DFF_863.Q ),
    .b(g35),
    .c(_00067_),
    .y(_00247_)
  );
  al_and3ftt _04830_ (
    .a(_00246_),
    .b(_00245_),
    .c(_00247_),
    .y(_00248_)
  );
  al_ao21ttf _04831_ (
    .a(_00244_),
    .b(_00248_),
    .c(_00060_),
    .y(_00249_)
  );
  al_nand3 _04832_ (
    .a(\DFF_498.Q ),
    .b(_00057_),
    .c(_00075_),
    .y(_00250_)
  );
  al_aoi21ttf _04833_ (
    .a(\DFF_150.Q ),
    .b(_00078_),
    .c(_00250_),
    .y(_00251_)
  );
  al_aoi21ttf _04834_ (
    .a(\DFF_766.Q ),
    .b(_00072_),
    .c(_00251_),
    .y(_00252_)
  );
  al_or3fft _04835_ (
    .a(_00081_),
    .b(\DFF_774.Q ),
    .c(_00082_),
    .y(_00253_)
  );
  al_aoi21ttf _04836_ (
    .a(\DFF_161.Q ),
    .b(_00085_),
    .c(_00253_),
    .y(_00254_)
  );
  al_inv _04837_ (
    .a(\DFF_137.Q ),
    .y(_00255_)
  );
  al_nand3fft _04838_ (
    .a(\DFF_1242.Q ),
    .b(_00255_),
    .c(_00089_),
    .y(_00256_)
  );
  al_ao21ttf _04839_ (
    .a(\DFF_190.Q ),
    .b(_00087_),
    .c(_00256_),
    .y(_00257_)
  );
  al_and3ftt _04840_ (
    .a(_00257_),
    .b(_00252_),
    .c(_00254_),
    .y(_00258_)
  );
  al_nand3 _04841_ (
    .a(_00028_),
    .b(\DFF_155.Q ),
    .c(_00047_),
    .y(_00259_)
  );
  al_aoi21 _04842_ (
    .a(\DFF_1282.Q ),
    .b(_00212_),
    .c(_00035_),
    .y(_00260_)
  );
  al_inv _04843_ (
    .a(\DFF_223.Q ),
    .y(_00261_)
  );
  al_and3 _04844_ (
    .a(\DFF_706.Q ),
    .b(_00024_),
    .c(_00022_),
    .y(_00262_)
  );
  al_aoi21 _04845_ (
    .a(\DFF_1357.Q ),
    .b(_00137_),
    .c(_00262_),
    .y(_00263_)
  );
  al_aoi21ftf _04846_ (
    .a(_00261_),
    .b(_00215_),
    .c(_00263_),
    .y(_00264_)
  );
  al_nand3 _04847_ (
    .a(_00259_),
    .b(_00260_),
    .c(_00264_),
    .y(_00265_)
  );
  al_ao21ttf _04848_ (
    .a(_00040_),
    .b(_00233_),
    .c(_00265_),
    .y(_00266_)
  );
  al_and3 _04849_ (
    .a(_00258_),
    .b(_00249_),
    .c(_00266_),
    .y(_00267_)
  );
  al_oai21ftt _04850_ (
    .a(g54),
    .b(g56),
    .c(\DFF_621.Q ),
    .y(_00268_)
  );
  al_nand3 _04851_ (
    .a(\DFF_781.Q ),
    .b(_00023_),
    .c(_00022_),
    .y(_00269_)
  );
  al_inv _04852_ (
    .a(\DFF_852.Q ),
    .y(_00270_)
  );
  al_nand3 _04853_ (
    .a(\DFF_790.Q ),
    .b(\DFF_1289.Q ),
    .c(_00047_),
    .y(_00271_)
  );
  al_ao21ftf _04854_ (
    .a(_00270_),
    .b(_00045_),
    .c(_00271_),
    .y(_00272_)
  );
  al_nand3ftt _04855_ (
    .a(\DFF_1125.Q ),
    .b(_00024_),
    .c(_00022_),
    .y(_00273_)
  );
  al_ao21ttf _04856_ (
    .a(\DFF_608.Q ),
    .b(_00137_),
    .c(_00273_),
    .y(_00274_)
  );
  al_nor3ftt _04857_ (
    .a(_00269_),
    .b(_00274_),
    .c(_00272_),
    .y(_00275_)
  );
  al_ao21 _04858_ (
    .a(_00233_),
    .b(_00040_),
    .c(_00275_),
    .y(_00276_)
  );
  al_aoi21ftf _04859_ (
    .a(\DFF_119.Q ),
    .b(g35),
    .c(_00061_),
    .y(_00277_)
  );
  al_inv _04860_ (
    .a(\DFF_142.Q ),
    .y(_00278_)
  );
  al_ao21ftf _04861_ (
    .a(_00066_),
    .b(_00278_),
    .c(_00192_),
    .y(_00279_)
  );
  al_and2ft _04862_ (
    .a(\DFF_74.Q ),
    .b(g35),
    .y(_00280_)
  );
  al_ao21ftf _04863_ (
    .a(_00280_),
    .b(_00063_),
    .c(_00279_),
    .y(_00281_)
  );
  al_inv _04864_ (
    .a(\DFF_1235.Q ),
    .y(_00282_)
  );
  al_ao21ftf _04865_ (
    .a(_00066_),
    .b(_00282_),
    .c(_00067_),
    .y(_00283_)
  );
  al_aoi21ftf _04866_ (
    .a(_00188_),
    .b(\DFF_1253.Q ),
    .c(_00283_),
    .y(_00284_)
  );
  al_nand3fft _04867_ (
    .a(_00277_),
    .b(_00281_),
    .c(_00284_),
    .y(_00285_)
  );
  al_nand3 _04868_ (
    .a(\DFF_196.Q ),
    .b(_00057_),
    .c(_00075_),
    .y(_00286_)
  );
  al_aoi21ttf _04869_ (
    .a(\DFF_829.Q ),
    .b(_00078_),
    .c(_00286_),
    .y(_00287_)
  );
  al_aoi21ttf _04870_ (
    .a(\DFF_1193.Q ),
    .b(_00085_),
    .c(_00287_),
    .y(_00288_)
  );
  al_or3fft _04871_ (
    .a(_00081_),
    .b(\DFF_403.Q ),
    .c(_00082_),
    .y(_00289_)
  );
  al_ao21ttf _04872_ (
    .a(\DFF_855.Q ),
    .b(_00072_),
    .c(_00289_),
    .y(_00290_)
  );
  al_inv _04873_ (
    .a(\DFF_296.Q ),
    .y(_00291_)
  );
  al_nand3fft _04874_ (
    .a(\DFF_1242.Q ),
    .b(_00291_),
    .c(_00089_),
    .y(_00292_)
  );
  al_aoi21ttf _04875_ (
    .a(\DFF_80.Q ),
    .b(_00087_),
    .c(_00292_),
    .y(_00293_)
  );
  al_and3ftt _04876_ (
    .a(_00290_),
    .b(_00293_),
    .c(_00288_),
    .y(_00294_)
  );
  al_aoi21ttf _04877_ (
    .a(_00060_),
    .b(_00285_),
    .c(_00294_),
    .y(_00295_)
  );
  al_nand3 _04878_ (
    .a(_00268_),
    .b(_00276_),
    .c(_00295_),
    .y(_00296_)
  );
  al_ao21 _04879_ (
    .a(_00276_),
    .b(_00295_),
    .c(_00268_),
    .y(_00297_)
  );
  al_nand3 _04880_ (
    .a(_00267_),
    .b(_00296_),
    .c(_00297_),
    .y(_00298_)
  );
  al_ao21 _04881_ (
    .a(_00296_),
    .b(_00297_),
    .c(_00267_),
    .y(_00299_)
  );
  al_nand3 _04882_ (
    .a(_00298_),
    .b(_00299_),
    .c(_00241_),
    .y(_00300_)
  );
  al_ao21 _04883_ (
    .a(_00298_),
    .b(_00299_),
    .c(_00241_),
    .y(_00301_)
  );
  al_ao21ttf _04884_ (
    .a(_00300_),
    .b(_00301_),
    .c(_00186_),
    .y(_00302_)
  );
  al_and2ft _04885_ (
    .a(_00185_),
    .b(_00184_),
    .y(_00303_)
  );
  al_nand3 _04886_ (
    .a(_00300_),
    .b(_00301_),
    .c(_00303_),
    .y(_00304_)
  );
  al_nand2 _04887_ (
    .a(_00302_),
    .b(_00304_),
    .y(\DFF_1074.D )
  );
  al_nand3 _04888_ (
    .a(\DFF_748.Q ),
    .b(_00302_),
    .c(_00304_),
    .y(g34972)
  );
  al_nand3 _04889_ (
    .a(\DFF_748.Q ),
    .b(_00099_),
    .c(_00117_),
    .y(g34913)
  );
  al_nor2 _04890_ (
    .a(\DFF_860.Q ),
    .b(\DFF_1361.Q ),
    .y(_00305_)
  );
  al_or3 _04891_ (
    .a(\DFF_551.Q ),
    .b(\DFF_351.Q ),
    .c(\DFF_411.Q ),
    .y(_00306_)
  );
  al_or3fft _04892_ (
    .a(\DFF_154.Q ),
    .b(\DFF_1139.Q ),
    .c(_00306_),
    .y(_00307_)
  );
  al_or3 _04893_ (
    .a(\DFF_1204.Q ),
    .b(\DFF_1324.Q ),
    .c(\DFF_891.Q ),
    .y(_00308_)
  );
  al_aoi21 _04894_ (
    .a(_00305_),
    .b(_00307_),
    .c(_00308_),
    .y(g31521)
  );
  al_and2 _04895_ (
    .a(\DFF_449.Q ),
    .b(\DFF_846.Q ),
    .y(g25114)
  );
  al_nand3 _04896_ (
    .a(_00116_),
    .b(_00106_),
    .c(_00099_),
    .y(\DFF_619.D )
  );
  al_and2ft _04897_ (
    .a(g35),
    .b(\DFF_800.Q ),
    .y(\DFF_999.D )
  );
  al_and2ft _04898_ (
    .a(g35),
    .b(\DFF_1402.Q ),
    .y(\DFF_1165.D )
  );
  al_or2 _04899_ (
    .a(g23190),
    .b(\DFF_1229.D ),
    .y(g34925)
  );
  al_and2ft _04900_ (
    .a(g35),
    .b(\DFF_231.Q ),
    .y(\DFF_1402.D )
  );
  al_and2ft _04901_ (
    .a(g35),
    .b(\DFF_1292.Q ),
    .y(\DFF_1353.D )
  );
  al_nand3 _04902_ (
    .a(\DFF_748.Q ),
    .b(_00180_),
    .c(_00164_),
    .y(g34923)
  );
  al_inv _04903_ (
    .a(\DFF_736.Q ),
    .y(_00309_)
  );
  al_inv _04904_ (
    .a(\DFF_353.Q ),
    .y(_00310_)
  );
  al_nor2 _04905_ (
    .a(\DFF_47.Q ),
    .b(g73),
    .y(_00311_)
  );
  al_nand2 _04906_ (
    .a(\DFF_47.Q ),
    .b(g73),
    .y(_00312_)
  );
  al_nand2ft _04907_ (
    .a(_00311_),
    .b(_00312_),
    .y(_00313_)
  );
  al_nand2ft _04908_ (
    .a(\DFF_1145.Q ),
    .b(g72),
    .y(_00314_)
  );
  al_nand2ft _04909_ (
    .a(g72),
    .b(\DFF_1145.Q ),
    .y(_00315_)
  );
  al_and3 _04910_ (
    .a(_00314_),
    .b(_00315_),
    .c(_00313_),
    .y(_00316_)
  );
  al_and2 _04911_ (
    .a(_00310_),
    .b(_00316_),
    .y(_00317_)
  );
  al_aoi21 _04912_ (
    .a(\DFF_252.Q ),
    .b(_00317_),
    .c(_00309_),
    .y(g33894)
  );
  al_nand2 _04913_ (
    .a(_00238_),
    .b(_00223_),
    .y(\DFF_790.D )
  );
  al_inv _04914_ (
    .a(\DFF_591.Q ),
    .y(_00318_)
  );
  al_and3 _04915_ (
    .a(_00318_),
    .b(\DFF_353.Q ),
    .c(_00316_),
    .y(_00319_)
  );
  al_and2ft _04916_ (
    .a(\DFF_1010.Q ),
    .b(\DFF_1233.Q ),
    .y(_00320_)
  );
  al_and3 _04917_ (
    .a(\DFF_622.Q ),
    .b(_00320_),
    .c(_00319_),
    .y(_00321_)
  );
  al_inv _04918_ (
    .a(\DFF_622.Q ),
    .y(_00322_)
  );
  al_and3 _04919_ (
    .a(\DFF_591.Q ),
    .b(_00322_),
    .c(_00317_),
    .y(_00323_)
  );
  al_and2ft _04920_ (
    .a(\DFF_671.Q ),
    .b(\DFF_996.Q ),
    .y(_00324_)
  );
  al_ao21 _04921_ (
    .a(_00324_),
    .b(_00323_),
    .c(_00321_),
    .y(_00325_)
  );
  al_and3 _04922_ (
    .a(\DFF_591.Q ),
    .b(\DFF_622.Q ),
    .c(_00317_),
    .y(_00326_)
  );
  al_nand2ft _04923_ (
    .a(\DFF_759.Q ),
    .b(\DFF_620.Q ),
    .y(_00327_)
  );
  al_and3 _04924_ (
    .a(\DFF_591.Q ),
    .b(\DFF_353.Q ),
    .c(_00316_),
    .y(_00328_)
  );
  al_and2ft _04925_ (
    .a(\DFF_265.Q ),
    .b(\DFF_886.Q ),
    .y(_00329_)
  );
  al_nand3 _04926_ (
    .a(\DFF_622.Q ),
    .b(_00329_),
    .c(_00328_),
    .y(_00330_)
  );
  al_ao21ftf _04927_ (
    .a(_00327_),
    .b(_00326_),
    .c(_00330_),
    .y(_00331_)
  );
  al_and2ft _04928_ (
    .a(\DFF_402.Q ),
    .b(\DFF_505.Q ),
    .y(_00332_)
  );
  al_and3 _04929_ (
    .a(_00322_),
    .b(_00332_),
    .c(_00328_),
    .y(_00333_)
  );
  al_and3 _04930_ (
    .a(_00318_),
    .b(\DFF_622.Q ),
    .c(_00317_),
    .y(_00334_)
  );
  al_and2ft _04931_ (
    .a(\DFF_500.Q ),
    .b(\DFF_18.Q ),
    .y(_00335_)
  );
  al_aoi21 _04932_ (
    .a(_00335_),
    .b(_00334_),
    .c(_00333_),
    .y(_00336_)
  );
  al_and2ft _04933_ (
    .a(\DFF_1141.Q ),
    .b(\DFF_1047.Q ),
    .y(_00337_)
  );
  al_nand3 _04934_ (
    .a(_00322_),
    .b(_00337_),
    .c(_00319_),
    .y(_00338_)
  );
  al_and3 _04935_ (
    .a(_00318_),
    .b(_00322_),
    .c(_00317_),
    .y(_00339_)
  );
  al_nand2 _04936_ (
    .a(g25259),
    .b(_00339_),
    .y(_00340_)
  );
  al_and3 _04937_ (
    .a(_00338_),
    .b(_00340_),
    .c(_00336_),
    .y(_00341_)
  );
  al_nand3fft _04938_ (
    .a(_00325_),
    .b(_00331_),
    .c(_00341_),
    .y(\DFF_1181.D )
  );
  al_ao21 _04939_ (
    .a(\DFF_994.Q ),
    .b(g99),
    .c(g134),
    .y(_00342_)
  );
  al_and2 _04940_ (
    .a(g113),
    .b(_00342_),
    .y(_00343_)
  );
  al_or3fft _04941_ (
    .a(_00316_),
    .b(_00343_),
    .c(\DFF_1181.D ),
    .y(g34383)
  );
  al_and2ft _04942_ (
    .a(g35),
    .b(\DFF_611.Q ),
    .y(\DFF_1101.D )
  );
  al_or2 _04943_ (
    .a(g23190),
    .b(\DFF_1222.D ),
    .y(g34917)
  );
  al_and2ft _04944_ (
    .a(g35),
    .b(\DFF_799.Q ),
    .y(\DFF_908.D )
  );
  al_nor2 _04945_ (
    .a(\DFF_363.Q ),
    .b(\DFF_1103.Q ),
    .y(_00344_)
  );
  al_and3ftt _04946_ (
    .a(\DFF_90.Q ),
    .b(\DFF_698.Q ),
    .c(\DFF_1133.Q ),
    .y(_00345_)
  );
  al_and3ftt _04947_ (
    .a(\DFF_1057.Q ),
    .b(_00345_),
    .c(_00344_),
    .y(_00346_)
  );
  al_nand3ftt _04948_ (
    .a(\DFF_563.Q ),
    .b(\DFF_214.Q ),
    .c(_00346_),
    .y(_00347_)
  );
  al_nand2 _04949_ (
    .a(\DFF_711.Q ),
    .b(_00347_),
    .y(_00348_)
  );
  al_inv _04950_ (
    .a(_00348_),
    .y(g27831)
  );
  al_and2ft _04951_ (
    .a(g35),
    .b(\DFF_980.Q ),
    .y(\DFF_1305.D )
  );
  al_and2ft _04952_ (
    .a(g35),
    .b(\DFF_501.Q ),
    .y(\DFF_200.D )
  );
  al_or2 _04953_ (
    .a(g23190),
    .b(\DFF_512.D ),
    .y(g34915)
  );
  al_nor2 _04954_ (
    .a(\DFF_201.Q ),
    .b(g73),
    .y(_00349_)
  );
  al_nand2 _04955_ (
    .a(\DFF_201.Q ),
    .b(g73),
    .y(_00350_)
  );
  al_nand2ft _04956_ (
    .a(_00349_),
    .b(_00350_),
    .y(_00351_)
  );
  al_nand2ft _04957_ (
    .a(\DFF_508.Q ),
    .b(g72),
    .y(_00352_)
  );
  al_nand2ft _04958_ (
    .a(g72),
    .b(\DFF_508.Q ),
    .y(_00353_)
  );
  al_and3 _04959_ (
    .a(_00352_),
    .b(_00353_),
    .c(_00351_),
    .y(_00354_)
  );
  al_inv _04960_ (
    .a(\DFF_411.Q ),
    .y(_00355_)
  );
  al_inv _04961_ (
    .a(\DFF_351.Q ),
    .y(_00356_)
  );
  al_and3 _04962_ (
    .a(\DFF_551.Q ),
    .b(_00356_),
    .c(_00354_),
    .y(_00357_)
  );
  al_and3 _04963_ (
    .a(\DFF_519.Q ),
    .b(\DFF_385.Q ),
    .c(\DFF_393.Q ),
    .y(_00358_)
  );
  al_and3 _04964_ (
    .a(_00355_),
    .b(_00358_),
    .c(_00357_),
    .y(_00359_)
  );
  al_and3 _04965_ (
    .a(\DFF_551.Q ),
    .b(\DFF_351.Q ),
    .c(_00354_),
    .y(_00360_)
  );
  al_and3 _04966_ (
    .a(\DFF_587.Q ),
    .b(\DFF_473.Q ),
    .c(\DFF_467.Q ),
    .y(_00361_)
  );
  al_and3 _04967_ (
    .a(\DFF_411.Q ),
    .b(_00361_),
    .c(_00360_),
    .y(_00362_)
  );
  al_and2 _04968_ (
    .a(\DFF_411.Q ),
    .b(_00354_),
    .y(_00363_)
  );
  al_and2ft _04969_ (
    .a(\DFF_551.Q ),
    .b(\DFF_351.Q ),
    .y(_00364_)
  );
  al_and3 _04970_ (
    .a(\DFF_271.Q ),
    .b(\DFF_522.Q ),
    .c(\DFF_54.Q ),
    .y(_00365_)
  );
  al_nand3 _04971_ (
    .a(_00364_),
    .b(_00365_),
    .c(_00363_),
    .y(_00366_)
  );
  al_nor2 _04972_ (
    .a(\DFF_551.Q ),
    .b(\DFF_351.Q ),
    .y(_00367_)
  );
  al_and3 _04973_ (
    .a(\DFF_411.Q ),
    .b(_00367_),
    .c(_00354_),
    .y(_00368_)
  );
  al_and3 _04974_ (
    .a(\DFF_575.Q ),
    .b(\DFF_289.Q ),
    .c(\DFF_910.Q ),
    .y(_00369_)
  );
  al_and2 _04975_ (
    .a(_00369_),
    .b(_00368_),
    .y(_00370_)
  );
  al_and3ftt _04976_ (
    .a(_00306_),
    .b(g26801),
    .c(_00354_),
    .y(_00371_)
  );
  al_and3 _04977_ (
    .a(_00355_),
    .b(_00364_),
    .c(_00354_),
    .y(_00372_)
  );
  al_and3 _04978_ (
    .a(\DFF_1150.Q ),
    .b(\DFF_1273.Q ),
    .c(\DFF_1068.Q ),
    .y(_00373_)
  );
  al_aoi21 _04979_ (
    .a(_00373_),
    .b(_00372_),
    .c(_00371_),
    .y(_00374_)
  );
  al_and3ftt _04980_ (
    .a(_00370_),
    .b(_00366_),
    .c(_00374_),
    .y(_00375_)
  );
  al_and3 _04981_ (
    .a(\DFF_20.Q ),
    .b(\DFF_916.Q ),
    .c(\DFF_104.Q ),
    .y(_00376_)
  );
  al_nand3 _04982_ (
    .a(\DFF_411.Q ),
    .b(_00376_),
    .c(_00357_),
    .y(_00377_)
  );
  al_and3 _04983_ (
    .a(\DFF_1408.Q ),
    .b(\DFF_245.Q ),
    .c(\DFF_199.Q ),
    .y(_00378_)
  );
  al_nand3 _04984_ (
    .a(_00355_),
    .b(_00378_),
    .c(_00360_),
    .y(_00379_)
  );
  al_and3 _04985_ (
    .a(_00377_),
    .b(_00379_),
    .c(_00375_),
    .y(_00380_)
  );
  al_nand3fft _04986_ (
    .a(_00359_),
    .b(_00362_),
    .c(_00380_),
    .y(\DFF_304.D )
  );
  al_or3fft _04987_ (
    .a(_00343_),
    .b(_00354_),
    .c(\DFF_304.D ),
    .y(g33659)
  );
  al_and2ft _04988_ (
    .a(g35),
    .b(\DFF_1381.Q ),
    .y(g21727)
  );
  al_nand3 _04989_ (
    .a(_00258_),
    .b(_00249_),
    .c(_00266_),
    .y(\DFF_547.D )
  );
  al_nand2 _04990_ (
    .a(_00276_),
    .b(_00295_),
    .y(\DFF_761.D )
  );
  al_nor2 _04991_ (
    .a(\DFF_115.Q ),
    .b(g73),
    .y(_00381_)
  );
  al_nand2 _04992_ (
    .a(\DFF_115.Q ),
    .b(g73),
    .y(_00382_)
  );
  al_nand2ft _04993_ (
    .a(_00381_),
    .b(_00382_),
    .y(_00383_)
  );
  al_nand2ft _04994_ (
    .a(\DFF_1084.Q ),
    .b(g72),
    .y(_00384_)
  );
  al_nand2ft _04995_ (
    .a(g72),
    .b(\DFF_1084.Q ),
    .y(_00385_)
  );
  al_and3 _04996_ (
    .a(_00384_),
    .b(_00385_),
    .c(_00383_),
    .y(_00386_)
  );
  al_inv _04997_ (
    .a(\DFF_1374.Q ),
    .y(_00387_)
  );
  al_and2 _04998_ (
    .a(\DFF_1379.Q ),
    .b(_00386_),
    .y(_00388_)
  );
  al_and3 _04999_ (
    .a(_00387_),
    .b(\DFF_1173.Q ),
    .c(_00388_),
    .y(_00389_)
  );
  al_and2 _05000_ (
    .a(\DFF_1347.Q ),
    .b(\DFF_443.Q ),
    .y(_00390_)
  );
  al_inv _05001_ (
    .a(\DFF_1379.Q ),
    .y(_00391_)
  );
  al_and2 _05002_ (
    .a(_00391_),
    .b(_00386_),
    .y(_00392_)
  );
  al_and2 _05003_ (
    .a(\DFF_1374.Q ),
    .b(\DFF_1173.Q ),
    .y(_00393_)
  );
  al_and2 _05004_ (
    .a(\DFF_118.Q ),
    .b(\DFF_139.Q ),
    .y(_00394_)
  );
  al_nand3 _05005_ (
    .a(_00393_),
    .b(_00394_),
    .c(_00392_),
    .y(_00395_)
  );
  al_ao21ttf _05006_ (
    .a(_00390_),
    .b(_00389_),
    .c(_00395_),
    .y(_00396_)
  );
  al_inv _05007_ (
    .a(\DFF_1173.Q ),
    .y(_00397_)
  );
  al_and3 _05008_ (
    .a(\DFF_1374.Q ),
    .b(_00397_),
    .c(_00392_),
    .y(_00398_)
  );
  al_and2 _05009_ (
    .a(\DFF_429.Q ),
    .b(\DFF_833.Q ),
    .y(_00399_)
  );
  al_nand2 _05010_ (
    .a(_00399_),
    .b(_00398_),
    .y(_00400_)
  );
  al_and3 _05011_ (
    .a(\DFF_1374.Q ),
    .b(_00397_),
    .c(_00388_),
    .y(_00401_)
  );
  al_and2 _05012_ (
    .a(\DFF_1312.Q ),
    .b(\DFF_536.Q ),
    .y(_00402_)
  );
  al_ao21ttf _05013_ (
    .a(_00401_),
    .b(_00402_),
    .c(_00400_),
    .y(_00403_)
  );
  al_and2 _05014_ (
    .a(\DFF_286.Q ),
    .b(\DFF_517.Q ),
    .y(_00404_)
  );
  al_nand3 _05015_ (
    .a(_00393_),
    .b(_00404_),
    .c(_00388_),
    .y(_00405_)
  );
  al_and3 _05016_ (
    .a(_00387_),
    .b(\DFF_1173.Q ),
    .c(_00392_),
    .y(_00406_)
  );
  al_nand2 _05017_ (
    .a(\DFF_1252.Q ),
    .b(\DFF_1283.Q ),
    .y(_00407_)
  );
  al_nand2ft _05018_ (
    .a(_00407_),
    .b(_00406_),
    .y(_00408_)
  );
  al_inv _05019_ (
    .a(g25114),
    .y(_00409_)
  );
  al_nor2 _05020_ (
    .a(\DFF_1374.Q ),
    .b(\DFF_1173.Q ),
    .y(_00410_)
  );
  al_and3 _05021_ (
    .a(\DFF_1379.Q ),
    .b(_00410_),
    .c(_00386_),
    .y(_00411_)
  );
  al_and2 _05022_ (
    .a(\DFF_952.Q ),
    .b(\DFF_878.Q ),
    .y(_00412_)
  );
  al_and2 _05023_ (
    .a(_00412_),
    .b(_00411_),
    .y(_00413_)
  );
  al_and3 _05024_ (
    .a(_00391_),
    .b(_00410_),
    .c(_00386_),
    .y(_00414_)
  );
  al_ao21ftt _05025_ (
    .a(_00409_),
    .b(_00414_),
    .c(_00413_),
    .y(_00415_)
  );
  al_nor3fft _05026_ (
    .a(_00405_),
    .b(_00408_),
    .c(_00415_),
    .y(_00416_)
  );
  al_nand3fft _05027_ (
    .a(_00396_),
    .b(_00403_),
    .c(_00416_),
    .y(\DFF_743.D )
  );
  al_or3fft _05028_ (
    .a(_00343_),
    .b(_00386_),
    .c(\DFF_743.D ),
    .y(g34425)
  );
  al_nor2 _05029_ (
    .a(\DFF_451.Q ),
    .b(g73),
    .y(_00417_)
  );
  al_nand2 _05030_ (
    .a(\DFF_451.Q ),
    .b(g73),
    .y(_00418_)
  );
  al_nand2ft _05031_ (
    .a(_00417_),
    .b(_00418_),
    .y(_00419_)
  );
  al_nand2ft _05032_ (
    .a(\DFF_951.Q ),
    .b(g72),
    .y(_00420_)
  );
  al_nand2ft _05033_ (
    .a(g72),
    .b(\DFF_951.Q ),
    .y(_00421_)
  );
  al_and3 _05034_ (
    .a(_00420_),
    .b(_00421_),
    .c(_00419_),
    .y(_00422_)
  );
  al_inv _05035_ (
    .a(\DFF_1020.Q ),
    .y(_00423_)
  );
  al_and2 _05036_ (
    .a(\DFF_428.Q ),
    .b(_00422_),
    .y(_00424_)
  );
  al_and3 _05037_ (
    .a(_00423_),
    .b(\DFF_1080.Q ),
    .c(_00424_),
    .y(_00425_)
  );
  al_and2ft _05038_ (
    .a(\DFF_681.Q ),
    .b(\DFF_297.Q ),
    .y(_00426_)
  );
  al_inv _05039_ (
    .a(\DFF_1080.Q ),
    .y(_00427_)
  );
  al_inv _05040_ (
    .a(\DFF_428.Q ),
    .y(_00428_)
  );
  al_and3 _05041_ (
    .a(\DFF_1020.Q ),
    .b(_00428_),
    .c(_00422_),
    .y(_00429_)
  );
  al_and2 _05042_ (
    .a(_00427_),
    .b(_00429_),
    .y(_00430_)
  );
  al_and2ft _05043_ (
    .a(\DFF_103.Q ),
    .b(\DFF_174.Q ),
    .y(_00431_)
  );
  al_inv _05044_ (
    .a(\DFF_1375.Q ),
    .y(_00432_)
  );
  al_and3fft _05045_ (
    .a(\DFF_1020.Q ),
    .b(\DFF_428.Q ),
    .c(\DFF_1080.Q ),
    .y(_00433_)
  );
  al_and2 _05046_ (
    .a(_00433_),
    .b(_00422_),
    .y(_00434_)
  );
  al_and3 _05047_ (
    .a(\DFF_1037.Q ),
    .b(_00432_),
    .c(_00434_),
    .y(_00435_)
  );
  al_aoi21 _05048_ (
    .a(_00431_),
    .b(_00430_),
    .c(_00435_),
    .y(_00436_)
  );
  al_ao21ttf _05049_ (
    .a(_00425_),
    .b(_00426_),
    .c(_00436_),
    .y(_00437_)
  );
  al_and2 _05050_ (
    .a(\DFF_1080.Q ),
    .b(_00429_),
    .y(_00438_)
  );
  al_and2ft _05051_ (
    .a(\DFF_1295.Q ),
    .b(\DFF_1236.Q ),
    .y(_00439_)
  );
  al_and3 _05052_ (
    .a(\DFF_1020.Q ),
    .b(_00427_),
    .c(_00424_),
    .y(_00440_)
  );
  al_and2ft _05053_ (
    .a(\DFF_148.Q ),
    .b(\DFF_793.Q ),
    .y(_00441_)
  );
  al_and2 _05054_ (
    .a(\DFF_1020.Q ),
    .b(\DFF_1080.Q ),
    .y(_00442_)
  );
  al_and3 _05055_ (
    .a(\DFF_428.Q ),
    .b(_00442_),
    .c(_00422_),
    .y(_00443_)
  );
  al_and2ft _05056_ (
    .a(\DFF_562.Q ),
    .b(\DFF_189.Q ),
    .y(_00444_)
  );
  al_and2 _05057_ (
    .a(_00444_),
    .b(_00443_),
    .y(_00445_)
  );
  al_aoi21 _05058_ (
    .a(_00441_),
    .b(_00440_),
    .c(_00445_),
    .y(_00446_)
  );
  al_ao21ttf _05059_ (
    .a(_00438_),
    .b(_00439_),
    .c(_00446_),
    .y(_00447_)
  );
  al_inv _05060_ (
    .a(\DFF_889.Q ),
    .y(_00448_)
  );
  al_and3 _05061_ (
    .a(_00423_),
    .b(_00427_),
    .c(_00424_),
    .y(_00449_)
  );
  al_nand3fft _05062_ (
    .a(\DFF_1091.Q ),
    .b(_00448_),
    .c(_00449_),
    .y(_00450_)
  );
  al_or3 _05063_ (
    .a(\DFF_1020.Q ),
    .b(\DFF_428.Q ),
    .c(\DFF_1080.Q ),
    .y(_00451_)
  );
  al_and2ft _05064_ (
    .a(_00451_),
    .b(_00422_),
    .y(_00452_)
  );
  al_aoi21ttf _05065_ (
    .a(g25167),
    .b(_00452_),
    .c(_00450_),
    .y(_00453_)
  );
  al_or3ftt _05066_ (
    .a(_00453_),
    .b(_00437_),
    .c(_00447_),
    .y(\DFF_379.D )
  );
  al_or3fft _05067_ (
    .a(_00343_),
    .b(_00422_),
    .c(\DFF_379.D ),
    .y(g34201)
  );
  al_nand3ftt _05068_ (
    .a(\DFF_934.Q ),
    .b(\DFF_1399.Q ),
    .c(_00342_),
    .y(g33874)
  );
  al_and2ft _05069_ (
    .a(g35),
    .b(\DFF_1314.Q ),
    .y(\DFF_800.D )
  );
  al_and3ftt _05070_ (
    .a(\DFF_894.Q ),
    .b(\DFF_849.Q ),
    .c(\DFF_207.Q ),
    .y(_00454_)
  );
  al_and2ft _05071_ (
    .a(\DFF_849.Q ),
    .b(\DFF_894.Q ),
    .y(_00455_)
  );
  al_and3 _05072_ (
    .a(\DFF_894.Q ),
    .b(\DFF_1006.Q ),
    .c(\DFF_849.Q ),
    .y(_00456_)
  );
  al_aoi21 _05073_ (
    .a(\DFF_609.Q ),
    .b(_00455_),
    .c(_00456_),
    .y(_00457_)
  );
  al_nand3fft _05074_ (
    .a(_00006_),
    .b(_00454_),
    .c(_00457_),
    .y(\DFF_417.D )
  );
  al_and2 _05075_ (
    .a(\DFF_1118.Q ),
    .b(_00342_),
    .y(_00458_)
  );
  al_or3fft _05076_ (
    .a(\DFF_997.Q ),
    .b(_00458_),
    .c(\DFF_417.D ),
    .y(g33636)
  );
  al_nand3 _05077_ (
    .a(\DFF_748.Q ),
    .b(_00238_),
    .c(_00223_),
    .y(g34927)
  );
  al_and2ft _05078_ (
    .a(g35),
    .b(\DFF_680.Q ),
    .y(\DFF_391.D )
  );
  al_and2ft _05079_ (
    .a(g35),
    .b(\DFF_445.Q ),
    .y(\DFF_680.D )
  );
  al_and3 _05080_ (
    .a(\DFF_635.Q ),
    .b(\DFF_270.Q ),
    .c(\DFF_1373.Q ),
    .y(_00459_)
  );
  al_and2 _05081_ (
    .a(\DFF_604.Q ),
    .b(_00459_),
    .y(_00460_)
  );
  al_and3ftt _05082_ (
    .a(\DFF_412.Q ),
    .b(\DFF_62.Q ),
    .c(\DFF_452.Q ),
    .y(_00461_)
  );
  al_and3 _05083_ (
    .a(\DFF_894.Q ),
    .b(\DFF_849.Q ),
    .c(_00461_),
    .y(_00462_)
  );
  al_nand3 _05084_ (
    .a(_00460_),
    .b(_00462_),
    .c(_00392_),
    .y(_00463_)
  );
  al_and3ftt _05085_ (
    .a(\DFF_847.Q ),
    .b(\DFF_914.Q ),
    .c(\DFF_218.Q ),
    .y(_00464_)
  );
  al_and3 _05086_ (
    .a(\DFF_1199.Q ),
    .b(\DFF_892.Q ),
    .c(_00464_),
    .y(_00465_)
  );
  al_and3 _05087_ (
    .a(\DFF_99.Q ),
    .b(\DFF_1326.Q ),
    .c(\DFF_1029.Q ),
    .y(_00466_)
  );
  al_nand3 _05088_ (
    .a(\DFF_1107.Q ),
    .b(_00466_),
    .c(_00465_),
    .y(_00467_)
  );
  al_ao21ftf _05089_ (
    .a(_00467_),
    .b(_00388_),
    .c(_00463_),
    .y(\DFF_796.D )
  );
  al_or3fft _05090_ (
    .a(_00343_),
    .b(_00386_),
    .c(\DFF_796.D ),
    .y(g34221)
  );
  al_nand2 _05091_ (
    .a(\DFF_748.Q ),
    .b(_00267_),
    .y(g34921)
  );
  al_and2ft _05092_ (
    .a(g35),
    .b(\DFF_932.Q ),
    .y(\DFF_1292.D )
  );
  al_nand3 _05093_ (
    .a(\DFF_748.Q ),
    .b(_00276_),
    .c(_00295_),
    .y(g34919)
  );
  al_and2ft _05094_ (
    .a(g35),
    .b(\DFF_1319.Q ),
    .y(\DFF_611.D )
  );
  al_nand2 _05095_ (
    .a(_00180_),
    .b(_00164_),
    .y(\DFF_355.D )
  );
  al_and3ftt _05096_ (
    .a(\DFF_892.Q ),
    .b(\DFF_1199.Q ),
    .c(\DFF_78.Q ),
    .y(_00468_)
  );
  al_and3fft _05097_ (
    .a(\DFF_1199.Q ),
    .b(\DFF_892.Q ),
    .c(\DFF_313.Q ),
    .y(_00469_)
  );
  al_and2ft _05098_ (
    .a(\DFF_1199.Q ),
    .b(\DFF_892.Q ),
    .y(_00470_)
  );
  al_and3 _05099_ (
    .a(\DFF_1199.Q ),
    .b(\DFF_922.Q ),
    .c(\DFF_892.Q ),
    .y(_00471_)
  );
  al_aoi21 _05100_ (
    .a(\DFF_684.Q ),
    .b(_00470_),
    .c(_00471_),
    .y(_00472_)
  );
  al_nand3fft _05101_ (
    .a(_00468_),
    .b(_00469_),
    .c(_00472_),
    .y(\DFF_1424.D )
  );
  al_and2 _05102_ (
    .a(\DFF_981.Q ),
    .b(_00342_),
    .y(_00473_)
  );
  al_or3fft _05103_ (
    .a(\DFF_1100.Q ),
    .b(_00473_),
    .c(\DFF_1424.D ),
    .y(g33935)
  );
  al_and2ft _05104_ (
    .a(g35),
    .b(\DFF_177.Q ),
    .y(\DFF_501.D )
  );
  al_and2ft _05105_ (
    .a(g35),
    .b(\DFF_399.Q ),
    .y(\DFF_1381.D )
  );
  al_inv _05106_ (
    .a(\DFF_582.Q ),
    .y(_00474_)
  );
  al_and3ftt _05107_ (
    .a(\DFF_447.Q ),
    .b(\DFF_591.Q ),
    .c(\DFF_96.Q ),
    .y(_00475_)
  );
  al_or3 _05108_ (
    .a(\DFF_1045.Q ),
    .b(\DFF_292.Q ),
    .c(\DFF_533.Q ),
    .y(_00476_)
  );
  al_and3 _05109_ (
    .a(\DFF_1393.Q ),
    .b(\DFF_798.Q ),
    .c(\DFF_1232.Q ),
    .y(_00477_)
  );
  al_and2ft _05110_ (
    .a(\DFF_1161.Q ),
    .b(_00477_),
    .y(_00478_)
  );
  al_or2 _05111_ (
    .a(\DFF_591.Q ),
    .b(\DFF_786.Q ),
    .y(_00479_)
  );
  al_or3 _05112_ (
    .a(\DFF_353.Q ),
    .b(\DFF_1145.Q ),
    .c(_00479_),
    .y(_00480_)
  );
  al_and3fft _05113_ (
    .a(\DFF_47.Q ),
    .b(_00480_),
    .c(_00478_),
    .y(_00481_)
  );
  al_nand2 _05114_ (
    .a(\DFF_142.Q ),
    .b(\DFF_21.Q ),
    .y(_00482_)
  );
  al_nand2 _05115_ (
    .a(\DFF_135.Q ),
    .b(\DFF_656.Q ),
    .y(_00483_)
  );
  al_oai21ttf _05116_ (
    .a(\DFF_135.Q ),
    .b(\DFF_656.Q ),
    .c(\DFF_194.Q ),
    .y(_00484_)
  );
  al_ao21ttf _05117_ (
    .a(\DFF_194.Q ),
    .b(_00483_),
    .c(_00484_),
    .y(_00485_)
  );
  al_nand3 _05118_ (
    .a(_00482_),
    .b(_00485_),
    .c(_00481_),
    .y(_00486_)
  );
  al_and2 _05119_ (
    .a(\DFF_1390.Q ),
    .b(_00486_),
    .y(_00487_)
  );
  al_aoi21ttf _05120_ (
    .a(_00475_),
    .b(_00476_),
    .c(_00487_),
    .y(_00488_)
  );
  al_nand2 _05121_ (
    .a(\DFF_1060.Q ),
    .b(_00475_),
    .y(_00489_)
  );
  al_nand3ftt _05122_ (
    .a(_00489_),
    .b(\DFF_1339.Q ),
    .c(_00488_),
    .y(_00490_)
  );
  al_and3fft _05123_ (
    .a(_00474_),
    .b(_00490_),
    .c(\DFF_409.Q ),
    .y(_00491_)
  );
  al_ao21 _05124_ (
    .a(\DFF_318.Q ),
    .b(_00491_),
    .c(\DFF_555.Q ),
    .y(_00492_)
  );
  al_and3 _05125_ (
    .a(\DFF_555.Q ),
    .b(\DFF_318.Q ),
    .c(_00488_),
    .y(_00493_)
  );
  al_nand2 _05126_ (
    .a(_00493_),
    .b(_00491_),
    .y(_00494_)
  );
  al_and2 _05127_ (
    .a(g35),
    .b(_00488_),
    .y(_00495_)
  );
  al_nand3 _05128_ (
    .a(_00495_),
    .b(_00494_),
    .c(_00492_),
    .y(_00496_)
  );
  al_ao21ftf _05129_ (
    .a(g35),
    .b(\DFF_318.Q ),
    .c(_00496_),
    .y(\DFF_555.D )
  );
  al_or3 _05130_ (
    .a(\DFF_244.Q ),
    .b(\DFF_958.Q ),
    .c(\DFF_289.Q ),
    .y(_00497_)
  );
  al_and2ft _05131_ (
    .a(\DFF_575.Q ),
    .b(\DFF_910.Q ),
    .y(_00498_)
  );
  al_and2ft _05132_ (
    .a(\DFF_1384.Q ),
    .b(\DFF_1389.Q ),
    .y(_00499_)
  );
  al_nand3ftt _05133_ (
    .a(_00497_),
    .b(_00498_),
    .c(_00499_),
    .y(_00500_)
  );
  al_ao21ftt _05134_ (
    .a(_00497_),
    .b(_00498_),
    .c(\DFF_938.Q ),
    .y(_00501_)
  );
  al_nand3 _05135_ (
    .a(g35),
    .b(_00500_),
    .c(_00501_),
    .y(_00502_)
  );
  al_ao21ftf _05136_ (
    .a(g35),
    .b(\DFF_307.Q ),
    .c(_00502_),
    .y(\DFF_938.D )
  );
  al_and3ftt _05137_ (
    .a(\DFF_880.Q ),
    .b(\DFF_339.Q ),
    .c(g35),
    .y(\DFF_880.D )
  );
  al_inv _05138_ (
    .a(\DFF_980.Q ),
    .y(_00503_)
  );
  al_or3 _05139_ (
    .a(\DFF_613.Q ),
    .b(\DFF_234.Q ),
    .c(\DFF_159.Q ),
    .y(_00504_)
  );
  al_or3 _05140_ (
    .a(\DFF_1002.Q ),
    .b(\DFF_1073.Q ),
    .c(_00504_),
    .y(_00505_)
  );
  al_nand2ft _05141_ (
    .a(\DFF_250.Q ),
    .b(\DFF_159.Q ),
    .y(_00506_)
  );
  al_oai21ftt _05142_ (
    .a(_00503_),
    .b(_00505_),
    .c(_00506_),
    .y(_00507_)
  );
  al_mux2h _05143_ (
    .a(\DFF_613.Q ),
    .b(_00507_),
    .s(g35),
    .y(\DFF_1073.D )
  );
  al_and2ft _05144_ (
    .a(\DFF_410.Q ),
    .b(\DFF_584.Q ),
    .y(_00508_)
  );
  al_nor2 _05145_ (
    .a(\DFF_1150.Q ),
    .b(\DFF_1068.Q ),
    .y(_00509_)
  );
  al_nand3 _05146_ (
    .a(_00499_),
    .b(_00508_),
    .c(_00509_),
    .y(_00510_)
  );
  al_ao21 _05147_ (
    .a(_00508_),
    .b(_00509_),
    .c(\DFF_419.Q ),
    .y(_00511_)
  );
  al_nand3 _05148_ (
    .a(g35),
    .b(_00511_),
    .c(_00510_),
    .y(_00512_)
  );
  al_ao21ftf _05149_ (
    .a(g35),
    .b(\DFF_957.Q ),
    .c(_00512_),
    .y(\DFF_419.D )
  );
  al_inv _05150_ (
    .a(\DFF_1233.Q ),
    .y(_00513_)
  );
  al_inv _05151_ (
    .a(\DFF_209.Q ),
    .y(_00514_)
  );
  al_and2ft _05152_ (
    .a(\DFF_956.Q ),
    .b(\DFF_1390.Q ),
    .y(_00515_)
  );
  al_oa21 _05153_ (
    .a(\DFF_1039.Q ),
    .b(\DFF_1343.Q ),
    .c(\DFF_1159.Q ),
    .y(_00516_)
  );
  al_ao21 _05154_ (
    .a(_00515_),
    .b(_00516_),
    .c(g134),
    .y(_00517_)
  );
  al_aoi21ftf _05155_ (
    .a(\DFF_948.Q ),
    .b(\DFF_403.Q ),
    .c(_00517_),
    .y(_00518_)
  );
  al_nand3ftt _05156_ (
    .a(\DFF_1270.Q ),
    .b(\DFF_1319.Q ),
    .c(\DFF_1067.Q ),
    .y(_00519_)
  );
  al_inv _05157_ (
    .a(\DFF_146.Q ),
    .y(_00520_)
  );
  al_and2ft _05158_ (
    .a(\DFF_1148.Q ),
    .b(\DFF_717.Q ),
    .y(_00521_)
  );
  al_nor2 _05159_ (
    .a(\DFF_1194.Q ),
    .b(\DFF_1313.Q ),
    .y(_00522_)
  );
  al_and3ftt _05160_ (
    .a(\DFF_1371.Q ),
    .b(\DFF_740.Q ),
    .c(\DFF_990.Q ),
    .y(_00523_)
  );
  al_and3ftt _05161_ (
    .a(\DFF_375.Q ),
    .b(_00523_),
    .c(_00522_),
    .y(_00524_)
  );
  al_ao21 _05162_ (
    .a(_00521_),
    .b(_00524_),
    .c(_00520_),
    .y(_00525_)
  );
  al_nand3 _05163_ (
    .a(_00519_),
    .b(_00518_),
    .c(_00525_),
    .y(_00526_)
  );
  al_nand3fft _05164_ (
    .a(_00513_),
    .b(_00514_),
    .c(_00526_),
    .y(_00527_)
  );
  al_inv _05165_ (
    .a(\DFF_1389.Q ),
    .y(_00528_)
  );
  al_aoi21ftf _05166_ (
    .a(_00519_),
    .b(_00528_),
    .c(_00518_),
    .y(_00529_)
  );
  al_aoi21ftf _05167_ (
    .a(\DFF_481.Q ),
    .b(_00519_),
    .c(_00529_),
    .y(_00530_)
  );
  al_aoi21ftf _05168_ (
    .a(\DFF_457.Q ),
    .b(_00527_),
    .c(g35),
    .y(_00531_)
  );
  al_ao21ftf _05169_ (
    .a(_00527_),
    .b(_00530_),
    .c(_00531_),
    .y(_00532_)
  );
  al_ao21ftf _05170_ (
    .a(g35),
    .b(\DFF_625.Q ),
    .c(_00532_),
    .y(\DFF_457.D )
  );
  al_and3 _05171_ (
    .a(\DFF_871.Q ),
    .b(\DFF_1275.Q ),
    .c(\DFF_1017.Q ),
    .y(_00533_)
  );
  al_and3 _05172_ (
    .a(\DFF_901.Q ),
    .b(\DFF_1117.Q ),
    .c(_00533_),
    .y(_00534_)
  );
  al_nand2 _05173_ (
    .a(\DFF_1275.Q ),
    .b(\DFF_431.Q ),
    .y(_00535_)
  );
  al_nand2 _05174_ (
    .a(\DFF_431.Q ),
    .b(_00534_),
    .y(_00536_)
  );
  al_aoi21ftf _05175_ (
    .a(_00534_),
    .b(_00535_),
    .c(_00536_),
    .y(_00537_)
  );
  al_mux2h _05176_ (
    .a(\DFF_901.Q ),
    .b(_00537_),
    .s(g35),
    .y(\DFF_431.D )
  );
  al_mux2l _05177_ (
    .a(\DFF_382.Q ),
    .b(\DFF_496.Q ),
    .s(g72),
    .y(_00538_)
  );
  al_mux2l _05178_ (
    .a(\DFF_362.Q ),
    .b(\DFF_346.Q ),
    .s(g72),
    .y(_00539_)
  );
  al_mux2l _05179_ (
    .a(_00538_),
    .b(_00539_),
    .s(g73),
    .y(_00540_)
  );
  al_mux2h _05180_ (
    .a(\DFF_252.Q ),
    .b(_00540_),
    .s(g35),
    .y(\DFF_357.D )
  );
  al_and2 _05181_ (
    .a(\DFF_199.Q ),
    .b(g35),
    .y(\DFF_830.D )
  );
  al_inv _05182_ (
    .a(\DFF_552.Q ),
    .y(_00541_)
  );
  al_nor2 _05183_ (
    .a(\DFF_845.Q ),
    .b(\DFF_746.Q ),
    .y(_00542_)
  );
  al_inv _05184_ (
    .a(_00542_),
    .y(_00543_)
  );
  al_oai21ftt _05185_ (
    .a(\DFF_1364.Q ),
    .b(_00451_),
    .c(_00542_),
    .y(_00544_)
  );
  al_and3ftt _05186_ (
    .a(\DFF_893.Q ),
    .b(\DFF_962.Q ),
    .c(_00544_),
    .y(_00545_)
  );
  al_aoi21ftf _05187_ (
    .a(_00543_),
    .b(\DFF_1288.Q ),
    .c(_00545_),
    .y(_00546_)
  );
  al_nand3fft _05188_ (
    .a(_00432_),
    .b(_00541_),
    .c(_00546_),
    .y(_00547_)
  );
  al_nand2 _05189_ (
    .a(g35),
    .b(_00547_),
    .y(_00548_)
  );
  al_mux2l _05190_ (
    .a(\DFF_1075.Q ),
    .b(\DFF_882.Q ),
    .s(_00548_),
    .y(\DFF_882.D )
  );
  al_and2 _05191_ (
    .a(\DFF_498.Q ),
    .b(g35),
    .y(\DFF_498.D )
  );
  al_and3 _05192_ (
    .a(\DFF_1364.Q ),
    .b(\DFF_428.Q ),
    .c(_00442_),
    .y(_00549_)
  );
  al_aoi21ftt _05193_ (
    .a(\DFF_1020.Q ),
    .b(_00428_),
    .c(_00549_),
    .y(_00550_)
  );
  al_ao21ftt _05194_ (
    .a(\DFF_1240.Q ),
    .b(_00550_),
    .c(\DFF_470.Q ),
    .y(_00551_)
  );
  al_nor2ft _05195_ (
    .a(g35),
    .b(_00433_),
    .y(_00552_)
  );
  al_and2ft _05196_ (
    .a(g35),
    .b(\DFF_763.Q ),
    .y(_00553_)
  );
  al_ao21 _05197_ (
    .a(_00552_),
    .b(_00551_),
    .c(_00553_),
    .y(\DFF_470.D )
  );
  al_aoi21 _05198_ (
    .a(\DFF_68.Q ),
    .b(g35),
    .c(\DFF_1098.Q ),
    .y(_00554_)
  );
  al_inv _05199_ (
    .a(\DFF_1098.Q ),
    .y(_00555_)
  );
  al_and3ftt _05200_ (
    .a(g113),
    .b(\DFF_304.Q ),
    .c(_00342_),
    .y(_00556_)
  );
  al_nand3ftt _05201_ (
    .a(_00306_),
    .b(_00556_),
    .c(_00354_),
    .y(_00557_)
  );
  al_ao21ftf _05202_ (
    .a(_00555_),
    .b(\DFF_68.Q ),
    .c(_00557_),
    .y(_00558_)
  );
  al_aoi21 _05203_ (
    .a(g35),
    .b(_00558_),
    .c(_00554_),
    .y(\DFF_68.D )
  );
  al_inv _05204_ (
    .a(\DFF_1331.Q ),
    .y(_00559_)
  );
  al_inv _05205_ (
    .a(\DFF_148.Q ),
    .y(_00560_)
  );
  al_and2ft _05206_ (
    .a(\DFF_962.Q ),
    .b(\DFF_893.Q ),
    .y(_00561_)
  );
  al_and2 _05207_ (
    .a(_00561_),
    .b(_00544_),
    .y(_00562_)
  );
  al_aoi21ftf _05208_ (
    .a(_00543_),
    .b(\DFF_302.Q ),
    .c(_00562_),
    .y(_00563_)
  );
  al_nand3fft _05209_ (
    .a(_00559_),
    .b(_00560_),
    .c(_00563_),
    .y(_00564_)
  );
  al_aoi21 _05210_ (
    .a(\DFF_1395.Q ),
    .b(_00564_),
    .c(_00066_),
    .y(_00565_)
  );
  al_oai21 _05211_ (
    .a(\DFF_1395.Q ),
    .b(_00564_),
    .c(_00565_),
    .y(_00566_)
  );
  al_aoi21ftf _05212_ (
    .a(\DFF_818.Q ),
    .b(_00066_),
    .c(_00566_),
    .y(\DFF_1395.D )
  );
  al_and2 _05213_ (
    .a(\DFF_1304.Q ),
    .b(\DFF_407.Q ),
    .y(_00567_)
  );
  al_nand3 _05214_ (
    .a(_00555_),
    .b(_00567_),
    .c(_00557_),
    .y(_00568_)
  );
  al_ao21ftf _05215_ (
    .a(g35),
    .b(\DFF_1304.Q ),
    .c(_00568_),
    .y(\DFF_1098.D )
  );
  al_oa21ftt _05216_ (
    .a(g35),
    .b(\DFF_605.Q ),
    .c(\DFF_285.Q ),
    .y(_00569_)
  );
  al_nand2ft _05217_ (
    .a(\DFF_1367.Q ),
    .b(\DFF_668.Q ),
    .y(_00570_)
  );
  al_oa21ftf _05218_ (
    .a(\DFF_668.Q ),
    .b(\DFF_787.Q ),
    .c(\DFF_605.Q ),
    .y(_00571_)
  );
  al_ao21ftf _05219_ (
    .a(\DFF_285.Q ),
    .b(_00571_),
    .c(_00570_),
    .y(_00572_)
  );
  al_ao21 _05220_ (
    .a(g35),
    .b(_00572_),
    .c(_00569_),
    .y(\DFF_605.D )
  );
  al_or2 _05221_ (
    .a(_00066_),
    .b(_00481_),
    .y(_00573_)
  );
  al_mux2l _05222_ (
    .a(\DFF_988.Q ),
    .b(\DFF_194.Q ),
    .s(_00573_),
    .y(\DFF_194.D )
  );
  al_mux2l _05223_ (
    .a(g6748),
    .b(\DFF_1209.Q ),
    .s(g35),
    .y(\DFF_383.D )
  );
  al_nand3fft _05224_ (
    .a(\DFF_1131.Q ),
    .b(\DFF_416.Q ),
    .c(g35),
    .y(g28042)
  );
  al_inv _05225_ (
    .a(\DFF_993.Q ),
    .y(_00574_)
  );
  al_nor2 _05226_ (
    .a(\DFF_893.Q ),
    .b(\DFF_962.Q ),
    .y(_00575_)
  );
  al_and3 _05227_ (
    .a(_00002_),
    .b(_00575_),
    .c(_00544_),
    .y(_00576_)
  );
  al_and3ftt _05228_ (
    .a(g113),
    .b(\DFF_379.Q ),
    .c(_00342_),
    .y(_00577_)
  );
  al_aoi21ttf _05229_ (
    .a(_00577_),
    .b(_00449_),
    .c(_00576_),
    .y(_00578_)
  );
  al_or2 _05230_ (
    .a(_00066_),
    .b(_00578_),
    .y(_00579_)
  );
  al_and3fft _05231_ (
    .a(_00066_),
    .b(_00576_),
    .c(_00448_),
    .y(_00580_)
  );
  al_aoi21 _05232_ (
    .a(_00574_),
    .b(_00579_),
    .c(_00580_),
    .y(\DFF_889.D )
  );
  al_and2ft _05233_ (
    .a(g35),
    .b(\DFF_347.Q ),
    .y(_00581_)
  );
  al_nand2 _05234_ (
    .a(\DFF_1326.Q ),
    .b(\DFF_1029.Q ),
    .y(_00582_)
  );
  al_and3fft _05235_ (
    .a(\DFF_847.Q ),
    .b(\DFF_218.Q ),
    .c(\DFF_914.Q ),
    .y(_00583_)
  );
  al_nor3fft _05236_ (
    .a(\DFF_1107.Q ),
    .b(_00583_),
    .c(_00582_),
    .y(_00584_)
  );
  al_aoi21ttf _05237_ (
    .a(_00471_),
    .b(_00584_),
    .c(\DFF_99.Q ),
    .y(_00585_)
  );
  al_and3 _05238_ (
    .a(\DFF_1379.Q ),
    .b(_00393_),
    .c(_00386_),
    .y(_00586_)
  );
  al_and3ftt _05239_ (
    .a(g113),
    .b(\DFF_743.Q ),
    .c(_00342_),
    .y(_00587_)
  );
  al_nand3 _05240_ (
    .a(_00585_),
    .b(_00587_),
    .c(_00586_),
    .y(_00588_)
  );
  al_ao21 _05241_ (
    .a(_00585_),
    .b(_00588_),
    .c(\DFF_286.Q ),
    .y(_00589_)
  );
  al_aoi21 _05242_ (
    .a(\DFF_286.Q ),
    .b(_00585_),
    .c(_00066_),
    .y(_00590_)
  );
  al_ao21 _05243_ (
    .a(_00590_),
    .b(_00589_),
    .c(_00581_),
    .y(\DFF_286.D )
  );
  al_and2 _05244_ (
    .a(\DFF_519.Q ),
    .b(\DFF_385.Q ),
    .y(_00591_)
  );
  al_and2ft _05245_ (
    .a(\DFF_734.Q ),
    .b(\DFF_723.Q ),
    .y(_00592_)
  );
  al_nand3 _05246_ (
    .a(_00499_),
    .b(_00591_),
    .c(_00592_),
    .y(_00593_)
  );
  al_ao21 _05247_ (
    .a(_00592_),
    .b(_00591_),
    .c(\DFF_949.Q ),
    .y(_00594_)
  );
  al_nand3 _05248_ (
    .a(g35),
    .b(_00594_),
    .c(_00593_),
    .y(_00595_)
  );
  al_ao21ftf _05249_ (
    .a(g35),
    .b(\DFF_854.Q ),
    .c(_00595_),
    .y(\DFF_949.D )
  );
  al_and2 _05250_ (
    .a(\DFF_784.Q ),
    .b(\DFF_776.Q ),
    .y(_00596_)
  );
  al_and2ft _05251_ (
    .a(\DFF_587.Q ),
    .b(\DFF_467.Q ),
    .y(_00597_)
  );
  al_nand3 _05252_ (
    .a(_00499_),
    .b(_00596_),
    .c(_00597_),
    .y(_00598_)
  );
  al_ao21 _05253_ (
    .a(_00597_),
    .b(_00596_),
    .c(\DFF_1317.Q ),
    .y(_00599_)
  );
  al_nand3 _05254_ (
    .a(g35),
    .b(_00599_),
    .c(_00598_),
    .y(_00600_)
  );
  al_ao21ftf _05255_ (
    .a(g35),
    .b(\DFF_868.Q ),
    .c(_00600_),
    .y(\DFF_1317.D )
  );
  al_and3ftt _05256_ (
    .a(\DFF_331.Q ),
    .b(\DFF_43.Q ),
    .c(\DFF_1412.Q ),
    .y(_00601_)
  );
  al_and3 _05257_ (
    .a(\DFF_853.Q ),
    .b(_00601_),
    .c(_00393_),
    .y(_00602_)
  );
  al_and3 _05258_ (
    .a(\DFF_115.Q ),
    .b(\DFF_1084.Q ),
    .c(_00602_),
    .y(_00603_)
  );
  al_and2ft _05259_ (
    .a(g113),
    .b(_00342_),
    .y(_00604_)
  );
  al_nor2 _05260_ (
    .a(g73),
    .b(g72),
    .y(_00605_)
  );
  al_oai21ftt _05261_ (
    .a(_00605_),
    .b(_00604_),
    .c(\DFF_961.Q ),
    .y(_00606_)
  );
  al_nor3fft _05262_ (
    .a(g35),
    .b(_00606_),
    .c(_00603_),
    .y(_00607_)
  );
  al_nand3 _05263_ (
    .a(\DFF_1374.Q ),
    .b(\DFF_1173.Q ),
    .c(\DFF_853.Q ),
    .y(_00608_)
  );
  al_nor3fft _05264_ (
    .a(\DFF_1379.Q ),
    .b(_00601_),
    .c(_00608_),
    .y(_00609_)
  );
  al_oai21ftf _05265_ (
    .a(_00601_),
    .b(_00608_),
    .c(\DFF_1379.Q ),
    .y(_00610_)
  );
  al_and3ftt _05266_ (
    .a(_00609_),
    .b(_00610_),
    .c(_00607_),
    .y(\DFF_1379.D )
  );
  al_ao21ttf _05267_ (
    .a(\DFF_775.Q ),
    .b(\DFF_827.Q ),
    .c(g35),
    .y(_00611_)
  );
  al_and2 _05268_ (
    .a(\DFF_1156.Q ),
    .b(_00611_),
    .y(_00612_)
  );
  al_or3fft _05269_ (
    .a(\DFF_1076.Q ),
    .b(g35),
    .c(_00612_),
    .y(_00613_)
  );
  al_aoi21ftf _05270_ (
    .a(_00066_),
    .b(\DFF_1076.Q ),
    .c(_00612_),
    .y(_00614_)
  );
  al_nand2ft _05271_ (
    .a(_00614_),
    .b(_00613_),
    .y(\DFF_1076.D )
  );
  al_mux2l _05272_ (
    .a(\DFF_339.Q ),
    .b(\DFF_791.Q ),
    .s(g35),
    .y(\DFF_606.D )
  );
  al_nor2 _05273_ (
    .a(\DFF_456.Q ),
    .b(\DFF_1284.Q ),
    .y(_00615_)
  );
  al_or2 _05274_ (
    .a(\DFF_441.Q ),
    .b(\DFF_1260.Q ),
    .y(_00616_)
  );
  al_nor2 _05275_ (
    .a(\DFF_222.Q ),
    .b(\DFF_1302.Q ),
    .y(_00617_)
  );
  al_or2 _05276_ (
    .a(\DFF_243.Q ),
    .b(\DFF_778.Q ),
    .y(_00618_)
  );
  al_and3fft _05277_ (
    .a(_00616_),
    .b(_00618_),
    .c(_00617_),
    .y(_00619_)
  );
  al_aoi21 _05278_ (
    .a(_00615_),
    .b(_00619_),
    .c(_00066_),
    .y(_00620_)
  );
  al_nor2 _05279_ (
    .a(\DFF_287.Q ),
    .b(\DFF_52.Q ),
    .y(_00621_)
  );
  al_or2 _05280_ (
    .a(\DFF_1079.Q ),
    .b(\DFF_310.Q ),
    .y(_00622_)
  );
  al_oa21 _05281_ (
    .a(\DFF_361.Q ),
    .b(\DFF_1198.Q ),
    .c(g35),
    .y(_00623_)
  );
  al_aoi21 _05282_ (
    .a(g35),
    .b(_00622_),
    .c(_00623_),
    .y(_00624_)
  );
  al_oai21 _05283_ (
    .a(\DFF_1079.Q ),
    .b(\DFF_310.Q ),
    .c(_00623_),
    .y(_00625_)
  );
  al_ao21 _05284_ (
    .a(_00621_),
    .b(_00625_),
    .c(_00624_),
    .y(_00626_)
  );
  al_ao21ftf _05285_ (
    .a(_00621_),
    .b(g35),
    .c(_00624_),
    .y(_00627_)
  );
  al_oai21 _05286_ (
    .a(\DFF_332.Q ),
    .b(\DFF_716.Q ),
    .c(g35),
    .y(_00628_)
  );
  al_aoi21ftf _05287_ (
    .a(_00628_),
    .b(_00627_),
    .c(_00626_),
    .y(_00629_)
  );
  al_nand3fft _05288_ (
    .a(\DFF_243.Q ),
    .b(\DFF_778.Q ),
    .c(_00617_),
    .y(_00630_)
  );
  al_oai21ftf _05289_ (
    .a(_00618_),
    .b(_00617_),
    .c(_00616_),
    .y(_00631_)
  );
  al_nand3 _05290_ (
    .a(g35),
    .b(_00630_),
    .c(_00631_),
    .y(_00632_)
  );
  al_mux2h _05291_ (
    .a(_00619_),
    .b(_00632_),
    .s(_00615_),
    .y(_00633_)
  );
  al_or2ft _05292_ (
    .a(_00628_),
    .b(_00627_),
    .y(_00634_)
  );
  al_or3fft _05293_ (
    .a(_00620_),
    .b(_00633_),
    .c(_00634_),
    .y(_00635_)
  );
  al_ao21ftf _05294_ (
    .a(_00620_),
    .b(_00629_),
    .c(_00635_),
    .y(g28030)
  );
  al_inv _05295_ (
    .a(\DFF_1323.Q ),
    .y(_00636_)
  );
  al_aoi21ftf _05296_ (
    .a(_00636_),
    .b(_00081_),
    .c(_00517_),
    .y(_00637_)
  );
  al_nand3 _05297_ (
    .a(\DFF_1270.Q ),
    .b(\DFF_1319.Q ),
    .c(\DFF_1067.Q ),
    .y(_00638_)
  );
  al_nor2 _05298_ (
    .a(\DFF_1148.Q ),
    .b(\DFF_717.Q ),
    .y(_00639_)
  );
  al_ao21ttf _05299_ (
    .a(_00639_),
    .b(_00524_),
    .c(\DFF_372.Q ),
    .y(_00640_)
  );
  al_nand3 _05300_ (
    .a(_00638_),
    .b(_00637_),
    .c(_00640_),
    .y(_00641_)
  );
  al_nand3fft _05301_ (
    .a(\DFF_713.Q ),
    .b(\DFF_505.Q ),
    .c(_00641_),
    .y(_00642_)
  );
  al_nor2 _05302_ (
    .a(\DFF_1368.Q ),
    .b(\DFF_702.Q ),
    .y(_00643_)
  );
  al_nand2 _05303_ (
    .a(\DFF_1368.Q ),
    .b(\DFF_702.Q ),
    .y(_00644_)
  );
  al_nand2ft _05304_ (
    .a(_00643_),
    .b(_00644_),
    .y(_00645_)
  );
  al_mux2l _05305_ (
    .a(\DFF_1071.Q ),
    .b(_00645_),
    .s(_00642_),
    .y(_00646_)
  );
  al_mux2h _05306_ (
    .a(\DFF_702.Q ),
    .b(_00646_),
    .s(g35),
    .y(\DFF_1071.D )
  );
  al_nor2 _05307_ (
    .a(g35),
    .b(\DFF_1363.Q ),
    .y(_00647_)
  );
  al_nand3 _05308_ (
    .a(\DFF_659.Q ),
    .b(\DFF_360.Q ),
    .c(g25114),
    .y(_00648_)
  );
  al_nand2ft _05309_ (
    .a(\DFF_846.Q ),
    .b(\DFF_449.Q ),
    .y(_00649_)
  );
  al_or3fft _05310_ (
    .a(\DFF_773.Q ),
    .b(\DFF_537.Q ),
    .c(_00649_),
    .y(_00650_)
  );
  al_and3 _05311_ (
    .a(\DFF_141.Q ),
    .b(_00650_),
    .c(_00648_),
    .y(_00651_)
  );
  al_or2 _05312_ (
    .a(\DFF_449.Q ),
    .b(\DFF_846.Q ),
    .y(_00652_)
  );
  al_nand2 _05313_ (
    .a(\DFF_638.Q ),
    .b(\DFF_616.Q ),
    .y(_00653_)
  );
  al_nand2 _05314_ (
    .a(\DFF_100.Q ),
    .b(\DFF_281.Q ),
    .y(_00654_)
  );
  al_ao21 _05315_ (
    .a(_00653_),
    .b(_00654_),
    .c(_00652_),
    .y(_00655_)
  );
  al_nand2ft _05316_ (
    .a(\DFF_449.Q ),
    .b(\DFF_846.Q ),
    .y(_00656_)
  );
  al_nand2 _05317_ (
    .a(\DFF_923.Q ),
    .b(\DFF_765.Q ),
    .y(_00657_)
  );
  al_nand2 _05318_ (
    .a(\DFF_165.Q ),
    .b(\DFF_1325.Q ),
    .y(_00658_)
  );
  al_ao21 _05319_ (
    .a(_00657_),
    .b(_00658_),
    .c(_00656_),
    .y(_00659_)
  );
  al_nand3 _05320_ (
    .a(_00655_),
    .b(_00659_),
    .c(_00651_),
    .y(_00660_)
  );
  al_nand2 _05321_ (
    .a(\DFF_566.Q ),
    .b(\DFF_1040.Q ),
    .y(_00661_)
  );
  al_nand2 _05322_ (
    .a(\DFF_187.Q ),
    .b(\DFF_360.Q ),
    .y(_00662_)
  );
  al_ao21 _05323_ (
    .a(_00661_),
    .b(_00662_),
    .c(_00656_),
    .y(_00663_)
  );
  al_nand2 _05324_ (
    .a(\DFF_750.Q ),
    .b(\DFF_281.Q ),
    .y(_00664_)
  );
  al_ao21ttf _05325_ (
    .a(\DFF_390.Q ),
    .b(\DFF_616.Q ),
    .c(_00664_),
    .y(_00665_)
  );
  al_aoi21ftf _05326_ (
    .a(_00649_),
    .b(_00665_),
    .c(_00663_),
    .y(_00666_)
  );
  al_nor3fft _05327_ (
    .a(\DFF_1212.Q ),
    .b(\DFF_537.Q ),
    .c(_00652_),
    .y(_00667_)
  );
  al_nand2 _05328_ (
    .a(\DFF_165.Q ),
    .b(\DFF_602.Q ),
    .y(_00668_)
  );
  al_nand2 _05329_ (
    .a(\DFF_13.Q ),
    .b(\DFF_765.Q ),
    .y(_00669_)
  );
  al_ao21ttf _05330_ (
    .a(_00668_),
    .b(_00669_),
    .c(g25114),
    .y(_00670_)
  );
  al_nand3fft _05331_ (
    .a(\DFF_141.Q ),
    .b(_00667_),
    .c(_00670_),
    .y(_00671_)
  );
  al_ao21ftf _05332_ (
    .a(_00671_),
    .b(_00666_),
    .c(_00660_),
    .y(_00672_)
  );
  al_and3 _05333_ (
    .a(\DFF_566.Q ),
    .b(\DFF_141.Q ),
    .c(g25114),
    .y(_00673_)
  );
  al_nand2 _05334_ (
    .a(\DFF_1363.Q ),
    .b(_00673_),
    .y(_00674_)
  );
  al_or3fft _05335_ (
    .a(\DFF_906.Q ),
    .b(\DFF_497.Q ),
    .c(_00649_),
    .y(_00675_)
  );
  al_nor2 _05336_ (
    .a(\DFF_141.Q ),
    .b(\DFF_165.Q ),
    .y(_00676_)
  );
  al_nand2 _05337_ (
    .a(\DFF_141.Q ),
    .b(\DFF_165.Q ),
    .y(_00677_)
  );
  al_and3ftt _05338_ (
    .a(_00676_),
    .b(_00677_),
    .c(_00675_),
    .y(_00678_)
  );
  al_or3fft _05339_ (
    .a(\DFF_927.Q ),
    .b(\DFF_1095.Q ),
    .c(_00656_),
    .y(_00679_)
  );
  al_or3fft _05340_ (
    .a(\DFF_655.Q ),
    .b(\DFF_983.Q ),
    .c(_00652_),
    .y(_00680_)
  );
  al_nand3 _05341_ (
    .a(_00679_),
    .b(_00680_),
    .c(_00678_),
    .y(_00681_)
  );
  al_and2 _05342_ (
    .a(\DFF_906.Q ),
    .b(\DFF_1406.Q ),
    .y(_00682_)
  );
  al_or3fft _05343_ (
    .a(\DFF_655.Q ),
    .b(\DFF_1186.Q ),
    .c(_00649_),
    .y(_00683_)
  );
  al_aoi21ftf _05344_ (
    .a(_00652_),
    .b(_00682_),
    .c(_00683_),
    .y(_00684_)
  );
  al_nand3 _05345_ (
    .a(\DFF_927.Q ),
    .b(\DFF_950.Q ),
    .c(g25114),
    .y(_00685_)
  );
  al_ao21ftf _05346_ (
    .a(_00676_),
    .b(_00677_),
    .c(_00685_),
    .y(_00686_)
  );
  al_ao21ftf _05347_ (
    .a(_00686_),
    .b(_00684_),
    .c(_00681_),
    .y(_00687_)
  );
  al_nand3 _05348_ (
    .a(_00674_),
    .b(_00687_),
    .c(_00672_),
    .y(_00688_)
  );
  al_nand2 _05349_ (
    .a(g28753),
    .b(_00688_),
    .y(_00689_)
  );
  al_oa21ftf _05350_ (
    .a(\DFF_132.Q ),
    .b(g28753),
    .c(_00066_),
    .y(_00690_)
  );
  al_aoi21 _05351_ (
    .a(_00690_),
    .b(_00689_),
    .c(_00647_),
    .y(\DFF_132.D )
  );
  al_nor2 _05352_ (
    .a(\DFF_587.Q ),
    .b(\DFF_467.Q ),
    .y(_00691_)
  );
  al_nand3 _05353_ (
    .a(_00499_),
    .b(_00596_),
    .c(_00691_),
    .y(_00692_)
  );
  al_ao21 _05354_ (
    .a(_00691_),
    .b(_00596_),
    .c(\DFF_947.Q ),
    .y(_00693_)
  );
  al_nand3 _05355_ (
    .a(g35),
    .b(_00693_),
    .c(_00692_),
    .y(_00694_)
  );
  al_ao21ftf _05356_ (
    .a(g35),
    .b(\DFF_257.Q ),
    .c(_00694_),
    .y(\DFF_947.D )
  );
  al_inv _05357_ (
    .a(\DFF_845.Q ),
    .y(_00695_)
  );
  al_inv _05358_ (
    .a(\DFF_746.Q ),
    .y(_00696_)
  );
  al_nand3fft _05359_ (
    .a(_00695_),
    .b(_00696_),
    .c(_00549_),
    .y(_00697_)
  );
  al_and3ftt _05360_ (
    .a(g113),
    .b(\DFF_1220.Q ),
    .c(_00342_),
    .y(_00698_)
  );
  al_oa21ftf _05361_ (
    .a(\DFF_1104.Q ),
    .b(_00604_),
    .c(_00698_),
    .y(_00699_)
  );
  al_mux2l _05362_ (
    .a(\DFF_233.Q ),
    .b(_00699_),
    .s(_00697_),
    .y(_00700_)
  );
  al_mux2h _05363_ (
    .a(\DFF_1104.Q ),
    .b(_00700_),
    .s(g35),
    .y(\DFF_233.D )
  );
  al_or3 _05364_ (
    .a(\DFF_734.Q ),
    .b(\DFF_723.Q ),
    .c(\DFF_393.Q ),
    .y(_00701_)
  );
  al_nand3ftt _05365_ (
    .a(_00701_),
    .b(_00591_),
    .c(_00499_),
    .y(_00702_)
  );
  al_ao21ftt _05366_ (
    .a(_00701_),
    .b(_00591_),
    .c(\DFF_17.Q ),
    .y(_00703_)
  );
  al_nand3 _05367_ (
    .a(g35),
    .b(_00702_),
    .c(_00703_),
    .y(_00704_)
  );
  al_ao21ftf _05368_ (
    .a(g35),
    .b(\DFF_1201.Q ),
    .c(_00704_),
    .y(\DFF_17.D )
  );
  al_and2ft _05369_ (
    .a(\DFF_35.Q ),
    .b(\DFF_803.Q ),
    .y(_00705_)
  );
  al_and2ft _05370_ (
    .a(\DFF_522.Q ),
    .b(\DFF_271.Q ),
    .y(_00706_)
  );
  al_nand3 _05371_ (
    .a(_00499_),
    .b(_00705_),
    .c(_00706_),
    .y(_00707_)
  );
  al_ao21 _05372_ (
    .a(_00705_),
    .b(_00706_),
    .c(\DFF_134.Q ),
    .y(_00708_)
  );
  al_nand3 _05373_ (
    .a(g35),
    .b(_00708_),
    .c(_00707_),
    .y(_00709_)
  );
  al_ao21ftf _05374_ (
    .a(g35),
    .b(\DFF_1401.Q ),
    .c(_00709_),
    .y(\DFF_134.D )
  );
  al_mux2l _05375_ (
    .a(\DFF_140.Q ),
    .b(\DFF_1388.Q ),
    .s(g84),
    .y(_00710_)
  );
  al_and3ftt _05376_ (
    .a(\DFF_586.Q ),
    .b(\DFF_703.Q ),
    .c(\DFF_805.Q ),
    .y(_00711_)
  );
  al_or3fft _05377_ (
    .a(g35),
    .b(_00711_),
    .c(_00710_),
    .y(_00712_)
  );
  al_aoi21ftf _05378_ (
    .a(\DFF_703.Q ),
    .b(_00066_),
    .c(_00712_),
    .y(\DFF_1239.D )
  );
  al_and2 _05379_ (
    .a(\DFF_529.Q ),
    .b(\DFF_819.Q ),
    .y(_00713_)
  );
  al_and3 _05380_ (
    .a(\DFF_1293.Q ),
    .b(\DFF_1038.Q ),
    .c(_00713_),
    .y(_00714_)
  );
  al_aoi21 _05381_ (
    .a(\DFF_538.Q ),
    .b(_00714_),
    .c(_00066_),
    .y(_00715_)
  );
  al_nand2ft _05382_ (
    .a(g35),
    .b(\DFF_538.Q ),
    .y(_00716_)
  );
  al_ao21ftf _05383_ (
    .a(\DFF_840.Q ),
    .b(_00715_),
    .c(_00716_),
    .y(\DFF_224.D )
  );
  al_nand3fft _05384_ (
    .a(\DFF_941.Q ),
    .b(\DFF_445.Q ),
    .c(\DFF_507.Q ),
    .y(_00717_)
  );
  al_oa21 _05385_ (
    .a(\DFF_979.Q ),
    .b(\DFF_283.Q ),
    .c(\DFF_1237.Q ),
    .y(_00718_)
  );
  al_ao21 _05386_ (
    .a(_00515_),
    .b(_00718_),
    .c(g134),
    .y(_00719_)
  );
  al_aoi21ftf _05387_ (
    .a(\DFF_1242.Q ),
    .b(\DFF_137.Q ),
    .c(_00719_),
    .y(_00720_)
  );
  al_nand3 _05388_ (
    .a(_00717_),
    .b(_00720_),
    .c(_00348_),
    .y(_00721_)
  );
  al_nand3fft _05389_ (
    .a(\DFF_646.Q ),
    .b(\DFF_1054.Q ),
    .c(_00721_),
    .y(_00722_)
  );
  al_inv _05390_ (
    .a(\DFF_828.Q ),
    .y(_00723_)
  );
  al_aoi21ftf _05391_ (
    .a(_00717_),
    .b(_00528_),
    .c(_00720_),
    .y(_00724_)
  );
  al_ao21ftf _05392_ (
    .a(_00723_),
    .b(_00717_),
    .c(_00724_),
    .y(_00725_)
  );
  al_mux2l _05393_ (
    .a(\DFF_246.Q ),
    .b(_00725_),
    .s(_00722_),
    .y(_00726_)
  );
  al_mux2h _05394_ (
    .a(\DFF_1266.Q ),
    .b(_00726_),
    .s(g35),
    .y(\DFF_246.D )
  );
  al_inv _05395_ (
    .a(\DFF_599.Q ),
    .y(_00727_)
  );
  al_and2 _05396_ (
    .a(\DFF_46.Q ),
    .b(\DFF_1335.Q ),
    .y(_00728_)
  );
  al_and3 _05397_ (
    .a(\DFF_263.Q ),
    .b(\DFF_117.Q ),
    .c(_00728_),
    .y(_00729_)
  );
  al_aoi21 _05398_ (
    .a(\DFF_599.Q ),
    .b(_00729_),
    .c(_00066_),
    .y(_00730_)
  );
  al_ao21ftf _05399_ (
    .a(_00729_),
    .b(_00727_),
    .c(_00730_),
    .y(_00731_)
  );
  al_ao21ftf _05400_ (
    .a(g35),
    .b(\DFF_666.Q ),
    .c(_00731_),
    .y(\DFF_599.D )
  );
  al_aoi21 _05401_ (
    .a(\DFF_467.Q ),
    .b(g35),
    .c(\DFF_473.Q ),
    .y(_00732_)
  );
  al_and2 _05402_ (
    .a(\DFF_473.Q ),
    .b(\DFF_467.Q ),
    .y(_00733_)
  );
  al_nand3 _05403_ (
    .a(\DFF_411.Q ),
    .b(_00556_),
    .c(_00360_),
    .y(_00734_)
  );
  al_nand2ft _05404_ (
    .a(_00733_),
    .b(_00734_),
    .y(_00735_)
  );
  al_aoi21 _05405_ (
    .a(g35),
    .b(_00735_),
    .c(_00732_),
    .y(\DFF_467.D )
  );
  al_inv _05406_ (
    .a(\DFF_538.Q ),
    .y(_00736_)
  );
  al_ao21ftf _05407_ (
    .a(_00714_),
    .b(_00736_),
    .c(_00715_),
    .y(_00737_)
  );
  al_ao21ftf _05408_ (
    .a(g35),
    .b(\DFF_1303.Q ),
    .c(_00737_),
    .y(\DFF_538.D )
  );
  al_oai21ftf _05409_ (
    .a(\DFF_1256.Q ),
    .b(\DFF_817.Q ),
    .c(\DFF_205.Q ),
    .y(_00738_)
  );
  al_nand3ftt _05410_ (
    .a(\DFF_317.Q ),
    .b(g35),
    .c(_00738_),
    .y(_00739_)
  );
  al_ao21ftf _05411_ (
    .a(g35),
    .b(\DFF_817.Q ),
    .c(_00739_),
    .y(\DFF_205.D )
  );
  al_oa21ftt _05412_ (
    .a(g35),
    .b(\DFF_701.Q ),
    .c(\DFF_495.Q ),
    .y(_00740_)
  );
  al_nand2ft _05413_ (
    .a(\DFF_1385.Q ),
    .b(\DFF_631.Q ),
    .y(_00741_)
  );
  al_oa21ftf _05414_ (
    .a(\DFF_631.Q ),
    .b(\DFF_548.Q ),
    .c(\DFF_701.Q ),
    .y(_00742_)
  );
  al_ao21ftf _05415_ (
    .a(\DFF_495.Q ),
    .b(_00742_),
    .c(_00741_),
    .y(_00743_)
  );
  al_ao21 _05416_ (
    .a(g35),
    .b(_00743_),
    .c(_00740_),
    .y(\DFF_701.D )
  );
  al_and3ftt _05417_ (
    .a(g113),
    .b(\DFF_796.Q ),
    .c(_00342_),
    .y(_00744_)
  );
  al_nand3 _05418_ (
    .a(_00391_),
    .b(_00744_),
    .c(_00386_),
    .y(_00745_)
  );
  al_oa21ftt _05419_ (
    .a(g35),
    .b(_00745_),
    .c(\DFF_792.Q ),
    .y(\DFF_107.D )
  );
  al_and2ft _05420_ (
    .a(g35),
    .b(\DFF_934.Q ),
    .y(_00746_)
  );
  al_or3 _05421_ (
    .a(\DFF_1379.Q ),
    .b(\DFF_115.Q ),
    .c(\DFF_1084.Q ),
    .y(_00747_)
  );
  al_and2 _05422_ (
    .a(\DFF_186.Q ),
    .b(g35),
    .y(_00748_)
  );
  al_nand3fft _05423_ (
    .a(\DFF_853.Q ),
    .b(_00747_),
    .c(_00748_),
    .y(_00749_)
  );
  al_oai21ftf _05424_ (
    .a(_00410_),
    .b(_00749_),
    .c(_00746_),
    .y(\DFF_607.D )
  );
  al_nand3 _05425_ (
    .a(\DFF_607.Q ),
    .b(\DFF_724.Q ),
    .c(g35),
    .y(_00750_)
  );
  al_oa21 _05426_ (
    .a(g35),
    .b(\DFF_1296.Q ),
    .c(_00750_),
    .y(\DFF_79.D )
  );
  al_or2 _05427_ (
    .a(\DFF_1391.Q ),
    .b(\DFF_708.Q ),
    .y(_00751_)
  );
  al_mux2h _05428_ (
    .a(\DFF_597.Q ),
    .b(_00751_),
    .s(g35),
    .y(\DFF_1391.D )
  );
  al_nand3ftt _05429_ (
    .a(\DFF_1408.Q ),
    .b(\DFF_245.Q ),
    .c(\DFF_199.Q ),
    .y(_00752_)
  );
  al_aoi21ftf _05430_ (
    .a(\DFF_738.Q ),
    .b(_00752_),
    .c(g35),
    .y(_00753_)
  );
  al_ao21ftf _05431_ (
    .a(_00752_),
    .b(_00499_),
    .c(_00753_),
    .y(_00754_)
  );
  al_ao21ftf _05432_ (
    .a(g35),
    .b(\DFF_102.Q ),
    .c(_00754_),
    .y(\DFF_738.D )
  );
  al_inv _05433_ (
    .a(\DFF_233.Q ),
    .y(_00755_)
  );
  al_and2 _05434_ (
    .a(\DFF_893.Q ),
    .b(\DFF_962.Q ),
    .y(_00756_)
  );
  al_and2 _05435_ (
    .a(_00756_),
    .b(_00544_),
    .y(_00757_)
  );
  al_aoi21ftf _05436_ (
    .a(_00755_),
    .b(_00542_),
    .c(_00757_),
    .y(_00758_)
  );
  al_and2 _05437_ (
    .a(\DFF_623.Q ),
    .b(\DFF_562.Q ),
    .y(_00759_)
  );
  al_nand2 _05438_ (
    .a(_00759_),
    .b(_00758_),
    .y(_00760_)
  );
  al_nand2 _05439_ (
    .a(\DFF_933.Q ),
    .b(\DFF_1267.Q ),
    .y(_00761_)
  );
  al_nor2 _05440_ (
    .a(\DFF_933.Q ),
    .b(\DFF_1267.Q ),
    .y(_00762_)
  );
  al_nand2ft _05441_ (
    .a(_00762_),
    .b(_00761_),
    .y(_00763_)
  );
  al_mux2l _05442_ (
    .a(\DFF_1140.Q ),
    .b(_00763_),
    .s(_00760_),
    .y(_00764_)
  );
  al_mux2h _05443_ (
    .a(\DFF_1267.Q ),
    .b(_00764_),
    .s(g35),
    .y(\DFF_1140.D )
  );
  al_and3ftt _05444_ (
    .a(\DFF_1199.Q ),
    .b(\DFF_892.Q ),
    .c(\DFF_684.Q ),
    .y(_00765_)
  );
  al_aoi21ttf _05445_ (
    .a(_00765_),
    .b(_00584_),
    .c(\DFF_160.Q ),
    .y(_00766_)
  );
  al_inv _05446_ (
    .a(\DFF_664.Q ),
    .y(_00767_)
  );
  al_nand2ft _05447_ (
    .a(\DFF_536.Q ),
    .b(\DFF_1312.Q ),
    .y(_00768_)
  );
  al_nand2 _05448_ (
    .a(\DFF_81.Q ),
    .b(\DFF_19.Q ),
    .y(_00769_)
  );
  al_nand2 _05449_ (
    .a(\DFF_102.Q ),
    .b(\DFF_1300.Q ),
    .y(_00770_)
  );
  al_ao21 _05450_ (
    .a(_00769_),
    .b(_00770_),
    .c(_00768_),
    .y(_00771_)
  );
  al_nor2 _05451_ (
    .a(\DFF_1312.Q ),
    .b(\DFF_536.Q ),
    .y(_00772_)
  );
  al_nand3 _05452_ (
    .a(\DFF_1052.Q ),
    .b(\DFF_369.Q ),
    .c(_00772_),
    .y(_00773_)
  );
  al_and3 _05453_ (
    .a(_00767_),
    .b(_00773_),
    .c(_00771_),
    .y(_00774_)
  );
  al_nand2 _05454_ (
    .a(\DFF_321.Q ),
    .b(\DFF_873.Q ),
    .y(_00775_)
  );
  al_nand2 _05455_ (
    .a(\DFF_1420.Q ),
    .b(\DFF_309.Q ),
    .y(_00776_)
  );
  al_ao21ttf _05456_ (
    .a(_00775_),
    .b(_00776_),
    .c(_00402_),
    .y(_00777_)
  );
  al_nand2ft _05457_ (
    .a(\DFF_1312.Q ),
    .b(\DFF_536.Q ),
    .y(_00778_)
  );
  al_nand2 _05458_ (
    .a(\DFF_738.Q ),
    .b(\DFF_290.Q ),
    .y(_00779_)
  );
  al_ao21ttf _05459_ (
    .a(\DFF_1259.Q ),
    .b(\DFF_34.Q ),
    .c(_00779_),
    .y(_00780_)
  );
  al_ao21ftf _05460_ (
    .a(_00778_),
    .b(_00780_),
    .c(_00777_),
    .y(_00781_)
  );
  al_nand3 _05461_ (
    .a(\DFF_72.Q ),
    .b(\DFF_1300.Q ),
    .c(_00402_),
    .y(_00782_)
  );
  al_or3fft _05462_ (
    .a(\DFF_633.Q ),
    .b(\DFF_369.Q ),
    .c(_00778_),
    .y(_00783_)
  );
  al_and3 _05463_ (
    .a(\DFF_664.Q ),
    .b(_00783_),
    .c(_00782_),
    .y(_00784_)
  );
  al_nand2 _05464_ (
    .a(\DFF_707.Q ),
    .b(\DFF_34.Q ),
    .y(_00785_)
  );
  al_nand2 _05465_ (
    .a(\DFF_982.Q ),
    .b(\DFF_290.Q ),
    .y(_00786_)
  );
  al_ao21ttf _05466_ (
    .a(_00785_),
    .b(_00786_),
    .c(_00772_),
    .y(_00787_)
  );
  al_nand2 _05467_ (
    .a(\DFF_227.Q ),
    .b(\DFF_873.Q ),
    .y(_00788_)
  );
  al_nand2 _05468_ (
    .a(\DFF_1420.Q ),
    .b(\DFF_12.Q ),
    .y(_00789_)
  );
  al_ao21 _05469_ (
    .a(_00788_),
    .b(_00789_),
    .c(_00768_),
    .y(_00790_)
  );
  al_nand3 _05470_ (
    .a(_00787_),
    .b(_00790_),
    .c(_00784_),
    .y(_00791_)
  );
  al_ao21ftf _05471_ (
    .a(_00781_),
    .b(_00774_),
    .c(_00791_),
    .y(_00792_)
  );
  al_and3 _05472_ (
    .a(\DFF_664.Q ),
    .b(\DFF_81.Q ),
    .c(_00402_),
    .y(_00793_)
  );
  al_nor3fft _05473_ (
    .a(\DFF_468.Q ),
    .b(\DFF_108.Q ),
    .c(_00778_),
    .y(_00794_)
  );
  al_and3 _05474_ (
    .a(\DFF_220.Q ),
    .b(\DFF_626.Q ),
    .c(_00772_),
    .y(_00795_)
  );
  al_nor2 _05475_ (
    .a(\DFF_1420.Q ),
    .b(\DFF_664.Q ),
    .y(_00796_)
  );
  al_nand2 _05476_ (
    .a(\DFF_1420.Q ),
    .b(\DFF_664.Q ),
    .y(_00797_)
  );
  al_nand2ft _05477_ (
    .a(_00796_),
    .b(_00797_),
    .y(_00798_)
  );
  al_nand3 _05478_ (
    .a(\DFF_942.Q ),
    .b(\DFF_105.Q ),
    .c(_00402_),
    .y(_00799_)
  );
  al_and3ftt _05479_ (
    .a(_00795_),
    .b(_00799_),
    .c(_00798_),
    .y(_00800_)
  );
  al_nor3fft _05480_ (
    .a(\DFF_220.Q ),
    .b(\DFF_1177.Q ),
    .c(_00778_),
    .y(_00801_)
  );
  al_and3 _05481_ (
    .a(\DFF_468.Q ),
    .b(\DFF_628.Q ),
    .c(_00772_),
    .y(_00802_)
  );
  al_or3fft _05482_ (
    .a(\DFF_942.Q ),
    .b(\DFF_1244.Q ),
    .c(_00768_),
    .y(_00803_)
  );
  al_and3ftt _05483_ (
    .a(_00796_),
    .b(_00797_),
    .c(_00803_),
    .y(_00804_)
  );
  al_nand3fft _05484_ (
    .a(_00801_),
    .b(_00802_),
    .c(_00804_),
    .y(_00805_)
  );
  al_ao21ftf _05485_ (
    .a(_00794_),
    .b(_00800_),
    .c(_00805_),
    .y(_00806_)
  );
  al_aoi21ttf _05486_ (
    .a(\DFF_1356.Q ),
    .b(_00793_),
    .c(_00806_),
    .y(_00807_)
  );
  al_ao21ttf _05487_ (
    .a(_00792_),
    .b(_00807_),
    .c(_00766_),
    .y(_00808_)
  );
  al_nand2 _05488_ (
    .a(_00793_),
    .b(_00766_),
    .y(_00809_)
  );
  al_nand3 _05489_ (
    .a(\DFF_58.Q ),
    .b(_00809_),
    .c(_00808_),
    .y(_00810_)
  );
  al_ao21 _05490_ (
    .a(\DFF_58.Q ),
    .b(_00809_),
    .c(_00808_),
    .y(_00811_)
  );
  al_nand3 _05491_ (
    .a(g35),
    .b(_00810_),
    .c(_00811_),
    .y(_00812_)
  );
  al_aoi21ftf _05492_ (
    .a(\DFF_1134.Q ),
    .b(_00066_),
    .c(_00812_),
    .y(\DFF_58.D )
  );
  al_mux2l _05493_ (
    .a(\DFF_1282.Q ),
    .b(\DFF_1289.Q ),
    .s(g35),
    .y(\DFF_1282.D )
  );
  al_oai21ftf _05494_ (
    .a(\DFF_503.Q ),
    .b(\DFF_569.Q ),
    .c(\DFF_1392.Q ),
    .y(_00813_)
  );
  al_nand3ftt _05495_ (
    .a(\DFF_630.Q ),
    .b(g35),
    .c(_00813_),
    .y(_00814_)
  );
  al_ao21ftf _05496_ (
    .a(g35),
    .b(\DFF_569.Q ),
    .c(_00814_),
    .y(\DFF_1392.D )
  );
  al_nand2 _05497_ (
    .a(_00577_),
    .b(_00440_),
    .y(_00815_)
  );
  al_ao21 _05498_ (
    .a(_00563_),
    .b(_00815_),
    .c(_00066_),
    .y(_00816_)
  );
  al_inv _05499_ (
    .a(\DFF_793.Q ),
    .y(_00817_)
  );
  al_and3fft _05500_ (
    .a(_00066_),
    .b(_00563_),
    .c(_00817_),
    .y(_00818_)
  );
  al_aoi21 _05501_ (
    .a(_00559_),
    .b(_00816_),
    .c(_00818_),
    .y(\DFF_793.D )
  );
  al_and2ft _05502_ (
    .a(g35),
    .b(\DFF_1153.Q ),
    .y(_00819_)
  );
  al_inv _05503_ (
    .a(\DFF_1039.Q ),
    .y(_00820_)
  );
  al_nand2ft _05504_ (
    .a(\DFF_990.Q ),
    .b(\DFF_67.Q ),
    .y(_00821_)
  );
  al_nand2ft _05505_ (
    .a(\DFF_67.Q ),
    .b(\DFF_990.Q ),
    .y(_00822_)
  );
  al_nand2 _05506_ (
    .a(_00821_),
    .b(_00822_),
    .y(_00823_)
  );
  al_nand3 _05507_ (
    .a(\DFF_1343.Q ),
    .b(\DFF_577.Q ),
    .c(\DFF_316.Q ),
    .y(_00824_)
  );
  al_mux2l _05508_ (
    .a(\DFF_1343.Q ),
    .b(_00824_),
    .s(_00823_),
    .y(_00825_)
  );
  al_ao21ttf _05509_ (
    .a(_00821_),
    .b(_00822_),
    .c(\DFF_211.Q ),
    .y(_00826_)
  );
  al_and3 _05510_ (
    .a(_00820_),
    .b(_00826_),
    .c(_00825_),
    .y(_00827_)
  );
  al_inv _05511_ (
    .a(\DFF_1153.Q ),
    .y(_00828_)
  );
  al_or2 _05512_ (
    .a(\DFF_408.Q ),
    .b(\DFF_990.Q ),
    .y(_00829_)
  );
  al_ao21ttf _05513_ (
    .a(_00828_),
    .b(_00827_),
    .c(_00829_),
    .y(_00830_)
  );
  al_aoi21ftt _05514_ (
    .a(\DFF_577.Q ),
    .b(_00827_),
    .c(_00830_),
    .y(_00831_)
  );
  al_aoi21ftf _05515_ (
    .a(\DFF_577.Q ),
    .b(_00830_),
    .c(g35),
    .y(_00832_)
  );
  al_ao21ftt _05516_ (
    .a(_00831_),
    .b(_00832_),
    .c(_00819_),
    .y(\DFF_577.D )
  );
  al_and2 _05517_ (
    .a(\DFF_64.Q ),
    .b(g35),
    .y(\DFF_64.D )
  );
  al_aoi21 _05518_ (
    .a(\DFF_292.Q ),
    .b(\DFF_533.Q ),
    .c(\DFF_1045.Q ),
    .y(_00833_)
  );
  al_oa21 _05519_ (
    .a(\DFF_292.Q ),
    .b(\DFF_533.Q ),
    .c(g35),
    .y(_00834_)
  );
  al_and3ftt _05520_ (
    .a(_00833_),
    .b(_00475_),
    .c(_00834_),
    .y(\DFF_252.D )
  );
  al_inv _05521_ (
    .a(\DFF_283.Q ),
    .y(_00835_)
  );
  al_nand2ft _05522_ (
    .a(\DFF_606.Q ),
    .b(\DFF_698.Q ),
    .y(_00836_)
  );
  al_nand2ft _05523_ (
    .a(\DFF_698.Q ),
    .b(\DFF_606.Q ),
    .y(_00837_)
  );
  al_ao21ttf _05524_ (
    .a(_00836_),
    .b(_00837_),
    .c(\DFF_1144.Q ),
    .y(_00838_)
  );
  al_nand2 _05525_ (
    .a(_00836_),
    .b(_00837_),
    .y(_00839_)
  );
  al_nand3 _05526_ (
    .a(\DFF_979.Q ),
    .b(\DFF_368.Q ),
    .c(\DFF_421.Q ),
    .y(_00840_)
  );
  al_mux2l _05527_ (
    .a(\DFF_979.Q ),
    .b(_00840_),
    .s(_00839_),
    .y(_00841_)
  );
  al_and3 _05528_ (
    .a(_00835_),
    .b(_00838_),
    .c(_00841_),
    .y(_00842_)
  );
  al_inv _05529_ (
    .a(\DFF_788.Q ),
    .y(_00843_)
  );
  al_or2 _05530_ (
    .a(\DFF_698.Q ),
    .b(\DFF_511.Q ),
    .y(_00844_)
  );
  al_aoi21ttf _05531_ (
    .a(_00843_),
    .b(_00842_),
    .c(_00844_),
    .y(_00845_)
  );
  al_aoi21ftf _05532_ (
    .a(\DFF_421.Q ),
    .b(_00842_),
    .c(_00845_),
    .y(_00846_)
  );
  al_ao21ftf _05533_ (
    .a(\DFF_70.Q ),
    .b(_00842_),
    .c(_00846_),
    .y(_00847_)
  );
  al_ao21ftt _05534_ (
    .a(\DFF_368.Q ),
    .b(_00842_),
    .c(_00847_),
    .y(_00848_)
  );
  al_and2ft _05535_ (
    .a(\DFF_131.Q ),
    .b(_00842_),
    .y(_00849_)
  );
  al_mux2l _05536_ (
    .a(\DFF_131.Q ),
    .b(_00849_),
    .s(_00848_),
    .y(_00850_)
  );
  al_mux2h _05537_ (
    .a(\DFF_368.Q ),
    .b(_00850_),
    .s(g35),
    .y(\DFF_131.D )
  );
  al_nand3fft _05538_ (
    .a(\DFF_1324.Q ),
    .b(\DFF_891.Q ),
    .c(_00305_),
    .y(_00851_)
  );
  al_nor2 _05539_ (
    .a(\DFF_154.Q ),
    .b(_00306_),
    .y(_00852_)
  );
  al_ao21ftt _05540_ (
    .a(_00851_),
    .b(_00852_),
    .c(_00066_),
    .y(_00853_)
  );
  al_mux2l _05541_ (
    .a(\DFF_282.Q ),
    .b(\DFF_1152.Q ),
    .s(_00853_),
    .y(\DFF_1152.D )
  );
  al_and2ft _05542_ (
    .a(g35),
    .b(\DFF_1328.Q ),
    .y(_00854_)
  );
  al_and2ft _05543_ (
    .a(\DFF_993.Q ),
    .b(\DFF_889.Q ),
    .y(_00855_)
  );
  al_nand2 _05544_ (
    .a(_00855_),
    .b(_00576_),
    .y(_00856_)
  );
  al_nand2ft _05545_ (
    .a(\DFF_1050.Q ),
    .b(\DFF_1328.Q ),
    .y(_00857_)
  );
  al_nand2ft _05546_ (
    .a(\DFF_1328.Q ),
    .b(\DFF_1050.Q ),
    .y(_00858_)
  );
  al_or3fft _05547_ (
    .a(_00857_),
    .b(_00858_),
    .c(_00856_),
    .y(_00859_)
  );
  al_aoi21ftf _05548_ (
    .a(\DFF_301.Q ),
    .b(_00856_),
    .c(g35),
    .y(_00860_)
  );
  al_ao21 _05549_ (
    .a(_00859_),
    .b(_00860_),
    .c(_00854_),
    .y(\DFF_301.D )
  );
  al_or3 _05550_ (
    .a(\DFF_1338.Q ),
    .b(\DFF_944.Q ),
    .c(\DFF_418.Q ),
    .y(_00861_)
  );
  al_or3 _05551_ (
    .a(\DFF_992.Q ),
    .b(\DFF_389.Q ),
    .c(_00861_),
    .y(_00862_)
  );
  al_or3 _05552_ (
    .a(\DFF_485.Q ),
    .b(\DFF_1286.Q ),
    .c(_00862_),
    .y(_00863_)
  );
  al_nor2 _05553_ (
    .a(\DFF_31.Q ),
    .b(\DFF_885.Q ),
    .y(_00864_)
  );
  al_ao21ttf _05554_ (
    .a(\DFF_31.Q ),
    .b(\DFF_885.Q ),
    .c(g35),
    .y(_00865_)
  );
  al_ao21 _05555_ (
    .a(_00864_),
    .b(_00863_),
    .c(_00865_),
    .y(_00866_)
  );
  al_mux2l _05556_ (
    .a(\DFF_282.Q ),
    .b(\DFF_1230.Q ),
    .s(\DFF_1340.Q ),
    .y(_00867_)
  );
  al_inv _05557_ (
    .a(_00867_),
    .y(_00868_)
  );
  al_mux2h _05558_ (
    .a(\DFF_31.Q ),
    .b(_00868_),
    .s(g35),
    .y(_00869_)
  );
  al_mux2l _05559_ (
    .a(_00869_),
    .b(_00867_),
    .s(_00866_),
    .y(\DFF_919.D )
  );
  al_and3fft _05560_ (
    .a(\DFF_622.Q ),
    .b(\DFF_353.Q ),
    .c(\DFF_786.Q ),
    .y(_00870_)
  );
  al_nand3 _05561_ (
    .a(\DFF_47.Q ),
    .b(\DFF_1145.Q ),
    .c(_00870_),
    .y(_00871_)
  );
  al_nor3fft _05562_ (
    .a(\DFF_1161.Q ),
    .b(_00477_),
    .c(_00871_),
    .y(_00872_)
  );
  al_nor2 _05563_ (
    .a(\DFF_1365.Q ),
    .b(\DFF_573.Q ),
    .y(_00873_)
  );
  al_inv _05564_ (
    .a(_00873_),
    .y(_00874_)
  );
  al_mux2l _05565_ (
    .a(_00874_),
    .b(\DFF_1044.Q ),
    .s(_00872_),
    .y(_00875_)
  );
  al_mux2h _05566_ (
    .a(\DFF_1365.Q ),
    .b(_00875_),
    .s(g35),
    .y(\DFF_1044.D )
  );
  al_nand3fft _05567_ (
    .a(\DFF_1091.Q ),
    .b(_00448_),
    .c(_00576_),
    .y(_00876_)
  );
  al_and2ft _05568_ (
    .a(\DFF_769.Q ),
    .b(\DFF_1141.Q ),
    .y(_00877_)
  );
  al_inv _05569_ (
    .a(\DFF_570.Q ),
    .y(_00878_)
  );
  al_aoi21 _05570_ (
    .a(_00878_),
    .b(_00876_),
    .c(_00066_),
    .y(_00879_)
  );
  al_ao21ftf _05571_ (
    .a(_00876_),
    .b(_00877_),
    .c(_00879_),
    .y(_00880_)
  );
  al_ao21ftf _05572_ (
    .a(g35),
    .b(\DFF_1026.Q ),
    .c(_00880_),
    .y(\DFF_570.D )
  );
  al_and3 _05573_ (
    .a(\DFF_305.Q ),
    .b(\DFF_1001.Q ),
    .c(\DFF_401.Q ),
    .y(_00881_)
  );
  al_and2 _05574_ (
    .a(\DFF_181.Q ),
    .b(_00881_),
    .y(_00882_)
  );
  al_and2 _05575_ (
    .a(\DFF_5.Q ),
    .b(g35),
    .y(_00883_)
  );
  al_aoi21ttf _05576_ (
    .a(_00883_),
    .b(_00882_),
    .c(\DFF_423.Q ),
    .y(\DFF_347.D )
  );
  al_nand2ft _05577_ (
    .a(\DFF_466.Q ),
    .b(\DFF_572.Q ),
    .y(_00884_)
  );
  al_nand3 _05578_ (
    .a(\DFF_636.Q ),
    .b(g35),
    .c(_00884_),
    .y(_00885_)
  );
  al_nand2ft _05579_ (
    .a(\DFF_1333.Q ),
    .b(\DFF_572.Q ),
    .y(_00886_)
  );
  al_mux2l _05580_ (
    .a(\DFF_636.Q ),
    .b(\DFF_572.Q ),
    .s(g35),
    .y(_00887_)
  );
  al_aoi21ftf _05581_ (
    .a(_00887_),
    .b(_00886_),
    .c(_00885_),
    .y(\DFF_415.D )
  );
  al_nor2 _05582_ (
    .a(\DFF_49.Q ),
    .b(g35),
    .y(_00888_)
  );
  al_inv _05583_ (
    .a(\DFF_998.Q ),
    .y(_00889_)
  );
  al_inv _05584_ (
    .a(g84),
    .y(_00890_)
  );
  al_nand2 _05585_ (
    .a(\DFF_1321.Q ),
    .b(\DFF_97.Q ),
    .y(_00891_)
  );
  al_nand2 _05586_ (
    .a(\DFF_712.Q ),
    .b(\DFF_1321.Q ),
    .y(_00892_)
  );
  al_mux2l _05587_ (
    .a(_00891_),
    .b(_00892_),
    .s(_00890_),
    .y(_00893_)
  );
  al_or3fft _05588_ (
    .a(\DFF_838.Q ),
    .b(_00889_),
    .c(_00893_),
    .y(_00894_)
  );
  al_nor2 _05589_ (
    .a(\DFF_1321.Q ),
    .b(\DFF_97.Q ),
    .y(_00895_)
  );
  al_nor2 _05590_ (
    .a(\DFF_712.Q ),
    .b(\DFF_1321.Q ),
    .y(_00896_)
  );
  al_mux2l _05591_ (
    .a(_00895_),
    .b(_00896_),
    .s(_00890_),
    .y(_00897_)
  );
  al_nand3 _05592_ (
    .a(\DFF_998.Q ),
    .b(\DFF_1048.Q ),
    .c(_00897_),
    .y(_00898_)
  );
  al_and2 _05593_ (
    .a(_00898_),
    .b(_00894_),
    .y(_00899_)
  );
  al_and3 _05594_ (
    .a(\DFF_838.Q ),
    .b(\DFF_122.Q ),
    .c(\DFF_851.Q ),
    .y(_00900_)
  );
  al_and3fft _05595_ (
    .a(\DFF_122.Q ),
    .b(\DFF_851.Q ),
    .c(\DFF_1048.Q ),
    .y(_00901_)
  );
  al_mux2h _05596_ (
    .a(_00901_),
    .b(_00900_),
    .s(\DFF_49.Q ),
    .y(_00902_)
  );
  al_nand3ftt _05597_ (
    .a(_00902_),
    .b(\DFF_40.Q ),
    .c(_00899_),
    .y(_00903_)
  );
  al_aoi21ftf _05598_ (
    .a(\DFF_40.Q ),
    .b(_00902_),
    .c(g35),
    .y(_00904_)
  );
  al_aoi21 _05599_ (
    .a(_00904_),
    .b(_00903_),
    .c(_00888_),
    .y(\DFF_40.D )
  );
  al_and2ft _05600_ (
    .a(\DFF_1393.Q ),
    .b(\DFF_1161.Q ),
    .y(_00905_)
  );
  al_nand3 _05601_ (
    .a(\DFF_1232.Q ),
    .b(\DFF_269.Q ),
    .c(_00905_),
    .y(_00906_)
  );
  al_aoi21ttf _05602_ (
    .a(\DFF_1053.Q ),
    .b(\DFF_601.Q ),
    .c(\DFF_239.Q ),
    .y(_00907_)
  );
  al_oai21 _05603_ (
    .a(\DFF_1053.Q ),
    .b(\DFF_601.Q ),
    .c(_00907_),
    .y(_00908_)
  );
  al_and3 _05604_ (
    .a(\DFF_1053.Q ),
    .b(\DFF_601.Q ),
    .c(\DFF_542.Q ),
    .y(_00909_)
  );
  al_nand3fft _05605_ (
    .a(\DFF_1053.Q ),
    .b(\DFF_601.Q ),
    .c(\DFF_1108.Q ),
    .y(_00910_)
  );
  al_and3ftt _05606_ (
    .a(_00909_),
    .b(_00910_),
    .c(_00908_),
    .y(_00911_)
  );
  al_nand2ft _05607_ (
    .a(\DFF_237.Q ),
    .b(_00911_),
    .y(_00912_)
  );
  al_mux2l _05608_ (
    .a(\DFF_10.Q ),
    .b(\DFF_292.Q ),
    .s(\DFF_1053.Q ),
    .y(_00913_)
  );
  al_nand2ft _05609_ (
    .a(\DFF_1053.Q ),
    .b(\DFF_1315.Q ),
    .y(_00914_)
  );
  al_aoi21 _05610_ (
    .a(\DFF_1053.Q ),
    .b(\DFF_544.Q ),
    .c(\DFF_237.Q ),
    .y(_00915_)
  );
  al_nand3ftt _05611_ (
    .a(\DFF_1390.Q ),
    .b(_00914_),
    .c(_00915_),
    .y(_00916_)
  );
  al_aoi21 _05612_ (
    .a(\DFF_1045.Q ),
    .b(_00913_),
    .c(_00916_),
    .y(_00917_)
  );
  al_oa21 _05613_ (
    .a(\DFF_1045.Q ),
    .b(_00913_),
    .c(_00917_),
    .y(_00918_)
  );
  al_aoi21ftt _05614_ (
    .a(_00911_),
    .b(\DFF_237.Q ),
    .c(_00918_),
    .y(_00919_)
  );
  al_aoi21 _05615_ (
    .a(_00912_),
    .b(_00919_),
    .c(_00906_),
    .y(_00920_)
  );
  al_nand3 _05616_ (
    .a(g35),
    .b(\DFF_719.Q ),
    .c(_00906_),
    .y(_00921_)
  );
  al_ao21ttf _05617_ (
    .a(g35),
    .b(_00920_),
    .c(_00921_),
    .y(\DFF_719.D )
  );
  al_nand3ftt _05618_ (
    .a(\DFF_522.Q ),
    .b(\DFF_271.Q ),
    .c(\DFF_54.Q ),
    .y(_00922_)
  );
  al_aoi21ftf _05619_ (
    .a(\DFF_1351.Q ),
    .b(_00922_),
    .c(g35),
    .y(_00923_)
  );
  al_ao21ftf _05620_ (
    .a(_00922_),
    .b(_00499_),
    .c(_00923_),
    .y(_00924_)
  );
  al_ao21ftf _05621_ (
    .a(g35),
    .b(\DFF_1280.Q ),
    .c(_00924_),
    .y(\DFF_1351.D )
  );
  al_nor2 _05622_ (
    .a(\DFF_346.Q ),
    .b(\DFF_362.Q ),
    .y(_00925_)
  );
  al_and2ft _05623_ (
    .a(\DFF_382.Q ),
    .b(\DFF_771.Q ),
    .y(_00926_)
  );
  al_nand2 _05624_ (
    .a(\DFF_541.Q ),
    .b(\DFF_648.Q ),
    .y(_00927_)
  );
  al_and3fft _05625_ (
    .a(\DFF_496.Q ),
    .b(_00927_),
    .c(_00926_),
    .y(_00928_)
  );
  al_ao21 _05626_ (
    .a(_00925_),
    .b(_00928_),
    .c(\DFF_128.Q ),
    .y(_00929_)
  );
  al_nand3ftt _05627_ (
    .a(\DFF_771.Q ),
    .b(\DFF_382.Q ),
    .c(\DFF_496.Q ),
    .y(_00930_)
  );
  al_nor2 _05628_ (
    .a(\DFF_541.Q ),
    .b(\DFF_648.Q ),
    .y(_00931_)
  );
  al_and2 _05629_ (
    .a(\DFF_346.Q ),
    .b(\DFF_362.Q ),
    .y(_00932_)
  );
  al_nand3ftt _05630_ (
    .a(_00930_),
    .b(_00931_),
    .c(_00932_),
    .y(_00933_)
  );
  al_aoi21ttf _05631_ (
    .a(\DFF_128.Q ),
    .b(_00933_),
    .c(_00929_),
    .y(_00934_)
  );
  al_and3 _05632_ (
    .a(\DFF_1390.Q ),
    .b(_00486_),
    .c(_00934_),
    .y(_00935_)
  );
  al_and3 _05633_ (
    .a(\DFF_745.Q ),
    .b(\DFF_106.Q ),
    .c(\DFF_802.Q ),
    .y(_00936_)
  );
  al_and3 _05634_ (
    .a(\DFF_83.Q ),
    .b(_00936_),
    .c(_00935_),
    .y(_00937_)
  );
  al_oai21 _05635_ (
    .a(\DFF_83.Q ),
    .b(_00936_),
    .c(_00935_),
    .y(_00938_)
  );
  al_or3 _05636_ (
    .a(_00066_),
    .b(_00938_),
    .c(_00937_),
    .y(_00939_)
  );
  al_ao21ftf _05637_ (
    .a(g35),
    .b(\DFF_106.Q ),
    .c(_00939_),
    .y(\DFF_83.D )
  );
  al_oai21ftt _05638_ (
    .a(\DFF_1081.Q ),
    .b(\DFF_256.Q ),
    .c(\DFF_661.Q ),
    .y(_00940_)
  );
  al_nand2ft _05639_ (
    .a(\DFF_256.Q ),
    .b(\DFF_1081.Q ),
    .y(_00941_)
  );
  al_and3 _05640_ (
    .a(\DFF_74.Q ),
    .b(\DFF_50.Q ),
    .c(_00941_),
    .y(_00942_)
  );
  al_oa21ftt _05641_ (
    .a(\DFF_1081.Q ),
    .b(\DFF_256.Q ),
    .c(\DFF_28.Q ),
    .y(_00943_)
  );
  al_nand3 _05642_ (
    .a(\DFF_135.Q ),
    .b(\DFF_194.Q ),
    .c(\DFF_656.Q ),
    .y(_00944_)
  );
  al_aoi21ttf _05643_ (
    .a(\DFF_142.Q ),
    .b(\DFF_21.Q ),
    .c(_00944_),
    .y(_00945_)
  );
  al_or3 _05644_ (
    .a(\DFF_135.Q ),
    .b(\DFF_194.Q ),
    .c(\DFF_656.Q ),
    .y(_00946_)
  );
  al_and3 _05645_ (
    .a(_00945_),
    .b(_00946_),
    .c(_00481_),
    .y(_00947_)
  );
  al_nand2ft _05646_ (
    .a(\DFF_1081.Q ),
    .b(\DFF_515.Q ),
    .y(_00948_)
  );
  al_and3 _05647_ (
    .a(\DFF_876.Q ),
    .b(_00948_),
    .c(_00947_),
    .y(_00949_)
  );
  al_and2 _05648_ (
    .a(\DFF_175.Q ),
    .b(_00949_),
    .y(_00950_)
  );
  al_and3 _05649_ (
    .a(\DFF_328.Q ),
    .b(_00943_),
    .c(_00950_),
    .y(_00951_)
  );
  al_and3 _05650_ (
    .a(\DFF_157.Q ),
    .b(_00942_),
    .c(_00951_),
    .y(_00952_)
  );
  al_and3 _05651_ (
    .a(\DFF_896.Q ),
    .b(\DFF_789.Q ),
    .c(_00952_),
    .y(_00953_)
  );
  al_and3 _05652_ (
    .a(\DFF_1200.Q ),
    .b(\DFF_953.Q ),
    .c(_00953_),
    .y(_00954_)
  );
  al_oa21ftf _05653_ (
    .a(_00940_),
    .b(_00954_),
    .c(_00066_),
    .y(_00955_)
  );
  al_ao21ftf _05654_ (
    .a(_00940_),
    .b(_00954_),
    .c(_00955_),
    .y(_00956_)
  );
  al_ao21ftf _05655_ (
    .a(g35),
    .b(\DFF_1200.Q ),
    .c(_00956_),
    .y(\DFF_661.D )
  );
  al_oai21ftt _05656_ (
    .a(g35),
    .b(\DFF_827.Q ),
    .c(\DFF_775.Q ),
    .y(_00957_)
  );
  al_ao21ttf _05657_ (
    .a(\DFF_1156.Q ),
    .b(g35),
    .c(_00957_),
    .y(_00958_)
  );
  al_and3 _05658_ (
    .a(\DFF_775.Q ),
    .b(\DFF_827.Q ),
    .c(g35),
    .y(_00959_)
  );
  al_aoi21ttf _05659_ (
    .a(\DFF_1156.Q ),
    .b(_00959_),
    .c(_00958_),
    .y(\DFF_1156.D )
  );
  al_or2 _05660_ (
    .a(\DFF_1039.Q ),
    .b(\DFF_1343.Q ),
    .y(_00960_)
  );
  al_nand3 _05661_ (
    .a(\DFF_1419.Q ),
    .b(\DFF_1153.Q ),
    .c(\DFF_1227.Q ),
    .y(_00961_)
  );
  al_and3ftt _05662_ (
    .a(_00961_),
    .b(_00821_),
    .c(_00822_),
    .y(_00962_)
  );
  al_ao21 _05663_ (
    .a(_00829_),
    .b(_00962_),
    .c(_00960_),
    .y(_00963_)
  );
  al_nand3ftt _05664_ (
    .a(\DFF_202.Q ),
    .b(\DFF_1407.Q ),
    .c(\DFF_67.Q ),
    .y(_00964_)
  );
  al_and3ftt _05665_ (
    .a(_00964_),
    .b(\DFF_60.Q ),
    .c(_00963_),
    .y(_00965_)
  );
  al_and3 _05666_ (
    .a(\DFF_60.Q ),
    .b(_00964_),
    .c(_00521_),
    .y(_00966_)
  );
  al_nand3 _05667_ (
    .a(\DFF_614.Q ),
    .b(\DFF_1189.Q ),
    .c(_00966_),
    .y(_00967_)
  );
  al_oai21ftf _05668_ (
    .a(\DFF_1159.Q ),
    .b(_00967_),
    .c(_00066_),
    .y(_00968_)
  );
  al_oai21ttf _05669_ (
    .a(\DFF_1159.Q ),
    .b(_00965_),
    .c(_00968_),
    .y(_00969_)
  );
  al_ao21ftf _05670_ (
    .a(g35),
    .b(\DFF_202.Q ),
    .c(_00969_),
    .y(\DFF_1159.D )
  );
  al_aoi21ftf _05671_ (
    .a(\DFF_948.Q ),
    .b(\DFF_595.Q ),
    .c(_00517_),
    .y(_00970_)
  );
  al_and3ftt _05672_ (
    .a(\DFF_1319.Q ),
    .b(\DFF_1270.Q ),
    .c(\DFF_1067.Q ),
    .y(_00971_)
  );
  al_and2 _05673_ (
    .a(\DFF_1148.Q ),
    .b(\DFF_717.Q ),
    .y(_00972_)
  );
  al_ao21ttf _05674_ (
    .a(_00972_),
    .b(_00524_),
    .c(\DFF_1110.Q ),
    .y(_00973_)
  );
  al_nand3ftt _05675_ (
    .a(_00971_),
    .b(_00970_),
    .c(_00973_),
    .y(_00974_)
  );
  al_and2ft _05676_ (
    .a(\DFF_1143.Q ),
    .b(\DFF_265.Q ),
    .y(_00975_)
  );
  al_aoi21ftf _05677_ (
    .a(\DFF_1389.Q ),
    .b(_00971_),
    .c(_00970_),
    .y(_00976_)
  );
  al_ao21ftf _05678_ (
    .a(_00971_),
    .b(\DFF_481.Q ),
    .c(_00976_),
    .y(_00977_)
  );
  al_or3fft _05679_ (
    .a(_00974_),
    .b(_00975_),
    .c(_00977_),
    .y(_00978_)
  );
  al_ao21 _05680_ (
    .a(_00975_),
    .b(_00974_),
    .c(\DFF_1025.Q ),
    .y(_00979_)
  );
  al_nand3 _05681_ (
    .a(g35),
    .b(_00979_),
    .c(_00978_),
    .y(_00980_)
  );
  al_ao21ftf _05682_ (
    .a(g35),
    .b(\DFF_959.Q ),
    .c(_00980_),
    .y(\DFF_1025.D )
  );
  al_or3ftt _05683_ (
    .a(_00503_),
    .b(\DFF_1272.Q ),
    .c(_00505_),
    .y(_00981_)
  );
  al_ao21ftf _05684_ (
    .a(_00503_),
    .b(_00505_),
    .c(_00981_),
    .y(_00982_)
  );
  al_mux2h _05685_ (
    .a(\DFF_530.Q ),
    .b(_00982_),
    .s(g35),
    .y(\DFF_1411.D )
  );
  al_and3 _05686_ (
    .a(\DFF_785.Q ),
    .b(\DFF_5.Q ),
    .c(_00404_),
    .y(_00983_)
  );
  al_nand2 _05687_ (
    .a(_00983_),
    .b(_00585_),
    .y(_00984_)
  );
  al_or3fft _05688_ (
    .a(\DFF_274.Q ),
    .b(g35),
    .c(_00984_),
    .y(_00985_)
  );
  al_or2 _05689_ (
    .a(\DFF_441.Q ),
    .b(g35),
    .y(_00986_)
  );
  al_and2ft _05690_ (
    .a(\DFF_274.Q ),
    .b(g35),
    .y(_00987_)
  );
  al_ao21ttf _05691_ (
    .a(_00983_),
    .b(_00585_),
    .c(_00987_),
    .y(_00988_)
  );
  al_and3 _05692_ (
    .a(_00986_),
    .b(_00988_),
    .c(_00985_),
    .y(\DFF_274.D )
  );
  al_oai21ftt _05693_ (
    .a(\DFF_358.Q ),
    .b(\DFF_718.Q ),
    .c(\DFF_63.Q ),
    .y(_00989_)
  );
  al_nand2 _05694_ (
    .a(\DFF_660.Q ),
    .b(\DFF_358.Q ),
    .y(_00990_)
  );
  al_nor2 _05695_ (
    .a(\DFF_63.Q ),
    .b(\DFF_660.Q ),
    .y(_00991_)
  );
  al_nand3ftt _05696_ (
    .a(_00991_),
    .b(_00989_),
    .c(_00990_),
    .y(_00992_)
  );
  al_nor2 _05697_ (
    .a(\DFF_660.Q ),
    .b(\DFF_358.Q ),
    .y(_00993_)
  );
  al_nand2ft _05698_ (
    .a(\DFF_718.Q ),
    .b(\DFF_63.Q ),
    .y(_00994_)
  );
  al_and2ft _05699_ (
    .a(\DFF_63.Q ),
    .b(\DFF_718.Q ),
    .y(_00995_)
  );
  al_and3fft _05700_ (
    .a(\DFF_807.Q ),
    .b(_00995_),
    .c(_00994_),
    .y(_00996_)
  );
  al_ao21ftf _05701_ (
    .a(_00993_),
    .b(_00990_),
    .c(_00996_),
    .y(_00997_)
  );
  al_aoi21 _05702_ (
    .a(_00992_),
    .b(_00997_),
    .c(g135),
    .y(_00998_)
  );
  al_and2ft _05703_ (
    .a(\DFF_331.Q ),
    .b(\DFF_43.Q ),
    .y(_00999_)
  );
  al_nor3fft _05704_ (
    .a(\DFF_674.Q ),
    .b(_00999_),
    .c(_00608_),
    .y(_01000_)
  );
  al_aoi21 _05705_ (
    .a(_01000_),
    .b(_00998_),
    .c(_00066_),
    .y(\DFF_1299.D )
  );
  al_and3ftt _05706_ (
    .a(\DFF_214.Q ),
    .b(\DFF_563.Q ),
    .c(\DFF_600.Q ),
    .y(_01001_)
  );
  al_nand3fft _05707_ (
    .a(\DFF_24.Q ),
    .b(\DFF_296.Q ),
    .c(_00718_),
    .y(_01002_)
  );
  al_ao21ftf _05708_ (
    .a(\DFF_24.Q ),
    .b(_00718_),
    .c(\DFF_296.Q ),
    .y(_01003_)
  );
  al_nand3 _05709_ (
    .a(_01001_),
    .b(_01002_),
    .c(_01003_),
    .y(_01004_)
  );
  al_nor2 _05710_ (
    .a(\DFF_98.Q ),
    .b(\DFF_580.Q ),
    .y(_01005_)
  );
  al_ao21 _05711_ (
    .a(_01001_),
    .b(_01005_),
    .c(\DFF_1290.Q ),
    .y(_01006_)
  );
  al_nand3 _05712_ (
    .a(g35),
    .b(_01006_),
    .c(_01004_),
    .y(_01007_)
  );
  al_ao21ftf _05713_ (
    .a(_00255_),
    .b(_00066_),
    .c(_01007_),
    .y(\DFF_1290.D )
  );
  al_nor2 _05714_ (
    .a(\DFF_726.Q ),
    .b(g35),
    .y(_01008_)
  );
  al_nand3fft _05715_ (
    .a(_00817_),
    .b(\DFF_1331.Q ),
    .c(_00563_),
    .y(_01009_)
  );
  al_or2 _05716_ (
    .a(\DFF_726.Q ),
    .b(\DFF_442.Q ),
    .y(_01010_)
  );
  al_nand2 _05717_ (
    .a(\DFF_726.Q ),
    .b(\DFF_442.Q ),
    .y(_01011_)
  );
  al_or3fft _05718_ (
    .a(_01010_),
    .b(_01011_),
    .c(_01009_),
    .y(_01012_)
  );
  al_aoi21 _05719_ (
    .a(\DFF_818.Q ),
    .b(_01009_),
    .c(_00066_),
    .y(_01013_)
  );
  al_aoi21 _05720_ (
    .a(_01012_),
    .b(_01013_),
    .c(_01008_),
    .y(\DFF_818.D )
  );
  al_and2 _05721_ (
    .a(\DFF_144.Q ),
    .b(g35),
    .y(\DFF_144.D )
  );
  al_nand3 _05722_ (
    .a(_00355_),
    .b(_00556_),
    .c(_00360_),
    .y(_01014_)
  );
  al_ao21 _05723_ (
    .a(\DFF_1408.Q ),
    .b(\DFF_245.Q ),
    .c(\DFF_199.Q ),
    .y(_01015_)
  );
  al_or2ft _05724_ (
    .a(g35),
    .b(_00378_),
    .y(_01016_)
  );
  al_nand3ftt _05725_ (
    .a(_01016_),
    .b(_01015_),
    .c(_01014_),
    .y(_01017_)
  );
  al_ao21ftf _05726_ (
    .a(g35),
    .b(\DFF_1408.Q ),
    .c(_01017_),
    .y(\DFF_199.D )
  );
  al_nand3 _05727_ (
    .a(_00441_),
    .b(_00975_),
    .c(_00563_),
    .y(_01018_)
  );
  al_ao21 _05728_ (
    .a(_00441_),
    .b(_00563_),
    .c(\DFF_425.Q ),
    .y(_01019_)
  );
  al_nand3 _05729_ (
    .a(g35),
    .b(_01018_),
    .c(_01019_),
    .y(_01020_)
  );
  al_ao21ftf _05730_ (
    .a(g35),
    .b(\DFF_1171.Q ),
    .c(_01020_),
    .y(\DFF_425.D )
  );
  al_or3 _05731_ (
    .a(\DFF_909.Q ),
    .b(\DFF_565.Q ),
    .c(\DFF_1234.Q ),
    .y(_01021_)
  );
  al_nor2 _05732_ (
    .a(\DFF_1416.Q ),
    .b(\DFF_1049.Q ),
    .y(_01022_)
  );
  al_nand3fft _05733_ (
    .a(\DFF_704.Q ),
    .b(\DFF_480.Q ),
    .c(_01022_),
    .y(_01023_)
  );
  al_or2 _05734_ (
    .a(\DFF_1389.Q ),
    .b(\DFF_1224.Q ),
    .y(_01024_)
  );
  al_oai21ttf _05735_ (
    .a(_01021_),
    .b(_01023_),
    .c(_01024_),
    .y(_01025_)
  );
  al_aoi21ftf _05736_ (
    .a(_00528_),
    .b(\DFF_1224.Q ),
    .c(_01025_),
    .y(_01026_)
  );
  al_mux2h _05737_ (
    .a(\DFF_858.Q ),
    .b(_01026_),
    .s(g35),
    .y(\DFF_1234.D )
  );
  al_aoi21 _05738_ (
    .a(\DFF_1408.Q ),
    .b(g35),
    .c(\DFF_245.Q ),
    .y(_01027_)
  );
  al_inv _05739_ (
    .a(\DFF_245.Q ),
    .y(_01028_)
  );
  al_ao21ftf _05740_ (
    .a(_01028_),
    .b(\DFF_1408.Q ),
    .c(_01014_),
    .y(_01029_)
  );
  al_aoi21 _05741_ (
    .a(g35),
    .b(_01029_),
    .c(_01027_),
    .y(\DFF_1408.D )
  );
  al_ao21 _05742_ (
    .a(_00759_),
    .b(_00758_),
    .c(_00066_),
    .y(_01030_)
  );
  al_mux2l _05743_ (
    .a(\DFF_933.Q ),
    .b(\DFF_1267.Q ),
    .s(_01030_),
    .y(\DFF_1267.D )
  );
  al_and2 _05744_ (
    .a(g35),
    .b(\DFF_507.Q ),
    .y(\DFF_507.D )
  );
  al_oai21ftf _05745_ (
    .a(\DFF_630.Q ),
    .b(\DFF_1396.Q ),
    .c(\DFF_539.Q ),
    .y(_01031_)
  );
  al_nand3ftt _05746_ (
    .a(\DFF_503.Q ),
    .b(g35),
    .c(_01031_),
    .y(_01032_)
  );
  al_ao21ftf _05747_ (
    .a(g35),
    .b(\DFF_1396.Q ),
    .c(_01032_),
    .y(\DFF_539.D )
  );
  al_and2ft _05748_ (
    .a(g35),
    .b(\DFF_915.Q ),
    .y(_01033_)
  );
  al_and3 _05749_ (
    .a(\DFF_1056.Q ),
    .b(\DFF_230.Q ),
    .c(\DFF_732.Q ),
    .y(_01034_)
  );
  al_and3fft _05750_ (
    .a(\DFF_1056.Q ),
    .b(\DFF_230.Q ),
    .c(\DFF_1279.Q ),
    .y(_01035_)
  );
  al_mux2h _05751_ (
    .a(_01035_),
    .b(_01034_),
    .s(\DFF_915.Q ),
    .y(_01036_)
  );
  al_mux2l _05752_ (
    .a(\DFF_1105.Q ),
    .b(\DFF_1147.Q ),
    .s(g84),
    .y(_01037_)
  );
  al_and2ft _05753_ (
    .a(\DFF_1257.Q ),
    .b(\DFF_732.Q ),
    .y(_01038_)
  );
  al_nand3 _05754_ (
    .a(\DFF_940.Q ),
    .b(_01037_),
    .c(_01038_),
    .y(_01039_)
  );
  al_and2 _05755_ (
    .a(\DFF_1279.Q ),
    .b(\DFF_1257.Q ),
    .y(_01040_)
  );
  al_nand3fft _05756_ (
    .a(\DFF_940.Q ),
    .b(_01037_),
    .c(_01040_),
    .y(_01041_)
  );
  al_and2 _05757_ (
    .a(_01039_),
    .b(_01041_),
    .y(_01042_)
  );
  al_ao21ftf _05758_ (
    .a(_01036_),
    .b(_01042_),
    .c(\DFF_850.Q ),
    .y(_01043_)
  );
  al_oa21ttf _05759_ (
    .a(\DFF_850.Q ),
    .b(_01036_),
    .c(_00066_),
    .y(_01044_)
  );
  al_ao21 _05760_ (
    .a(_01044_),
    .b(_01043_),
    .c(_01033_),
    .y(\DFF_850.D )
  );
  al_and2ft _05761_ (
    .a(\DFF_1408.Q ),
    .b(\DFF_199.Q ),
    .y(_01045_)
  );
  al_and2 _05762_ (
    .a(\DFF_120.Q ),
    .b(\DFF_27.Q ),
    .y(_01046_)
  );
  al_nand3 _05763_ (
    .a(_00499_),
    .b(_01045_),
    .c(_01046_),
    .y(_01047_)
  );
  al_ao21 _05764_ (
    .a(_01045_),
    .b(_01046_),
    .c(\DFF_102.Q ),
    .y(_01048_)
  );
  al_nand3 _05765_ (
    .a(g35),
    .b(_01048_),
    .c(_01047_),
    .y(_01049_)
  );
  al_ao21ftf _05766_ (
    .a(g35),
    .b(\DFF_1052.Q ),
    .c(_01049_),
    .y(\DFF_102.D )
  );
  al_and2 _05767_ (
    .a(\DFF_1161.Q ),
    .b(_00477_),
    .y(_01050_)
  );
  al_or3ftt _05768_ (
    .a(\DFF_237.Q ),
    .b(\DFF_1315.Q ),
    .c(\DFF_1108.Q ),
    .y(_01051_)
  );
  al_aoi21ttf _05769_ (
    .a(\DFF_1390.Q ),
    .b(_00479_),
    .c(_00478_),
    .y(_01052_)
  );
  al_ao21ftf _05770_ (
    .a(\DFF_1390.Q ),
    .b(_01051_),
    .c(_01052_),
    .y(_01053_)
  );
  al_nand2 _05771_ (
    .a(g35),
    .b(_01053_),
    .y(_01054_)
  );
  al_ao21ftt _05772_ (
    .a(_01050_),
    .b(\DFF_1250.Q ),
    .c(_01054_),
    .y(_01055_)
  );
  al_aoi21ftf _05773_ (
    .a(\DFF_238.Q ),
    .b(_00066_),
    .c(_01055_),
    .y(\DFF_1250.D )
  );
  al_and3ftt _05774_ (
    .a(_00019_),
    .b(_00575_),
    .c(_00544_),
    .y(_01056_)
  );
  al_and3ftt _05775_ (
    .a(_00451_),
    .b(_00604_),
    .c(_00422_),
    .y(_01057_)
  );
  al_aoi21ttf _05776_ (
    .a(\DFF_379.Q ),
    .b(_01057_),
    .c(_01056_),
    .y(_01058_)
  );
  al_oai21ftf _05777_ (
    .a(\DFF_1344.Q ),
    .b(\DFF_1064.Q ),
    .c(\DFF_794.Q ),
    .y(_01059_)
  );
  al_and2 _05778_ (
    .a(g35),
    .b(_01059_),
    .y(_01060_)
  );
  al_inv _05779_ (
    .a(\DFF_1064.Q ),
    .y(_01061_)
  );
  al_nor2 _05780_ (
    .a(\DFF_164.Q ),
    .b(g35),
    .y(_01062_)
  );
  al_nor2 _05781_ (
    .a(_00066_),
    .b(_01056_),
    .y(_01063_)
  );
  al_ao21 _05782_ (
    .a(_01061_),
    .b(_01063_),
    .c(_01062_),
    .y(_01064_)
  );
  al_aoi21 _05783_ (
    .a(_01060_),
    .b(_01058_),
    .c(_01064_),
    .y(\DFF_1064.D )
  );
  al_nor2 _05784_ (
    .a(g35),
    .b(\DFF_531.Q ),
    .y(_01065_)
  );
  al_and3 _05785_ (
    .a(g35),
    .b(_00516_),
    .c(_00718_),
    .y(_01066_)
  );
  al_aoi21 _05786_ (
    .a(_00044_),
    .b(_01066_),
    .c(_01065_),
    .y(\DFF_899.D )
  );
  al_nand3 _05787_ (
    .a(\DFF_563.Q ),
    .b(\DFF_214.Q ),
    .c(\DFF_675.Q ),
    .y(_01067_)
  );
  al_aoi21 _05788_ (
    .a(\DFF_416.Q ),
    .b(_01067_),
    .c(_00066_),
    .y(_01068_)
  );
  al_ao21ftf _05789_ (
    .a(_01067_),
    .b(\DFF_606.Q ),
    .c(_01068_),
    .y(_01069_)
  );
  al_aoi21ftf _05790_ (
    .a(\DFF_133.Q ),
    .b(_00066_),
    .c(_01069_),
    .y(\DFF_416.D )
  );
  al_and2ft _05791_ (
    .a(\DFF_199.Q ),
    .b(\DFF_1408.Q ),
    .y(_01070_)
  );
  al_nand3 _05792_ (
    .a(_00499_),
    .b(_01046_),
    .c(_01070_),
    .y(_01071_)
  );
  al_ao21 _05793_ (
    .a(_01070_),
    .b(_01046_),
    .c(\DFF_626.Q ),
    .y(_01072_)
  );
  al_nand3 _05794_ (
    .a(g35),
    .b(_01072_),
    .c(_01071_),
    .y(_01073_)
  );
  al_ao21ftf _05795_ (
    .a(g35),
    .b(\DFF_105.Q ),
    .c(_01073_),
    .y(\DFF_626.D )
  );
  al_oai21 _05796_ (
    .a(\DFF_754.Q ),
    .b(\DFF_323.Q ),
    .c(g35),
    .y(_01074_)
  );
  al_ao21ftf _05797_ (
    .a(g35),
    .b(\DFF_195.Q ),
    .c(_01074_),
    .y(\DFF_323.D )
  );
  al_nor2 _05798_ (
    .a(\DFF_1163.Q ),
    .b(\DFF_1213.Q ),
    .y(_01075_)
  );
  al_nand3fft _05799_ (
    .a(\DFF_322.Q ),
    .b(\DFF_814.Q ),
    .c(_01075_),
    .y(_01076_)
  );
  al_or3 _05800_ (
    .a(\DFF_1179.Q ),
    .b(\DFF_1418.Q ),
    .c(\DFF_1277.Q ),
    .y(_01077_)
  );
  al_or3 _05801_ (
    .a(\DFF_520.Q ),
    .b(_01077_),
    .c(_01076_),
    .y(_01078_)
  );
  al_nor2 _05802_ (
    .a(\DFF_499.Q ),
    .b(\DFF_1140.Q ),
    .y(_01079_)
  );
  al_and3fft _05803_ (
    .a(\DFF_1031.Q ),
    .b(\DFF_488.Q ),
    .c(_01079_),
    .y(_01080_)
  );
  al_or3 _05804_ (
    .a(\DFF_1071.Q ),
    .b(\DFF_444.Q ),
    .c(\DFF_825.Q ),
    .y(_01081_)
  );
  al_and3fft _05805_ (
    .a(\DFF_841.Q ),
    .b(_01081_),
    .c(_01080_),
    .y(_01082_)
  );
  al_nand3fft _05806_ (
    .a(\DFF_1182.Q ),
    .b(_01078_),
    .c(_01082_),
    .y(_01083_)
  );
  al_mux2h _05807_ (
    .a(\DFF_364.Q ),
    .b(_01083_),
    .s(g35),
    .y(\DFF_1182.D )
  );
  al_mux2h _05808_ (
    .a(\DFF_998.Q ),
    .b(_00898_),
    .s(g35),
    .y(\DFF_879.D )
  );
  al_and2ft _05809_ (
    .a(g35),
    .b(\DFF_1327.Q ),
    .y(_01084_)
  );
  al_inv _05810_ (
    .a(\DFF_690.Q ),
    .y(_01085_)
  );
  al_and3fft _05811_ (
    .a(\DFF_432.Q ),
    .b(\DFF_1341.Q ),
    .c(\DFF_366.Q ),
    .y(_01086_)
  );
  al_nand3fft _05812_ (
    .a(\DFF_386.Q ),
    .b(\DFF_1192.Q ),
    .c(_01086_),
    .y(_01087_)
  );
  al_or3ftt _05813_ (
    .a(_01085_),
    .b(\DFF_1327.Q ),
    .c(_01087_),
    .y(_01088_)
  );
  al_and3 _05814_ (
    .a(\DFF_1065.Q ),
    .b(\DFF_432.Q ),
    .c(\DFF_1341.Q ),
    .y(_01089_)
  );
  al_and3 _05815_ (
    .a(\DFF_386.Q ),
    .b(\DFF_1192.Q ),
    .c(_01089_),
    .y(_01090_)
  );
  al_nand2 _05816_ (
    .a(\DFF_1327.Q ),
    .b(\DFF_690.Q ),
    .y(_01091_)
  );
  al_ao21ftf _05817_ (
    .a(_01091_),
    .b(_01090_),
    .c(_01088_),
    .y(_01092_)
  );
  al_inv _05818_ (
    .a(\DFF_0.Q ),
    .y(_01093_)
  );
  al_nand2 _05819_ (
    .a(\DFF_1327.Q ),
    .b(\DFF_502.Q ),
    .y(_01094_)
  );
  al_mux2l _05820_ (
    .a(_01091_),
    .b(_01094_),
    .s(g84),
    .y(_01095_)
  );
  al_or3fft _05821_ (
    .a(_01093_),
    .b(\DFF_1065.Q ),
    .c(_01095_),
    .y(_01096_)
  );
  al_nand3fft _05822_ (
    .a(\DFF_1327.Q ),
    .b(\DFF_690.Q ),
    .c(g84),
    .y(_01097_)
  );
  al_nor2 _05823_ (
    .a(\DFF_1327.Q ),
    .b(\DFF_502.Q ),
    .y(_01098_)
  );
  al_ao21ftf _05824_ (
    .a(g84),
    .b(_01098_),
    .c(_01097_),
    .y(_01099_)
  );
  al_nand3 _05825_ (
    .a(\DFF_0.Q ),
    .b(\DFF_366.Q ),
    .c(_01099_),
    .y(_01100_)
  );
  al_and2 _05826_ (
    .a(_01100_),
    .b(_01096_),
    .y(_01101_)
  );
  al_ao21 _05827_ (
    .a(\DFF_502.Q ),
    .b(_01101_),
    .c(_01092_),
    .y(_01102_)
  );
  al_aoi21 _05828_ (
    .a(\DFF_502.Q ),
    .b(_01092_),
    .c(_00066_),
    .y(_01103_)
  );
  al_ao21 _05829_ (
    .a(_01103_),
    .b(_01102_),
    .c(_01084_),
    .y(\DFF_502.D )
  );
  al_and2ft _05830_ (
    .a(\DFF_584.Q ),
    .b(\DFF_410.Q ),
    .y(_01104_)
  );
  al_and2ft _05831_ (
    .a(\DFF_1068.Q ),
    .b(\DFF_1150.Q ),
    .y(_01105_)
  );
  al_nand3 _05832_ (
    .a(_00499_),
    .b(_01104_),
    .c(_01105_),
    .y(_01106_)
  );
  al_ao21 _05833_ (
    .a(_01104_),
    .b(_01105_),
    .c(\DFF_730.Q ),
    .y(_01107_)
  );
  al_nand3 _05834_ (
    .a(g35),
    .b(_01107_),
    .c(_01106_),
    .y(_01108_)
  );
  al_ao21ftf _05835_ (
    .a(g35),
    .b(\DFF_1032.Q ),
    .c(_01108_),
    .y(\DFF_730.D )
  );
  al_ao21ftf _05836_ (
    .a(\DFF_1161.Q ),
    .b(_00477_),
    .c(g35),
    .y(_01109_)
  );
  al_mux2l _05837_ (
    .a(\DFF_10.Q ),
    .b(\DFF_427.Q ),
    .s(_01109_),
    .y(\DFF_427.D )
  );
  al_and2 _05838_ (
    .a(\DFF_916.Q ),
    .b(g35),
    .y(\DFF_1316.D )
  );
  al_nand2 _05839_ (
    .a(g35),
    .b(_00642_),
    .y(_01110_)
  );
  al_mux2l _05840_ (
    .a(\DFF_1368.Q ),
    .b(\DFF_702.Q ),
    .s(_01110_),
    .y(\DFF_702.D )
  );
  al_nand3 _05841_ (
    .a(_00499_),
    .b(_00509_),
    .c(_01104_),
    .y(_01111_)
  );
  al_ao21 _05842_ (
    .a(_01104_),
    .b(_00509_),
    .c(\DFF_957.Q ),
    .y(_01112_)
  );
  al_nand3 _05843_ (
    .a(g35),
    .b(_01112_),
    .c(_01111_),
    .y(_01113_)
  );
  al_ao21ftf _05844_ (
    .a(g35),
    .b(\DFF_1174.Q ),
    .c(_01113_),
    .y(\DFF_957.D )
  );
  al_and2ft _05845_ (
    .a(\DFF_385.Q ),
    .b(\DFF_519.Q ),
    .y(_01114_)
  );
  al_nand3ftt _05846_ (
    .a(_00701_),
    .b(_00499_),
    .c(_01114_),
    .y(_01115_)
  );
  al_ao21ftt _05847_ (
    .a(_00701_),
    .b(_01114_),
    .c(\DFF_241.Q ),
    .y(_01116_)
  );
  al_nand3 _05848_ (
    .a(g35),
    .b(_01115_),
    .c(_01116_),
    .y(_01117_)
  );
  al_ao21ftf _05849_ (
    .a(g35),
    .b(\DFF_93.Q ),
    .c(_01117_),
    .y(\DFF_241.D )
  );
  al_and2ft _05850_ (
    .a(\DFF_703.Q ),
    .b(\DFF_586.Q ),
    .y(_01118_)
  );
  al_nand3 _05851_ (
    .a(\DFF_1298.Q ),
    .b(_00710_),
    .c(_01118_),
    .y(_01119_)
  );
  al_mux2h _05852_ (
    .a(\DFF_1239.Q ),
    .b(_01119_),
    .s(g35),
    .y(\DFF_513.D )
  );
  al_inv _05853_ (
    .a(\DFF_1122.Q ),
    .y(_01120_)
  );
  al_and2 _05854_ (
    .a(\DFF_563.Q ),
    .b(\DFF_214.Q ),
    .y(_01121_)
  );
  al_ao21 _05855_ (
    .a(_01121_),
    .b(_00346_),
    .c(_01120_),
    .y(_01122_)
  );
  al_nand3ftt _05856_ (
    .a(\DFF_445.Q ),
    .b(\DFF_941.Q ),
    .c(\DFF_507.Q ),
    .y(_01123_)
  );
  al_aoi21ftf _05857_ (
    .a(\DFF_1242.Q ),
    .b(\DFF_1046.Q ),
    .c(_00719_),
    .y(_01124_)
  );
  al_nand3 _05858_ (
    .a(_01123_),
    .b(_01124_),
    .c(_01122_),
    .y(_01125_)
  );
  al_nand3fft _05859_ (
    .a(\DFF_620.Q ),
    .b(\DFF_111.Q ),
    .c(_01125_),
    .y(_01126_)
  );
  al_nand2 _05860_ (
    .a(g35),
    .b(_01126_),
    .y(_01127_)
  );
  al_mux2l _05861_ (
    .a(\DFF_455.Q ),
    .b(\DFF_832.Q ),
    .s(_01127_),
    .y(\DFF_832.D )
  );
  al_inv _05862_ (
    .a(\DFF_620.Q ),
    .y(_01128_)
  );
  al_nand3 _05863_ (
    .a(\DFF_759.Q ),
    .b(_01128_),
    .c(_01125_),
    .y(_01129_)
  );
  al_ao21ftf _05864_ (
    .a(_01123_),
    .b(_00528_),
    .c(_01124_),
    .y(_01130_)
  );
  al_ao21ftt _05865_ (
    .a(_00723_),
    .b(_01123_),
    .c(_01130_),
    .y(_01131_)
  );
  al_aoi21ftf _05866_ (
    .a(\DFF_1422.Q ),
    .b(_01129_),
    .c(g35),
    .y(_01132_)
  );
  al_oai21 _05867_ (
    .a(_01129_),
    .b(_01131_),
    .c(_01132_),
    .y(_01133_)
  );
  al_ao21ftf _05868_ (
    .a(g35),
    .b(\DFF_973.Q ),
    .c(_01133_),
    .y(\DFF_1422.D )
  );
  al_nand3 _05869_ (
    .a(\DFF_1360.Q ),
    .b(g35),
    .c(_00361_),
    .y(_01134_)
  );
  al_or2 _05870_ (
    .a(\DFF_742.Q ),
    .b(g35),
    .y(_01135_)
  );
  al_or3ftt _05871_ (
    .a(g35),
    .b(\DFF_1360.Q ),
    .c(_00361_),
    .y(_01136_)
  );
  al_and3 _05872_ (
    .a(_01135_),
    .b(_01134_),
    .c(_01136_),
    .y(\DFF_1360.D )
  );
  al_oai21ftf _05873_ (
    .a(\DFF_85.Q ),
    .b(\DFF_235.Q ),
    .c(\DFF_396.Q ),
    .y(_01137_)
  );
  al_nand3ftt _05874_ (
    .a(\DFF_376.Q ),
    .b(g35),
    .c(_01137_),
    .y(_01138_)
  );
  al_ao21ftf _05875_ (
    .a(g35),
    .b(\DFF_235.Q ),
    .c(_01138_),
    .y(\DFF_396.D )
  );
  al_nand3 _05876_ (
    .a(_00513_),
    .b(\DFF_1010.Q ),
    .c(_00526_),
    .y(_01139_)
  );
  al_aoi21ftf _05877_ (
    .a(\DFF_1247.Q ),
    .b(_01139_),
    .c(g35),
    .y(_01140_)
  );
  al_ao21ftf _05878_ (
    .a(_01139_),
    .b(_00530_),
    .c(_01140_),
    .y(_01141_)
  );
  al_ao21ftf _05879_ (
    .a(g35),
    .b(\DFF_65.Q ),
    .c(_01141_),
    .y(\DFF_1247.D )
  );
  al_nor2 _05880_ (
    .a(\DFF_1192.Q ),
    .b(g35),
    .y(_01142_)
  );
  al_mux2h _05881_ (
    .a(_01086_),
    .b(_01089_),
    .s(\DFF_1192.Q ),
    .y(_01143_)
  );
  al_nand3ftt _05882_ (
    .a(_01143_),
    .b(\DFF_386.Q ),
    .c(_01101_),
    .y(_01144_)
  );
  al_aoi21ftf _05883_ (
    .a(\DFF_386.Q ),
    .b(_01143_),
    .c(g35),
    .y(_01145_)
  );
  al_aoi21 _05884_ (
    .a(_01145_),
    .b(_01144_),
    .c(_01142_),
    .y(\DFF_386.D )
  );
  al_aoi21ftf _05885_ (
    .a(\DFF_1242.Q ),
    .b(\DFF_1136.Q ),
    .c(_00719_),
    .y(_01146_)
  );
  al_and3 _05886_ (
    .a(\DFF_941.Q ),
    .b(\DFF_445.Q ),
    .c(\DFF_507.Q ),
    .y(_01147_)
  );
  al_nor2 _05887_ (
    .a(\DFF_563.Q ),
    .b(\DFF_214.Q ),
    .y(_01148_)
  );
  al_ao21ttf _05888_ (
    .a(_01148_),
    .b(_00346_),
    .c(\DFF_295.Q ),
    .y(_01149_)
  );
  al_nand3ftt _05889_ (
    .a(_01147_),
    .b(_01146_),
    .c(_01149_),
    .y(_01150_)
  );
  al_nand2ft _05890_ (
    .a(\DFF_1413.Q ),
    .b(\DFF_671.Q ),
    .y(_01151_)
  );
  al_aoi21ftf _05891_ (
    .a(\DFF_1389.Q ),
    .b(_01147_),
    .c(_01146_),
    .y(_01152_)
  );
  al_ao21ftf _05892_ (
    .a(_01147_),
    .b(_00723_),
    .c(_01152_),
    .y(_01153_)
  );
  al_and3fft _05893_ (
    .a(_01151_),
    .b(_01153_),
    .c(_01150_),
    .y(_01154_)
  );
  al_ao21ftt _05894_ (
    .a(_01151_),
    .b(_01150_),
    .c(\DFF_641.Q ),
    .y(_01155_)
  );
  al_or3fft _05895_ (
    .a(g35),
    .b(_01155_),
    .c(_01154_),
    .y(_01156_)
  );
  al_ao21ftf _05896_ (
    .a(g35),
    .b(\DFF_809.Q ),
    .c(_01156_),
    .y(\DFF_641.D )
  );
  al_or3 _05897_ (
    .a(\DFF_1374.Q ),
    .b(\DFF_807.Q ),
    .c(\DFF_1173.Q ),
    .y(_01157_)
  );
  al_and3fft _05898_ (
    .a(\DFF_718.Q ),
    .b(_01157_),
    .c(_00991_),
    .y(_01158_)
  );
  al_and3ftt _05899_ (
    .a(\DFF_358.Q ),
    .b(\DFF_853.Q ),
    .c(g35),
    .y(_01159_)
  );
  al_nor3fft _05900_ (
    .a(\DFF_674.Q ),
    .b(_00999_),
    .c(_00747_),
    .y(_01160_)
  );
  al_nand3 _05901_ (
    .a(_01159_),
    .b(_01160_),
    .c(_01158_),
    .y(_01161_)
  );
  al_ao21ftf _05902_ (
    .a(g35),
    .b(\DFF_1374.Q ),
    .c(_01161_),
    .y(\DFF_934.D )
  );
  al_nand3ftt _05903_ (
    .a(\DFF_1204.Q ),
    .b(\DFF_527.Q ),
    .c(g35),
    .y(_01162_)
  );
  al_ao21ftf _05904_ (
    .a(g35),
    .b(\DFF_434.Q ),
    .c(_01162_),
    .y(\DFF_1204.D )
  );
  al_nor3ftt _05905_ (
    .a(\DFF_918.Q ),
    .b(_00499_),
    .c(_00369_),
    .y(_01163_)
  );
  al_oa21ftt _05906_ (
    .a(\DFF_918.Q ),
    .b(_00369_),
    .c(_00499_),
    .y(_01164_)
  );
  al_nor3ftt _05907_ (
    .a(g35),
    .b(_01163_),
    .c(_01164_),
    .y(\DFF_918.D )
  );
  al_oa21ttf _05908_ (
    .a(\DFF_366.Q ),
    .b(\DFF_1065.Q ),
    .c(\DFF_1341.Q ),
    .y(_01165_)
  );
  al_nand3 _05909_ (
    .a(_01165_),
    .b(_01100_),
    .c(_01096_),
    .y(_01166_)
  );
  al_nand3fft _05910_ (
    .a(\DFF_366.Q ),
    .b(\DFF_1065.Q ),
    .c(\DFF_1341.Q ),
    .y(_01167_)
  );
  al_nand3 _05911_ (
    .a(g35),
    .b(_01167_),
    .c(_01166_),
    .y(_01168_)
  );
  al_aoi21ftf _05912_ (
    .a(\DFF_366.Q ),
    .b(_00066_),
    .c(_01168_),
    .y(\DFF_1341.D )
  );
  al_and2 _05913_ (
    .a(\DFF_657.Q ),
    .b(g35),
    .y(\DFF_657.D )
  );
  al_and2ft _05914_ (
    .a(\DFF_925.Q ),
    .b(\DFF_653.Q ),
    .y(_01169_)
  );
  al_and2ft _05915_ (
    .a(\DFF_20.Q ),
    .b(\DFF_916.Q ),
    .y(_01170_)
  );
  al_nand3 _05916_ (
    .a(_00499_),
    .b(_01169_),
    .c(_01170_),
    .y(_01171_)
  );
  al_ao21 _05917_ (
    .a(_01169_),
    .b(_01170_),
    .c(\DFF_59.Q ),
    .y(_01172_)
  );
  al_nand3 _05918_ (
    .a(g35),
    .b(_01172_),
    .c(_01171_),
    .y(_01173_)
  );
  al_ao21ftf _05919_ (
    .a(g35),
    .b(\DFF_634.Q ),
    .c(_01173_),
    .y(\DFF_59.D )
  );
  al_and2 _05920_ (
    .a(g35),
    .b(g6745),
    .y(\DFF_760.D )
  );
  al_ao21 _05921_ (
    .a(\DFF_1161.Q ),
    .b(_00477_),
    .c(_00066_),
    .y(_01174_)
  );
  al_mux2l _05922_ (
    .a(\DFF_719.Q ),
    .b(\DFF_23.Q ),
    .s(_01174_),
    .y(\DFF_23.D )
  );
  al_oa21ftt _05923_ (
    .a(\DFF_1081.Q ),
    .b(\DFF_256.Q ),
    .c(g35),
    .y(_01175_)
  );
  al_aoi21ttf _05924_ (
    .a(\DFF_142.Q ),
    .b(\DFF_21.Q ),
    .c(_00946_),
    .y(_01176_)
  );
  al_and3 _05925_ (
    .a(_00944_),
    .b(_01176_),
    .c(_00481_),
    .y(_01177_)
  );
  al_and3 _05926_ (
    .a(\DFF_876.Q ),
    .b(_00948_),
    .c(_01177_),
    .y(_01178_)
  );
  al_and3 _05927_ (
    .a(\DFF_175.Q ),
    .b(_00943_),
    .c(_01178_),
    .y(_01179_)
  );
  al_or3fft _05928_ (
    .a(\DFF_328.Q ),
    .b(_01175_),
    .c(_01179_),
    .y(_01180_)
  );
  al_nand2ft _05929_ (
    .a(g35),
    .b(\DFF_28.Q ),
    .y(_01181_)
  );
  al_nand3fft _05930_ (
    .a(\DFF_328.Q ),
    .b(_00066_),
    .c(_01179_),
    .y(_01182_)
  );
  al_nand3 _05931_ (
    .a(_01181_),
    .b(_01182_),
    .c(_01180_),
    .y(\DFF_328.D )
  );
  al_nand2ft _05932_ (
    .a(\DFF_7.Q ),
    .b(\DFF_109.Q ),
    .y(_01183_)
  );
  al_oa21ftt _05933_ (
    .a(\DFF_752.Q ),
    .b(\DFF_109.Q ),
    .c(\DFF_654.Q ),
    .y(_01184_)
  );
  al_and3 _05934_ (
    .a(\DFF_728.Q ),
    .b(\DFF_88.Q ),
    .c(_01184_),
    .y(_01185_)
  );
  al_nand3 _05935_ (
    .a(\DFF_506.Q ),
    .b(\DFF_560.Q ),
    .c(_01185_),
    .y(_01186_)
  );
  al_oa21ftt _05936_ (
    .a(\DFF_109.Q ),
    .b(\DFF_7.Q ),
    .c(\DFF_863.Q ),
    .y(_01187_)
  );
  al_and3fft _05937_ (
    .a(_00282_),
    .b(_01186_),
    .c(_01187_),
    .y(_01188_)
  );
  al_ao21ftt _05938_ (
    .a(_00065_),
    .b(_01183_),
    .c(_01188_),
    .y(_01189_)
  );
  al_and3 _05939_ (
    .a(\DFF_162.Q ),
    .b(_01183_),
    .c(_01188_),
    .y(_01190_)
  );
  al_oai21ftf _05940_ (
    .a(_01189_),
    .b(_01190_),
    .c(_00066_),
    .y(_01191_)
  );
  al_aoi21ftf _05941_ (
    .a(\DFF_1235.Q ),
    .b(_00066_),
    .c(_01191_),
    .y(\DFF_162.D )
  );
  al_or3ftt _05942_ (
    .a(_00305_),
    .b(\DFF_154.Q ),
    .c(_00306_),
    .y(_01192_)
  );
  al_or3fft _05943_ (
    .a(\DFF_1324.Q ),
    .b(\DFF_891.Q ),
    .c(_01192_),
    .y(_01193_)
  );
  al_mux2l _05944_ (
    .a(\DFF_1083.Q ),
    .b(\DFF_1230.Q ),
    .s(_01193_),
    .y(_01194_)
  );
  al_mux2h _05945_ (
    .a(\DFF_1187.Q ),
    .b(_01194_),
    .s(g35),
    .y(\DFF_1083.D )
  );
  al_nand3fft _05946_ (
    .a(\DFF_1413.Q ),
    .b(\DFF_996.Q ),
    .c(_01150_),
    .y(_01195_)
  );
  al_nand2 _05947_ (
    .a(\DFF_888.Q ),
    .b(\DFF_1086.Q ),
    .y(_01196_)
  );
  al_nor2 _05948_ (
    .a(\DFF_888.Q ),
    .b(\DFF_1086.Q ),
    .y(_01197_)
  );
  al_nand2ft _05949_ (
    .a(_01197_),
    .b(_01196_),
    .y(_01198_)
  );
  al_mux2l _05950_ (
    .a(\DFF_322.Q ),
    .b(_01198_),
    .s(_01195_),
    .y(_01199_)
  );
  al_mux2h _05951_ (
    .a(\DFF_1086.Q ),
    .b(_01199_),
    .s(g35),
    .y(\DFF_322.D )
  );
  al_oa21ttf _05952_ (
    .a(\DFF_1279.Q ),
    .b(\DFF_732.Q ),
    .c(\DFF_230.Q ),
    .y(_01200_)
  );
  al_nand3 _05953_ (
    .a(_01200_),
    .b(_01039_),
    .c(_01041_),
    .y(_01201_)
  );
  al_or3ftt _05954_ (
    .a(\DFF_230.Q ),
    .b(\DFF_1279.Q ),
    .c(\DFF_732.Q ),
    .y(_01202_)
  );
  al_nand3 _05955_ (
    .a(g35),
    .b(_01202_),
    .c(_01201_),
    .y(_01203_)
  );
  al_aoi21ftf _05956_ (
    .a(\DFF_1279.Q ),
    .b(_00066_),
    .c(_01203_),
    .y(\DFF_230.D )
  );
  al_and2ft _05957_ (
    .a(g35),
    .b(\DFF_1227.Q ),
    .y(_01204_)
  );
  al_ao21ftf _05958_ (
    .a(\DFF_1227.Q ),
    .b(_00827_),
    .c(_00831_),
    .y(_01205_)
  );
  al_ao21ftt _05959_ (
    .a(\DFF_316.Q ),
    .b(_00827_),
    .c(_01205_),
    .y(_01206_)
  );
  al_aoi21ftf _05960_ (
    .a(\DFF_316.Q ),
    .b(_01205_),
    .c(g35),
    .y(_01207_)
  );
  al_ao21 _05961_ (
    .a(_01206_),
    .b(_01207_),
    .c(_01204_),
    .y(\DFF_316.D )
  );
  al_and2 _05962_ (
    .a(\DFF_724.Q ),
    .b(g35),
    .y(_01208_)
  );
  al_nand3fft _05963_ (
    .a(\DFF_439.Q ),
    .b(g73),
    .c(g72),
    .y(_01209_)
  );
  al_mux2l _05964_ (
    .a(_01209_),
    .b(\DFF_56.Q ),
    .s(_01208_),
    .y(\DFF_816.D )
  );
  al_and3fft _05965_ (
    .a(\DFF_563.Q ),
    .b(\DFF_214.Q ),
    .c(\DFF_600.Q ),
    .y(_01210_)
  );
  al_and2ft _05966_ (
    .a(\DFF_1094.Q ),
    .b(\DFF_98.Q ),
    .y(_01211_)
  );
  al_and3 _05967_ (
    .a(\DFF_1274.Q ),
    .b(_01210_),
    .c(_01211_),
    .y(_01212_)
  );
  al_or2 _05968_ (
    .a(_00113_),
    .b(_01212_),
    .y(_01213_)
  );
  al_nand2 _05969_ (
    .a(_00113_),
    .b(_01212_),
    .y(_01214_)
  );
  al_nand3 _05970_ (
    .a(g35),
    .b(_01214_),
    .c(_01213_),
    .y(_01215_)
  );
  al_aoi21ftf _05971_ (
    .a(\DFF_1274.Q ),
    .b(_00066_),
    .c(_01215_),
    .y(\DFF_1136.D )
  );
  al_and2ft _05972_ (
    .a(g35),
    .b(\DFF_1312.Q ),
    .y(_01216_)
  );
  al_nand2 _05973_ (
    .a(\DFF_1312.Q ),
    .b(_00766_),
    .y(_01217_)
  );
  al_aoi21ftf _05974_ (
    .a(\DFF_536.Q ),
    .b(_01217_),
    .c(g35),
    .y(_01218_)
  );
  al_nand3 _05975_ (
    .a(_00587_),
    .b(_00766_),
    .c(_00401_),
    .y(_01219_)
  );
  al_aoi21ftf _05976_ (
    .a(_01217_),
    .b(\DFF_536.Q ),
    .c(_01219_),
    .y(_01220_)
  );
  al_ao21 _05977_ (
    .a(_01218_),
    .b(_01220_),
    .c(_01216_),
    .y(\DFF_536.D )
  );
  al_nand3fft _05978_ (
    .a(\DFF_1191.Q ),
    .b(\DFF_178.Q ),
    .c(_00342_),
    .y(_01221_)
  );
  al_or2ft _05979_ (
    .a(\DFF_417.Q ),
    .b(_01221_),
    .y(_01222_)
  );
  al_ao21 _05980_ (
    .a(_00462_),
    .b(_01222_),
    .c(_00066_),
    .y(_01223_)
  );
  al_nand2 _05981_ (
    .a(\DFF_894.Q ),
    .b(\DFF_849.Q ),
    .y(_01224_)
  );
  al_oai21ftf _05982_ (
    .a(_00461_),
    .b(_01224_),
    .c(\DFF_1311.Q ),
    .y(_01225_)
  );
  al_oa21ftf _05983_ (
    .a(\DFF_417.Q ),
    .b(_01221_),
    .c(_00066_),
    .y(_01226_)
  );
  al_ao21ttf _05984_ (
    .a(_01221_),
    .b(_01225_),
    .c(_01226_),
    .y(_01227_)
  );
  al_aoi21ftf _05985_ (
    .a(\DFF_747.Q ),
    .b(_01223_),
    .c(_01227_),
    .y(\DFF_1311.D )
  );
  al_nor2 _05986_ (
    .a(\DFF_844.Q ),
    .b(g35),
    .y(_01228_)
  );
  al_oa21ftt _05987_ (
    .a(\DFF_109.Q ),
    .b(\DFF_7.Q ),
    .c(\DFF_844.Q ),
    .y(_01229_)
  );
  al_oa21ftt _05988_ (
    .a(\DFF_109.Q ),
    .b(\DFF_7.Q ),
    .c(\DFF_89.Q ),
    .y(_01230_)
  );
  al_and2 _05989_ (
    .a(\DFF_506.Q ),
    .b(_01185_),
    .y(_01231_)
  );
  al_and3 _05990_ (
    .a(\DFF_560.Q ),
    .b(_01183_),
    .c(_01231_),
    .y(_01232_)
  );
  al_and3 _05991_ (
    .a(\DFF_863.Q ),
    .b(\DFF_1235.Q ),
    .c(_01232_),
    .y(_01233_)
  );
  al_and3 _05992_ (
    .a(\DFF_162.Q ),
    .b(_01183_),
    .c(_01233_),
    .y(_01234_)
  );
  al_and3 _05993_ (
    .a(\DFF_874.Q ),
    .b(\DFF_1090.Q ),
    .c(_01234_),
    .y(_01235_)
  );
  al_and3 _05994_ (
    .a(\DFF_966.Q ),
    .b(_01230_),
    .c(_01235_),
    .y(_01236_)
  );
  al_nand3 _05995_ (
    .a(\DFF_812.Q ),
    .b(\DFF_751.Q ),
    .c(_01236_),
    .y(_01237_)
  );
  al_or3fft _05996_ (
    .a(\DFF_119.Q ),
    .b(_01229_),
    .c(_01237_),
    .y(_01238_)
  );
  al_nand3 _05997_ (
    .a(\DFF_338.Q ),
    .b(_01183_),
    .c(_01238_),
    .y(_01239_)
  );
  al_oa21ttf _05998_ (
    .a(\DFF_338.Q ),
    .b(_01238_),
    .c(_00066_),
    .y(_01240_)
  );
  al_aoi21 _05999_ (
    .a(_01239_),
    .b(_01240_),
    .c(_01228_),
    .y(\DFF_338.D )
  );
  al_nand3 _06000_ (
    .a(_00499_),
    .b(_00592_),
    .c(_01114_),
    .y(_01241_)
  );
  al_ao21 _06001_ (
    .a(_00592_),
    .b(_01114_),
    .c(\DFF_1085.Q ),
    .y(_01242_)
  );
  al_nand3 _06002_ (
    .a(g35),
    .b(_01242_),
    .c(_01241_),
    .y(_01243_)
  );
  al_ao21ftf _06003_ (
    .a(g35),
    .b(\DFF_920.Q ),
    .c(_01243_),
    .y(\DFF_1085.D )
  );
  al_or2 _06004_ (
    .a(_00474_),
    .b(_00490_),
    .y(_01244_)
  );
  al_ao21ttf _06005_ (
    .a(\DFF_409.Q ),
    .b(_00488_),
    .c(_01244_),
    .y(_01245_)
  );
  al_nand3fft _06006_ (
    .a(_00066_),
    .b(_00491_),
    .c(_01245_),
    .y(_01246_)
  );
  al_ao21ftf _06007_ (
    .a(g35),
    .b(\DFF_582.Q ),
    .c(_01246_),
    .y(\DFF_409.D )
  );
  al_mux2l _06008_ (
    .a(\DFF_357.Q ),
    .b(\DFF_1103.Q ),
    .s(g35),
    .y(\DFF_339.D )
  );
  al_mux2h _06009_ (
    .a(\DFF_0.Q ),
    .b(_01100_),
    .s(g35),
    .y(\DFF_1124.D )
  );
  al_and2ft _06010_ (
    .a(\DFF_1190.Q ),
    .b(g35),
    .y(\DFF_1190.D )
  );
  al_and3 _06011_ (
    .a(\DFF_794.Q ),
    .b(\DFF_246.Q ),
    .c(\DFF_1064.Q ),
    .y(_01247_)
  );
  al_and3fft _06012_ (
    .a(\DFF_794.Q ),
    .b(\DFF_1064.Q ),
    .c(\DFF_1180.Q ),
    .y(_01248_)
  );
  al_nand3ftt _06013_ (
    .a(\DFF_1064.Q ),
    .b(\DFF_1344.Q ),
    .c(\DFF_32.Q ),
    .y(_01249_)
  );
  al_nand3ftt _06014_ (
    .a(\DFF_1344.Q ),
    .b(\DFF_564.Q ),
    .c(\DFF_794.Q ),
    .y(_01250_)
  );
  al_and3ftt _06015_ (
    .a(\DFF_1344.Q ),
    .b(\DFF_735.Q ),
    .c(\DFF_1064.Q ),
    .y(_01251_)
  );
  al_aoi21 _06016_ (
    .a(\DFF_864.Q ),
    .b(g25167),
    .c(_01251_),
    .y(_01252_)
  );
  al_and3 _06017_ (
    .a(_01249_),
    .b(_01250_),
    .c(_01252_),
    .y(_01253_)
  );
  al_nand3fft _06018_ (
    .a(_01247_),
    .b(_01248_),
    .c(_01253_),
    .y(_01254_)
  );
  al_mux2h _06019_ (
    .a(\DFF_1069.Q ),
    .b(_01254_),
    .s(_01056_),
    .y(_01255_)
  );
  al_mux2h _06020_ (
    .a(\DFF_794.Q ),
    .b(_01255_),
    .s(g35),
    .y(\DFF_1069.D )
  );
  al_nand2ft _06021_ (
    .a(\DFF_879.Q ),
    .b(\DFF_596.Q ),
    .y(_01256_)
  );
  al_and3fft _06022_ (
    .a(\DFF_1287.Q ),
    .b(\DFF_821.Q ),
    .c(\DFF_596.Q ),
    .y(_01257_)
  );
  al_oai21ftf _06023_ (
    .a(\DFF_1287.Q ),
    .b(_01256_),
    .c(_01257_),
    .y(_01258_)
  );
  al_mux2h _06024_ (
    .a(\DFF_596.Q ),
    .b(_01258_),
    .s(g35),
    .y(\DFF_1142.D )
  );
  al_inv _06025_ (
    .a(\DFF_774.Q ),
    .y(_01259_)
  );
  al_and3ftt _06026_ (
    .a(\DFF_717.Q ),
    .b(\DFF_1148.Q ),
    .c(\DFF_327.Q ),
    .y(_01260_)
  );
  al_and2ft _06027_ (
    .a(\DFF_167.Q ),
    .b(\DFF_182.Q ),
    .y(_01261_)
  );
  al_and3 _06028_ (
    .a(\DFF_169.Q ),
    .b(_01260_),
    .c(_01261_),
    .y(_01262_)
  );
  al_or2 _06029_ (
    .a(_01259_),
    .b(_01262_),
    .y(_01263_)
  );
  al_nand2 _06030_ (
    .a(_01259_),
    .b(_01262_),
    .y(_01264_)
  );
  al_nand3 _06031_ (
    .a(g35),
    .b(_01264_),
    .c(_01263_),
    .y(_01265_)
  );
  al_aoi21ftf _06032_ (
    .a(\DFF_169.Q ),
    .b(_00066_),
    .c(_01265_),
    .y(\DFF_774.D )
  );
  al_and2ft _06033_ (
    .a(\DFF_784.Q ),
    .b(\DFF_776.Q ),
    .y(_01266_)
  );
  al_nand3 _06034_ (
    .a(_00499_),
    .b(_00597_),
    .c(_01266_),
    .y(_01267_)
  );
  al_ao21 _06035_ (
    .a(_00597_),
    .b(_01266_),
    .c(\DFF_868.Q ),
    .y(_01268_)
  );
  al_nand3 _06036_ (
    .a(g35),
    .b(_01268_),
    .c(_01267_),
    .y(_01269_)
  );
  al_ao21ftf _06037_ (
    .a(g35),
    .b(\DFF_1128.Q ),
    .c(_01269_),
    .y(\DFF_868.D )
  );
  al_inv _06038_ (
    .a(\DFF_473.Q ),
    .y(_01270_)
  );
  al_nand3 _06039_ (
    .a(_01270_),
    .b(_00596_),
    .c(_00734_),
    .y(_01271_)
  );
  al_ao21ftf _06040_ (
    .a(g35),
    .b(\DFF_776.Q ),
    .c(_01271_),
    .y(\DFF_473.D )
  );
  al_and2 _06041_ (
    .a(_00542_),
    .b(_00549_),
    .y(_01272_)
  );
  al_oa21ftf _06042_ (
    .a(\DFF_763.Q ),
    .b(_00604_),
    .c(_00698_),
    .y(_01273_)
  );
  al_mux2h _06043_ (
    .a(\DFF_1112.Q ),
    .b(_01273_),
    .s(_01272_),
    .y(_01274_)
  );
  al_mux2h _06044_ (
    .a(\DFF_284.Q ),
    .b(_01274_),
    .s(g35),
    .y(\DFF_1112.D )
  );
  al_nand3ftt _06045_ (
    .a(\DFF_910.Q ),
    .b(\DFF_575.Q ),
    .c(\DFF_289.Q ),
    .y(_01275_)
  );
  al_aoi21ftf _06046_ (
    .a(\DFF_172.Q ),
    .b(_01275_),
    .c(g35),
    .y(_01276_)
  );
  al_ao21ftf _06047_ (
    .a(_01275_),
    .b(_00499_),
    .c(_01276_),
    .y(_01277_)
  );
  al_ao21ftf _06048_ (
    .a(g35),
    .b(\DFF_219.Q ),
    .c(_01277_),
    .y(\DFF_172.D )
  );
  al_aoi21ftf _06049_ (
    .a(\DFF_948.Q ),
    .b(\DFF_774.Q ),
    .c(_00517_),
    .y(_01278_)
  );
  al_nand3fft _06050_ (
    .a(\DFF_1270.Q ),
    .b(\DFF_1319.Q ),
    .c(\DFF_1067.Q ),
    .y(_01279_)
  );
  al_and2ft _06051_ (
    .a(\DFF_717.Q ),
    .b(\DFF_1148.Q ),
    .y(_01280_)
  );
  al_ao21ttf _06052_ (
    .a(_01280_),
    .b(_00524_),
    .c(\DFF_422.Q ),
    .y(_01281_)
  );
  al_nand3 _06053_ (
    .a(_01279_),
    .b(_01278_),
    .c(_01281_),
    .y(_01282_)
  );
  al_aoi21ftf _06054_ (
    .a(_01279_),
    .b(_00528_),
    .c(_01278_),
    .y(_01283_)
  );
  al_ao21ttf _06055_ (
    .a(\DFF_481.Q ),
    .b(_01279_),
    .c(_01283_),
    .y(_01284_)
  );
  al_or3fft _06056_ (
    .a(_00877_),
    .b(_01282_),
    .c(_01284_),
    .y(_01285_)
  );
  al_ao21 _06057_ (
    .a(_00877_),
    .b(_01282_),
    .c(\DFF_204.Q ),
    .y(_01286_)
  );
  al_nand3 _06058_ (
    .a(g35),
    .b(_01286_),
    .c(_01285_),
    .y(_01287_)
  );
  al_ao21ftf _06059_ (
    .a(g35),
    .b(\DFF_1135.Q ),
    .c(_01287_),
    .y(\DFF_204.D )
  );
  al_aoi21 _06060_ (
    .a(\DFF_248.Q ),
    .b(g35),
    .c(\DFF_883.Q ),
    .y(_01288_)
  );
  al_oa21ftt _06061_ (
    .a(g35),
    .b(\DFF_883.Q ),
    .c(\DFF_248.Q ),
    .y(_01289_)
  );
  al_aoi21 _06062_ (
    .a(g35),
    .b(_01289_),
    .c(_01288_),
    .y(\DFF_248.D )
  );
  al_nand3ftt _06063_ (
    .a(\DFF_575.Q ),
    .b(\DFF_289.Q ),
    .c(\DFF_910.Q ),
    .y(_01290_)
  );
  al_aoi21ftf _06064_ (
    .a(\DFF_84.Q ),
    .b(_01290_),
    .c(g35),
    .y(_01291_)
  );
  al_ao21ftf _06065_ (
    .a(_01290_),
    .b(_00499_),
    .c(_01291_),
    .y(_01292_)
  );
  al_ao21ftf _06066_ (
    .a(g35),
    .b(\DFF_44.Q ),
    .c(_01292_),
    .y(\DFF_84.D )
  );
  al_and2ft _06067_ (
    .a(g35),
    .b(\DFF_97.Q ),
    .y(_01293_)
  );
  al_inv _06068_ (
    .a(\DFF_712.Q ),
    .y(_01294_)
  );
  al_nand3fft _06069_ (
    .a(\DFF_49.Q ),
    .b(\DFF_40.Q ),
    .c(_00901_),
    .y(_01295_)
  );
  al_nand3 _06070_ (
    .a(\DFF_49.Q ),
    .b(\DFF_40.Q ),
    .c(_00900_),
    .y(_01296_)
  );
  al_mux2l _06071_ (
    .a(_01295_),
    .b(_01296_),
    .s(_01294_),
    .y(_01297_)
  );
  al_aoi21ftt _06072_ (
    .a(_00896_),
    .b(_00892_),
    .c(_01297_),
    .y(_01298_)
  );
  al_ao21ftf _06073_ (
    .a(_00895_),
    .b(_00891_),
    .c(_01298_),
    .y(_01299_)
  );
  al_ao21ftf _06074_ (
    .a(_00889_),
    .b(_00898_),
    .c(_01299_),
    .y(_01300_)
  );
  al_oa21ftf _06075_ (
    .a(\DFF_998.Q ),
    .b(_01299_),
    .c(_00066_),
    .y(_01301_)
  );
  al_ao21 _06076_ (
    .a(_01300_),
    .b(_01301_),
    .c(_01293_),
    .y(\DFF_998.D )
  );
  al_or2 _06077_ (
    .a(\DFF_1227.Q ),
    .b(_00831_),
    .y(_01302_)
  );
  al_nand3 _06078_ (
    .a(g35),
    .b(_01205_),
    .c(_01302_),
    .y(_01303_)
  );
  al_ao21ftf _06079_ (
    .a(g35),
    .b(\DFF_577.Q ),
    .c(_01303_),
    .y(\DFF_1227.D )
  );
  al_mux2l _06080_ (
    .a(\DFF_608.Q ),
    .b(\DFF_236.Q ),
    .s(g35),
    .y(\DFF_608.D )
  );
  al_oai21ftt _06081_ (
    .a(\DFF_1390.Q ),
    .b(\DFF_1253.Q ),
    .c(g35),
    .y(_01304_)
  );
  al_ao21ftf _06082_ (
    .a(g35),
    .b(\DFF_593.Q ),
    .c(_01304_),
    .y(\DFF_1253.D )
  );
  al_oai21ftf _06083_ (
    .a(\DFF_1269.Q ),
    .b(\DFF_48.Q ),
    .c(\DFF_760.Q ),
    .y(_01305_)
  );
  al_mux2h _06084_ (
    .a(\DFF_756.Q ),
    .b(_01305_),
    .s(g35),
    .y(\DFF_1269.D )
  );
  al_nand3ftt _06085_ (
    .a(\DFF_199.Q ),
    .b(\DFF_1408.Q ),
    .c(\DFF_245.Q ),
    .y(_01306_)
  );
  al_aoi21ftf _06086_ (
    .a(\DFF_19.Q ),
    .b(_01306_),
    .c(g35),
    .y(_01307_)
  );
  al_ao21ftf _06087_ (
    .a(_01306_),
    .b(_00499_),
    .c(_01307_),
    .y(_01308_)
  );
  al_ao21ftf _06088_ (
    .a(g35),
    .b(\DFF_626.Q ),
    .c(_01308_),
    .y(\DFF_19.D )
  );
  al_nor3ftt _06089_ (
    .a(\DFF_839.Q ),
    .b(_00499_),
    .c(_00365_),
    .y(_01309_)
  );
  al_oa21ftt _06090_ (
    .a(\DFF_839.Q ),
    .b(_00365_),
    .c(_00499_),
    .y(_01310_)
  );
  al_nor3ftt _06091_ (
    .a(g35),
    .b(_01309_),
    .c(_01310_),
    .y(\DFF_839.D )
  );
  al_or3 _06092_ (
    .a(\DFF_1304.Q ),
    .b(\DFF_1098.Q ),
    .c(\DFF_407.Q ),
    .y(_01311_)
  );
  al_and2ft _06093_ (
    .a(\DFF_598.Q ),
    .b(\DFF_68.Q ),
    .y(_01312_)
  );
  al_nand3ftt _06094_ (
    .a(_01311_),
    .b(_00499_),
    .c(_01312_),
    .y(_01313_)
  );
  al_ao21ftt _06095_ (
    .a(_01311_),
    .b(_01312_),
    .c(\DFF_1325.Q ),
    .y(_01314_)
  );
  al_nand3 _06096_ (
    .a(g35),
    .b(_01313_),
    .c(_01314_),
    .y(_01315_)
  );
  al_ao21ftf _06097_ (
    .a(g35),
    .b(\DFF_100.Q ),
    .c(_01315_),
    .y(\DFF_1325.D )
  );
  al_nand2 _06098_ (
    .a(\DFF_954.Q ),
    .b(\DFF_1275.Q ),
    .y(_01316_)
  );
  al_and3 _06099_ (
    .a(\DFF_954.Q ),
    .b(\DFF_431.Q ),
    .c(_00534_),
    .y(_01317_)
  );
  al_aoi21 _06100_ (
    .a(_01316_),
    .b(_00536_),
    .c(_01317_),
    .y(_01318_)
  );
  al_mux2h _06101_ (
    .a(\DFF_431.Q ),
    .b(_01318_),
    .s(g35),
    .y(\DFF_954.D )
  );
  al_and2 _06102_ (
    .a(g35),
    .b(_00745_),
    .y(_01319_)
  );
  al_ao21 _06103_ (
    .a(\DFF_635.Q ),
    .b(\DFF_270.Q ),
    .c(\DFF_1373.Q ),
    .y(_01320_)
  );
  al_nand3ftt _06104_ (
    .a(_00459_),
    .b(_01320_),
    .c(_01319_),
    .y(_01321_)
  );
  al_ao21ftf _06105_ (
    .a(g35),
    .b(\DFF_270.Q ),
    .c(_01321_),
    .y(\DFF_1373.D )
  );
  al_nand3 _06106_ (
    .a(\DFF_412.Q ),
    .b(\DFF_452.Q ),
    .c(_00460_),
    .y(_01322_)
  );
  al_and3 _06107_ (
    .a(\DFF_604.Q ),
    .b(\DFF_452.Q ),
    .c(_00459_),
    .y(_01323_)
  );
  al_and2 _06108_ (
    .a(\DFF_62.Q ),
    .b(_01323_),
    .y(_01324_)
  );
  al_and3ftt _06109_ (
    .a(_01324_),
    .b(g35),
    .c(_00745_),
    .y(_01325_)
  );
  al_ao21ftf _06110_ (
    .a(\DFF_62.Q ),
    .b(_01322_),
    .c(_01325_),
    .y(_01326_)
  );
  al_ao21ftf _06111_ (
    .a(g35),
    .b(\DFF_412.Q ),
    .c(_01326_),
    .y(\DFF_62.D )
  );
  al_inv _06112_ (
    .a(\DFF_449.Q ),
    .y(_01327_)
  );
  al_mux2l _06113_ (
    .a(\DFF_1285.Q ),
    .b(\DFF_1400.Q ),
    .s(\DFF_846.Q ),
    .y(_01328_)
  );
  al_aoi21 _06114_ (
    .a(\DFF_449.Q ),
    .b(_01328_),
    .c(\DFF_747.Q ),
    .y(_01329_)
  );
  al_ao21ftf _06115_ (
    .a(_01328_),
    .b(_01327_),
    .c(_01329_),
    .y(_01330_)
  );
  al_ao21ttf _06116_ (
    .a(_00462_),
    .b(_01330_),
    .c(g28753),
    .y(_01331_)
  );
  al_ao21 _06117_ (
    .a(\DFF_792.Q ),
    .b(_00009_),
    .c(\DFF_747.Q ),
    .y(_01332_)
  );
  al_and3 _06118_ (
    .a(g35),
    .b(_01332_),
    .c(_01331_),
    .y(\DFF_747.D )
  );
  al_mux2l _06119_ (
    .a(\DFF_518.Q ),
    .b(\DFF_639.Q ),
    .s(g84),
    .y(_01333_)
  );
  al_and2ft _06120_ (
    .a(\DFF_1238.Q ),
    .b(\DFF_539.Q ),
    .y(_01334_)
  );
  al_nand3 _06121_ (
    .a(\DFF_823.Q ),
    .b(_01333_),
    .c(_01334_),
    .y(_01335_)
  );
  al_and2 _06122_ (
    .a(\DFF_1238.Q ),
    .b(\DFF_1392.Q ),
    .y(_01336_)
  );
  al_nand3fft _06123_ (
    .a(\DFF_823.Q ),
    .b(_01333_),
    .c(_01336_),
    .y(_01337_)
  );
  al_and3 _06124_ (
    .a(\DFF_191.Q ),
    .b(\DFF_539.Q ),
    .c(\DFF_557.Q ),
    .y(_01338_)
  );
  al_and3fft _06125_ (
    .a(\DFF_191.Q ),
    .b(\DFF_557.Q ),
    .c(\DFF_1392.Q ),
    .y(_01339_)
  );
  al_nor3ftt _06126_ (
    .a(\DFF_1132.Q ),
    .b(_01339_),
    .c(_01338_),
    .y(_01340_)
  );
  al_nand3 _06127_ (
    .a(_01335_),
    .b(_01337_),
    .c(_01340_),
    .y(_01341_)
  );
  al_oai21ttf _06128_ (
    .a(_01339_),
    .b(_01338_),
    .c(\DFF_1132.Q ),
    .y(_01342_)
  );
  al_nand3 _06129_ (
    .a(g35),
    .b(_01342_),
    .c(_01341_),
    .y(_01343_)
  );
  al_aoi21ftf _06130_ (
    .a(\DFF_557.Q ),
    .b(_00066_),
    .c(_01343_),
    .y(\DFF_1132.D )
  );
  al_and2ft _06131_ (
    .a(\DFF_653.Q ),
    .b(\DFF_925.Q ),
    .y(_01344_)
  );
  al_nand3 _06132_ (
    .a(_00499_),
    .b(_01170_),
    .c(_01344_),
    .y(_01345_)
  );
  al_ao21 _06133_ (
    .a(_01170_),
    .b(_01344_),
    .c(\DFF_634.Q ),
    .y(_01346_)
  );
  al_nand3 _06134_ (
    .a(g35),
    .b(_01346_),
    .c(_01345_),
    .y(_01347_)
  );
  al_ao21ftf _06135_ (
    .a(g35),
    .b(\DFF_945.Q ),
    .c(_01347_),
    .y(\DFF_634.D )
  );
  al_and3ftt _06136_ (
    .a(\DFF_1232.Q ),
    .b(\DFF_1393.Q ),
    .c(\DFF_798.Q ),
    .y(_01348_)
  );
  al_or2ft _06137_ (
    .a(g35),
    .b(_01348_),
    .y(_01349_)
  );
  al_nand2ft _06138_ (
    .a(\DFF_900.Q ),
    .b(\DFF_866.Q ),
    .y(_01350_)
  );
  al_ao21 _06139_ (
    .a(_01350_),
    .b(_01348_),
    .c(_00066_),
    .y(_01351_)
  );
  al_ao21ftt _06140_ (
    .a(_01348_),
    .b(\DFF_447.Q ),
    .c(_01351_),
    .y(_01352_)
  );
  al_aoi21ftf _06141_ (
    .a(\DFF_622.Q ),
    .b(_01349_),
    .c(_01352_),
    .y(\DFF_447.D )
  );
  al_or2ft _06142_ (
    .a(g35),
    .b(_00369_),
    .y(_01353_)
  );
  al_mux2l _06143_ (
    .a(\DFF_918.Q ),
    .b(\DFF_651.Q ),
    .s(_01353_),
    .y(\DFF_651.D )
  );
  al_and2ft _06144_ (
    .a(\DFF_916.Q ),
    .b(\DFF_20.Q ),
    .y(_01354_)
  );
  al_nand3 _06145_ (
    .a(_00499_),
    .b(_01344_),
    .c(_01354_),
    .y(_01355_)
  );
  al_ao21 _06146_ (
    .a(_01344_),
    .b(_01354_),
    .c(\DFF_179.Q ),
    .y(_01356_)
  );
  al_nand3 _06147_ (
    .a(g35),
    .b(_01356_),
    .c(_01355_),
    .y(_01357_)
  );
  al_ao21ftf _06148_ (
    .a(g35),
    .b(\DFF_494.Q ),
    .c(_01357_),
    .y(\DFF_179.D )
  );
  al_inv _06149_ (
    .a(\DFF_54.Q ),
    .y(_01358_)
  );
  al_nand3 _06150_ (
    .a(_00364_),
    .b(_00556_),
    .c(_00363_),
    .y(_01359_)
  );
  al_and2ft _06151_ (
    .a(\DFF_35.Q ),
    .b(g35),
    .y(_01360_)
  );
  al_and3 _06152_ (
    .a(_01358_),
    .b(_01360_),
    .c(_01359_),
    .y(\DFF_35.D )
  );
  al_inv _06153_ (
    .a(\DFF_1070.Q ),
    .y(_01361_)
  );
  al_inv _06154_ (
    .a(\DFF_1295.Q ),
    .y(_01362_)
  );
  al_aoi21ftf _06155_ (
    .a(_00543_),
    .b(\DFF_931.Q ),
    .c(_00757_),
    .y(_01363_)
  );
  al_nand3fft _06156_ (
    .a(_01361_),
    .b(_01362_),
    .c(_01363_),
    .y(_01364_)
  );
  al_aoi21 _06157_ (
    .a(\DFF_888.Q ),
    .b(_01364_),
    .c(_00066_),
    .y(_01365_)
  );
  al_oai21 _06158_ (
    .a(\DFF_888.Q ),
    .b(_01364_),
    .c(_01365_),
    .y(_01366_)
  );
  al_aoi21ftf _06159_ (
    .a(\DFF_964.Q ),
    .b(_00066_),
    .c(_01366_),
    .y(\DFF_888.D )
  );
  al_or2 _06160_ (
    .a(\DFF_305.Q ),
    .b(\DFF_401.Q ),
    .y(_01367_)
  );
  al_ao21ttf _06161_ (
    .a(\DFF_1001.Q ),
    .b(\DFF_401.Q ),
    .c(_01367_),
    .y(_01368_)
  );
  al_and3fft _06162_ (
    .a(\DFF_181.Q ),
    .b(\DFF_642.Q ),
    .c(g35),
    .y(_01369_)
  );
  al_and3ftt _06163_ (
    .a(\DFF_785.Q ),
    .b(_01369_),
    .c(_01368_),
    .y(\DFF_1001.D )
  );
  al_oai21ftt _06164_ (
    .a(g35),
    .b(_01363_),
    .c(\DFF_1310.Q ),
    .y(_01370_)
  );
  al_and2ft _06165_ (
    .a(\DFF_1070.Q ),
    .b(\DFF_1236.Q ),
    .y(_01371_)
  );
  al_nand2 _06166_ (
    .a(_01371_),
    .b(_01363_),
    .y(_01372_)
  );
  al_nand3 _06167_ (
    .a(\DFF_1129.Q ),
    .b(g35),
    .c(_01372_),
    .y(_01373_)
  );
  al_and2ft _06168_ (
    .a(_01370_),
    .b(_01373_),
    .y(_01374_)
  );
  al_or2ft _06169_ (
    .a(_01370_),
    .b(_01373_),
    .y(_01375_)
  );
  al_nand2ft _06170_ (
    .a(_01374_),
    .b(_01375_),
    .y(\DFF_1129.D )
  );
  al_nor2 _06171_ (
    .a(\DFF_209.Q ),
    .b(g35),
    .y(_01376_)
  );
  al_and2 _06172_ (
    .a(\DFF_622.Q ),
    .b(_00319_),
    .y(_01377_)
  );
  al_and3ftt _06173_ (
    .a(_00525_),
    .b(_00604_),
    .c(_01377_),
    .y(_01378_)
  );
  al_oai21ftf _06174_ (
    .a(\DFF_1233.Q ),
    .b(\DFF_1010.Q ),
    .c(\DFF_1181.Q ),
    .y(_01379_)
  );
  al_nand3ftt _06175_ (
    .a(\DFF_1010.Q ),
    .b(\DFF_1233.Q ),
    .c(\DFF_1181.Q ),
    .y(_01380_)
  );
  al_nand3 _06176_ (
    .a(_01379_),
    .b(_01380_),
    .c(_01378_),
    .y(_01381_)
  );
  al_oa21ftf _06177_ (
    .a(\DFF_943.Q ),
    .b(_01378_),
    .c(_00066_),
    .y(_01382_)
  );
  al_aoi21 _06178_ (
    .a(_01381_),
    .b(_01382_),
    .c(_01376_),
    .y(\DFF_943.D )
  );
  al_aoi21 _06179_ (
    .a(\DFF_1062.Q ),
    .b(g35),
    .c(\DFF_969.Q ),
    .y(_01383_)
  );
  al_oa21ftt _06180_ (
    .a(g35),
    .b(\DFF_969.Q ),
    .c(\DFF_1062.Q ),
    .y(_01384_)
  );
  al_aoi21 _06181_ (
    .a(g35),
    .b(_01384_),
    .c(_01383_),
    .y(\DFF_1062.D )
  );
  al_mux2l _06182_ (
    .a(\DFF_133.Q ),
    .b(\DFF_208.Q ),
    .s(\DFF_675.Q ),
    .y(_01385_)
  );
  al_mux2h _06183_ (
    .a(\DFF_416.Q ),
    .b(_01385_),
    .s(g35),
    .y(\DFF_208.D )
  );
  al_nand2ft _06184_ (
    .a(\DFF_101.Q ),
    .b(\DFF_1352.Q ),
    .y(_01386_)
  );
  al_oai21ttf _06185_ (
    .a(\DFF_1335.Q ),
    .b(\DFF_117.Q ),
    .c(_00728_),
    .y(_01387_)
  );
  al_or2 _06186_ (
    .a(\DFF_263.Q ),
    .b(\DFF_101.Q ),
    .y(_01388_)
  );
  al_ao21ttf _06187_ (
    .a(\DFF_263.Q ),
    .b(\DFF_117.Q ),
    .c(_01388_),
    .y(_01389_)
  );
  al_and3 _06188_ (
    .a(_01386_),
    .b(_01389_),
    .c(_01387_),
    .y(_01390_)
  );
  al_and3ftt _06189_ (
    .a(_00729_),
    .b(g35),
    .c(_01390_),
    .y(\DFF_46.D )
  );
  al_oai21ftf _06190_ (
    .a(\DFF_317.Q ),
    .b(\DFF_166.Q ),
    .c(\DFF_259.Q ),
    .y(_01391_)
  );
  al_nand3ftt _06191_ (
    .a(\DFF_1256.Q ),
    .b(g35),
    .c(_01391_),
    .y(_01392_)
  );
  al_ao21ftf _06192_ (
    .a(g35),
    .b(\DFF_166.Q ),
    .c(_01392_),
    .y(\DFF_259.D )
  );
  al_or2ft _06193_ (
    .a(g35),
    .b(_00358_),
    .y(_01393_)
  );
  al_mux2l _06194_ (
    .a(\DFF_1138.Q ),
    .b(\DFF_14.Q ),
    .s(_01393_),
    .y(\DFF_14.D )
  );
  al_aoi21ftf _06195_ (
    .a(_00543_),
    .b(\DFF_284.Q ),
    .c(_00545_),
    .y(_01394_)
  );
  al_oai21ftt _06196_ (
    .a(g35),
    .b(_01394_),
    .c(\DFF_406.Q ),
    .y(_01395_)
  );
  al_and2ft _06197_ (
    .a(\DFF_387.Q ),
    .b(\DFF_297.Q ),
    .y(_01396_)
  );
  al_nand2 _06198_ (
    .a(_01396_),
    .b(_01394_),
    .y(_01397_)
  );
  al_nand3 _06199_ (
    .a(\DFF_804.Q ),
    .b(g35),
    .c(_01397_),
    .y(_01398_)
  );
  al_and2ft _06200_ (
    .a(_01395_),
    .b(_01398_),
    .y(_01399_)
  );
  al_or2ft _06201_ (
    .a(_01395_),
    .b(_01398_),
    .y(_01400_)
  );
  al_nand2ft _06202_ (
    .a(_01399_),
    .b(_01400_),
    .y(\DFF_804.D )
  );
  al_ao21ttf _06203_ (
    .a(_00983_),
    .b(_00585_),
    .c(\DFF_441.Q ),
    .y(_01401_)
  );
  al_nand2ft _06204_ (
    .a(\DFF_1360.Q ),
    .b(g35),
    .y(_01402_)
  );
  al_ao21 _06205_ (
    .a(_00983_),
    .b(_00585_),
    .c(_00066_),
    .y(_01403_)
  );
  al_ao21ftf _06206_ (
    .a(_01402_),
    .b(\DFF_693.Q ),
    .c(_01403_),
    .y(_01404_)
  );
  al_and3ftt _06207_ (
    .a(\DFF_693.Q ),
    .b(_01402_),
    .c(_01403_),
    .y(_01405_)
  );
  al_aoi21 _06208_ (
    .a(_01401_),
    .b(_01404_),
    .c(_01405_),
    .y(\DFF_441.D )
  );
  al_inv _06209_ (
    .a(\DFF_186.Q ),
    .y(_01406_)
  );
  al_nand3 _06210_ (
    .a(_01406_),
    .b(_00999_),
    .c(_00606_),
    .y(_01407_)
  );
  al_aoi21ttf _06211_ (
    .a(g35),
    .b(_01407_),
    .c(\DFF_674.Q ),
    .y(\DFF_186.D )
  );
  al_and2 _06212_ (
    .a(\DFF_598.Q ),
    .b(\DFF_68.Q ),
    .y(_01408_)
  );
  al_and2ft _06213_ (
    .a(\DFF_407.Q ),
    .b(\DFF_1304.Q ),
    .y(_01409_)
  );
  al_nand3 _06214_ (
    .a(_00499_),
    .b(_01408_),
    .c(_01409_),
    .y(_01410_)
  );
  al_ao21 _06215_ (
    .a(_01409_),
    .b(_01408_),
    .c(\DFF_1095.Q ),
    .y(_01411_)
  );
  al_nand3 _06216_ (
    .a(g35),
    .b(_01411_),
    .c(_01410_),
    .y(_01412_)
  );
  al_ao21ftf _06217_ (
    .a(g35),
    .b(\DFF_983.Q ),
    .c(_01412_),
    .y(\DFF_1095.D )
  );
  al_inv _06218_ (
    .a(\DFF_769.Q ),
    .y(_01413_)
  );
  al_inv _06219_ (
    .a(\DFF_1047.Q ),
    .y(_01414_)
  );
  al_nand3fft _06220_ (
    .a(_01413_),
    .b(_01414_),
    .c(_01282_),
    .y(_01415_)
  );
  al_aoi21ftf _06221_ (
    .a(\DFF_1026.Q ),
    .b(_01415_),
    .c(g35),
    .y(_01416_)
  );
  al_oai21 _06222_ (
    .a(_01284_),
    .b(_01415_),
    .c(_01416_),
    .y(_01417_)
  );
  al_ao21ftf _06223_ (
    .a(g35),
    .b(\DFF_204.Q ),
    .c(_01417_),
    .y(\DFF_1026.D )
  );
  al_and2ft _06224_ (
    .a(\DFF_1116.Q ),
    .b(\DFF_288.Q ),
    .y(_01418_)
  );
  al_and2ft _06225_ (
    .a(\DFF_883.Q ),
    .b(g35),
    .y(_01419_)
  );
  al_ao21ftf _06226_ (
    .a(\DFF_1124.Q ),
    .b(\DFF_288.Q ),
    .c(_01419_),
    .y(_01420_)
  );
  al_mux2l _06227_ (
    .a(_01419_),
    .b(_01420_),
    .s(\DFF_722.Q ),
    .y(_01421_)
  );
  al_ao21ftf _06228_ (
    .a(_00066_),
    .b(_01418_),
    .c(_01421_),
    .y(\DFF_883.D )
  );
  al_oa21ftt _06229_ (
    .a(g35),
    .b(\DFF_250.Q ),
    .c(\DFF_929.Q ),
    .y(_01422_)
  );
  al_or3 _06230_ (
    .a(\DFF_687.Q ),
    .b(\DFF_929.Q ),
    .c(\DFF_373.Q ),
    .y(_01423_)
  );
  al_or3 _06231_ (
    .a(\DFF_348.Q ),
    .b(\DFF_1225.Q ),
    .c(_01423_),
    .y(_01424_)
  );
  al_nor2 _06232_ (
    .a(_00503_),
    .b(_01424_),
    .y(_01425_)
  );
  al_ao21 _06233_ (
    .a(g35),
    .b(_01425_),
    .c(_01422_),
    .y(\DFF_348.D )
  );
  al_and3 _06234_ (
    .a(\DFF_1173.Q ),
    .b(\DFF_853.Q ),
    .c(_00601_),
    .y(_01426_)
  );
  al_oa21ftf _06235_ (
    .a(_00387_),
    .b(_01426_),
    .c(_00602_),
    .y(_01427_)
  );
  al_nand3 _06236_ (
    .a(g35),
    .b(_00606_),
    .c(_01427_),
    .y(_01428_)
  );
  al_ao21ftf _06237_ (
    .a(g35),
    .b(\DFF_1173.Q ),
    .c(_01428_),
    .y(\DFF_1374.D )
  );
  al_mux2l _06238_ (
    .a(\DFF_1016.Q ),
    .b(\DFF_440.Q ),
    .s(g35),
    .y(\DFF_436.D )
  );
  al_or2ft _06239_ (
    .a(g35),
    .b(_00373_),
    .y(_01429_)
  );
  al_mux2l _06240_ (
    .a(\DFF_644.Q ),
    .b(\DFF_1055.Q ),
    .s(_01429_),
    .y(\DFF_1055.D )
  );
  al_oai21ftt _06241_ (
    .a(\DFF_48.Q ),
    .b(\DFF_1269.Q ),
    .c(\DFF_756.Q ),
    .y(_01430_)
  );
  al_oa21 _06242_ (
    .a(\DFF_48.Q ),
    .b(\DFF_1269.Q ),
    .c(\DFF_760.Q ),
    .y(_01431_)
  );
  al_or3fft _06243_ (
    .a(g35),
    .b(_01430_),
    .c(_01431_),
    .y(_01432_)
  );
  al_aoi21ftf _06244_ (
    .a(\DFF_48.Q ),
    .b(_00066_),
    .c(_01432_),
    .y(\DFF_756.D )
  );
  al_mux2l _06245_ (
    .a(g6750),
    .b(\DFF_808.Q ),
    .s(g35),
    .y(\DFF_491.D )
  );
  al_and2 _06246_ (
    .a(\DFF_948.Q ),
    .b(g35),
    .y(\DFF_948.D )
  );
  al_oa21ftt _06247_ (
    .a(\DFF_605.Q ),
    .b(\DFF_787.Q ),
    .c(g35),
    .y(_01433_)
  );
  al_nand3fft _06248_ (
    .a(\DFF_1367.Q ),
    .b(\DFF_605.Q ),
    .c(g35),
    .y(_01434_)
  );
  al_aoi21ttf _06249_ (
    .a(_01434_),
    .b(_01433_),
    .c(\DFF_668.Q ),
    .y(\DFF_285.D )
  );
  al_inv _06250_ (
    .a(\DFF_928.Q ),
    .y(_01435_)
  );
  al_and2 _06251_ (
    .a(\DFF_387.Q ),
    .b(\DFF_681.Q ),
    .y(_01436_)
  );
  al_nand2 _06252_ (
    .a(_01436_),
    .b(_01394_),
    .y(_01437_)
  );
  al_aoi21 _06253_ (
    .a(\DFF_571.Q ),
    .b(_01437_),
    .c(_00066_),
    .y(_01438_)
  );
  al_oai21 _06254_ (
    .a(\DFF_571.Q ),
    .b(_01437_),
    .c(_01438_),
    .y(_01439_)
  );
  al_aoi21ftf _06255_ (
    .a(g35),
    .b(_01435_),
    .c(_01439_),
    .y(\DFF_571.D )
  );
  al_aoi21 _06256_ (
    .a(\DFF_385.Q ),
    .b(g35),
    .c(\DFF_393.Q ),
    .y(_01440_)
  );
  al_inv _06257_ (
    .a(\DFF_393.Q ),
    .y(_01441_)
  );
  al_nand3 _06258_ (
    .a(_00355_),
    .b(_00556_),
    .c(_00357_),
    .y(_01442_)
  );
  al_ao21ftf _06259_ (
    .a(_01441_),
    .b(\DFF_385.Q ),
    .c(_01442_),
    .y(_01443_)
  );
  al_aoi21 _06260_ (
    .a(g35),
    .b(_01443_),
    .c(_01440_),
    .y(\DFF_385.D )
  );
  al_nor2 _06261_ (
    .a(\DFF_1388.Q ),
    .b(g35),
    .y(_01444_)
  );
  al_inv _06262_ (
    .a(\DFF_140.Q ),
    .y(_01445_)
  );
  al_inv _06263_ (
    .a(\DFF_586.Q ),
    .y(_01446_)
  );
  al_and3fft _06264_ (
    .a(\DFF_762.Q ),
    .b(\DFF_36.Q ),
    .c(\DFF_805.Q ),
    .y(_01447_)
  );
  al_nand3fft _06265_ (
    .a(\DFF_1170.Q ),
    .b(\DFF_217.Q ),
    .c(_01447_),
    .y(_01448_)
  );
  al_or3fft _06266_ (
    .a(_01445_),
    .b(_01446_),
    .c(_01448_),
    .y(_01449_)
  );
  al_and3 _06267_ (
    .a(\DFF_762.Q ),
    .b(\DFF_36.Q ),
    .c(\DFF_1298.Q ),
    .y(_01450_)
  );
  al_and3 _06268_ (
    .a(\DFF_1170.Q ),
    .b(\DFF_217.Q ),
    .c(_01450_),
    .y(_01451_)
  );
  al_nand3fft _06269_ (
    .a(_01445_),
    .b(_01446_),
    .c(_01451_),
    .y(_01452_)
  );
  al_nand2 _06270_ (
    .a(\DFF_1388.Q ),
    .b(_01452_),
    .y(_01453_)
  );
  al_aoi21ftf _06271_ (
    .a(\DFF_1388.Q ),
    .b(_01449_),
    .c(_01453_),
    .y(_01454_)
  );
  al_aoi21ftf _06272_ (
    .a(_00710_),
    .b(_00711_),
    .c(_01119_),
    .y(_01455_)
  );
  al_or3fft _06273_ (
    .a(\DFF_703.Q ),
    .b(_01455_),
    .c(_01454_),
    .y(_01456_)
  );
  al_aoi21ftf _06274_ (
    .a(\DFF_703.Q ),
    .b(_01454_),
    .c(g35),
    .y(_01457_)
  );
  al_aoi21 _06275_ (
    .a(_01456_),
    .b(_01457_),
    .c(_01444_),
    .y(\DFF_703.D )
  );
  al_or2ft _06276_ (
    .a(g35),
    .b(g26801),
    .y(_01458_)
  );
  al_mux2l _06277_ (
    .a(\DFF_826.Q ),
    .b(\DFF_926.Q ),
    .s(_01458_),
    .y(\DFF_926.D )
  );
  al_and2ft _06278_ (
    .a(g35),
    .b(\DFF_149.Q ),
    .y(_01459_)
  );
  al_inv _06279_ (
    .a(\DFF_339.Q ),
    .y(_01460_)
  );
  al_and3 _06280_ (
    .a(\DFF_339.Q ),
    .b(\DFF_880.Q ),
    .c(\DFF_94.Q ),
    .y(_01461_)
  );
  al_and3 _06281_ (
    .a(\DFF_963.Q ),
    .b(\DFF_1241.Q ),
    .c(_01461_),
    .y(_01462_)
  );
  al_and3 _06282_ (
    .a(\DFF_303.Q ),
    .b(\DFF_280.Q ),
    .c(_01462_),
    .y(_01463_)
  );
  al_nand3 _06283_ (
    .a(\DFF_149.Q ),
    .b(\DFF_859.Q ),
    .c(_01463_),
    .y(_01464_)
  );
  al_ao21ftf _06284_ (
    .a(_01460_),
    .b(\DFF_867.Q ),
    .c(_01464_),
    .y(_01465_)
  );
  al_oa21ftf _06285_ (
    .a(\DFF_867.Q ),
    .b(_01464_),
    .c(_00066_),
    .y(_01466_)
  );
  al_ao21 _06286_ (
    .a(_01465_),
    .b(_01466_),
    .c(_01459_),
    .y(\DFF_867.D )
  );
  al_and2 _06287_ (
    .a(\DFF_734.Q ),
    .b(\DFF_723.Q ),
    .y(_01467_)
  );
  al_nand3 _06288_ (
    .a(_01441_),
    .b(_01467_),
    .c(_01442_),
    .y(_01468_)
  );
  al_ao21ftf _06289_ (
    .a(g35),
    .b(\DFF_723.Q ),
    .c(_01468_),
    .y(\DFF_393.D )
  );
  al_or2 _06290_ (
    .a(\DFF_421.Q ),
    .b(_00845_),
    .y(_01469_)
  );
  al_or3fft _06291_ (
    .a(g35),
    .b(_01469_),
    .c(_00846_),
    .y(_01470_)
  );
  al_ao21ftf _06292_ (
    .a(g35),
    .b(\DFF_788.Q ),
    .c(_01470_),
    .y(\DFF_421.D )
  );
  al_nand2 _06293_ (
    .a(\DFF_1275.Q ),
    .b(\DFF_1117.Q ),
    .y(_01471_)
  );
  al_nand2 _06294_ (
    .a(\DFF_1117.Q ),
    .b(_00533_),
    .y(_01472_)
  );
  al_aoi21ftf _06295_ (
    .a(_00533_),
    .b(_01471_),
    .c(_01472_),
    .y(_01473_)
  );
  al_mux2h _06296_ (
    .a(\DFF_1017.Q ),
    .b(_01473_),
    .s(g35),
    .y(\DFF_1117.D )
  );
  al_mux2l _06297_ (
    .a(\DFF_135.Q ),
    .b(\DFF_573.Q ),
    .s(_01054_),
    .y(\DFF_573.D )
  );
  al_or2 _06298_ (
    .a(\DFF_979.Q ),
    .b(\DFF_283.Q ),
    .y(_01474_)
  );
  al_nand3 _06299_ (
    .a(\DFF_788.Q ),
    .b(\DFF_131.Q ),
    .c(\DFF_70.Q ),
    .y(_01475_)
  );
  al_and3ftt _06300_ (
    .a(_01475_),
    .b(_00836_),
    .c(_00837_),
    .y(_01476_)
  );
  al_ao21 _06301_ (
    .a(_00844_),
    .b(_01476_),
    .c(_01474_),
    .y(_01477_)
  );
  al_nand3ftt _06302_ (
    .a(\DFF_208.Q ),
    .b(\DFF_133.Q ),
    .c(\DFF_606.Q ),
    .y(_01478_)
  );
  al_and3ftt _06303_ (
    .a(_01478_),
    .b(\DFF_675.Q ),
    .c(_01477_),
    .y(_01479_)
  );
  al_and2ft _06304_ (
    .a(\DFF_214.Q ),
    .b(\DFF_563.Q ),
    .y(_01480_)
  );
  al_and3 _06305_ (
    .a(\DFF_675.Q ),
    .b(_01478_),
    .c(_01480_),
    .y(_01481_)
  );
  al_nand3 _06306_ (
    .a(\DFF_936.Q ),
    .b(\DFF_277.Q ),
    .c(_01481_),
    .y(_01482_)
  );
  al_oai21ftf _06307_ (
    .a(\DFF_1237.Q ),
    .b(_01482_),
    .c(_00066_),
    .y(_01483_)
  );
  al_oai21ttf _06308_ (
    .a(\DFF_1237.Q ),
    .b(_01479_),
    .c(_01483_),
    .y(_01484_)
  );
  al_ao21ftf _06309_ (
    .a(g35),
    .b(\DFF_208.Q ),
    .c(_01484_),
    .y(\DFF_1237.D )
  );
  al_or3 _06310_ (
    .a(\DFF_439.Q ),
    .b(g73),
    .c(g72),
    .y(_01485_)
  );
  al_mux2l _06311_ (
    .a(_01485_),
    .b(\DFF_1330.Q ),
    .s(_01208_),
    .y(\DFF_1349.D )
  );
  al_inv _06312_ (
    .a(\DFF_1051.Q ),
    .y(_01486_)
  );
  al_nor2 _06313_ (
    .a(\DFF_583.Q ),
    .b(\DFF_1216.Q ),
    .y(_01487_)
  );
  al_and3ftt _06314_ (
    .a(\DFF_964.Q ),
    .b(_01486_),
    .c(_01487_),
    .y(_01488_)
  );
  al_nor2 _06315_ (
    .a(\DFF_301.Q ),
    .b(\DFF_818.Q ),
    .y(_01489_)
  );
  al_nand3fft _06316_ (
    .a(\DFF_45.Q ),
    .b(\DFF_928.Q ),
    .c(_01489_),
    .y(_01490_)
  );
  al_or3ftt _06317_ (
    .a(_01488_),
    .b(\DFF_364.Q ),
    .c(_01490_),
    .y(_01491_)
  );
  al_mux2h _06318_ (
    .a(\DFF_1301.Q ),
    .b(_01491_),
    .s(g35),
    .y(\DFF_364.D )
  );
  al_nor2 _06319_ (
    .a(\DFF_1341.Q ),
    .b(g35),
    .y(_01492_)
  );
  al_mux2l _06320_ (
    .a(\DFF_1065.Q ),
    .b(\DFF_366.Q ),
    .s(\DFF_1341.Q ),
    .y(_01493_)
  );
  al_nand3ftt _06321_ (
    .a(_01493_),
    .b(\DFF_432.Q ),
    .c(_01101_),
    .y(_01494_)
  );
  al_aoi21ftf _06322_ (
    .a(\DFF_432.Q ),
    .b(_01493_),
    .c(g35),
    .y(_01495_)
  );
  al_aoi21 _06323_ (
    .a(_01495_),
    .b(_01494_),
    .c(_01492_),
    .y(\DFF_432.D )
  );
  al_and2 _06324_ (
    .a(g35),
    .b(_00557_),
    .y(_01496_)
  );
  al_and3ftt _06325_ (
    .a(\DFF_407.Q ),
    .b(_00555_),
    .c(_01496_),
    .y(\DFF_407.D )
  );
  al_and2ft _06326_ (
    .a(\DFF_120.Q ),
    .b(\DFF_27.Q ),
    .y(_01497_)
  );
  al_nand3 _06327_ (
    .a(_00499_),
    .b(_01045_),
    .c(_01497_),
    .y(_01498_)
  );
  al_ao21 _06328_ (
    .a(_01045_),
    .b(_01497_),
    .c(\DFF_1052.Q ),
    .y(_01499_)
  );
  al_nand3 _06329_ (
    .a(g35),
    .b(_01499_),
    .c(_01498_),
    .y(_01500_)
  );
  al_ao21ftf _06330_ (
    .a(g35),
    .b(\DFF_321.Q ),
    .c(_01500_),
    .y(\DFF_1052.D )
  );
  al_and2 _06331_ (
    .a(\DFF_326.Q ),
    .b(\DFF_30.Q ),
    .y(_01501_)
  );
  al_and3 _06332_ (
    .a(\DFF_797.Q ),
    .b(\DFF_110.Q ),
    .c(_01501_),
    .y(_01502_)
  );
  al_and2 _06333_ (
    .a(\DFF_1320.Q ),
    .b(g35),
    .y(_01503_)
  );
  al_aoi21ttf _06334_ (
    .a(_01503_),
    .b(_01502_),
    .c(\DFF_543.Q ),
    .y(\DFF_731.D )
  );
  al_nand2 _06335_ (
    .a(\DFF_853.Q ),
    .b(_00601_),
    .y(_01504_)
  );
  al_and2 _06336_ (
    .a(g35),
    .b(_00606_),
    .y(_01505_)
  );
  al_nor2 _06337_ (
    .a(\DFF_853.Q ),
    .b(_00601_),
    .y(_01506_)
  );
  al_ao21ftf _06338_ (
    .a(_01506_),
    .b(_01504_),
    .c(_01505_),
    .y(_01507_)
  );
  al_aoi21ftf _06339_ (
    .a(\DFF_186.Q ),
    .b(_00066_),
    .c(_01507_),
    .y(\DFF_853.D )
  );
  al_mux2l _06340_ (
    .a(\DFF_1164.Q ),
    .b(\DFF_1045.Q ),
    .s(_00478_),
    .y(_01508_)
  );
  al_mux2h _06341_ (
    .a(\DFF_601.Q ),
    .b(_01508_),
    .s(g35),
    .y(\DFF_1045.D )
  );
  al_nand2ft _06342_ (
    .a(\DFF_1239.Q ),
    .b(\DFF_1405.Q ),
    .y(_01509_)
  );
  al_nand3 _06343_ (
    .a(\DFF_801.Q ),
    .b(g35),
    .c(_01509_),
    .y(_01510_)
  );
  al_nand2ft _06344_ (
    .a(\DFF_513.Q ),
    .b(\DFF_1405.Q ),
    .y(_01511_)
  );
  al_mux2l _06345_ (
    .a(\DFF_801.Q ),
    .b(\DFF_1405.Q ),
    .s(g35),
    .y(_01512_)
  );
  al_aoi21ftf _06346_ (
    .a(_01512_),
    .b(_01511_),
    .c(_01510_),
    .y(\DFF_578.D )
  );
  al_mux2l _06347_ (
    .a(\DFF_1407.Q ),
    .b(\DFF_202.Q ),
    .s(\DFF_60.Q ),
    .y(_01513_)
  );
  al_mux2h _06348_ (
    .a(\DFF_1131.Q ),
    .b(_01513_),
    .s(g35),
    .y(\DFF_202.D )
  );
  al_and3ftt _06349_ (
    .a(\DFF_1236.Q ),
    .b(\DFF_1070.Q ),
    .c(\DFF_641.Q ),
    .y(_01514_)
  );
  al_and3fft _06350_ (
    .a(\DFF_1070.Q ),
    .b(\DFF_1295.Q ),
    .c(\DFF_465.Q ),
    .y(_01515_)
  );
  al_and2ft _06351_ (
    .a(\DFF_1236.Q ),
    .b(\DFF_1295.Q ),
    .y(_01516_)
  );
  al_ao21 _06352_ (
    .a(\DFF_924.Q ),
    .b(_01516_),
    .c(_01515_),
    .y(_01517_)
  );
  al_inv _06353_ (
    .a(\DFF_1394.Q ),
    .y(_01518_)
  );
  al_and3 _06354_ (
    .a(\DFF_1070.Q ),
    .b(\DFF_1295.Q ),
    .c(\DFF_255.Q ),
    .y(_01519_)
  );
  al_aoi21 _06355_ (
    .a(\DFF_809.Q ),
    .b(_00439_),
    .c(_01519_),
    .y(_01520_)
  );
  al_aoi21ftf _06356_ (
    .a(_01518_),
    .b(_01371_),
    .c(_01520_),
    .y(_01521_)
  );
  al_nand3fft _06357_ (
    .a(_01514_),
    .b(_01517_),
    .c(_01521_),
    .y(_01522_)
  );
  al_mux2h _06358_ (
    .a(\DFF_1310.Q ),
    .b(_01522_),
    .s(_01363_),
    .y(_01523_)
  );
  al_mux2h _06359_ (
    .a(\DFF_1295.Q ),
    .b(_01523_),
    .s(g35),
    .y(\DFF_1310.D )
  );
  al_nand3ftt _06360_ (
    .a(\DFF_440.Q ),
    .b(g113),
    .c(\DFF_1016.Q ),
    .y(_01524_)
  );
  al_oai21ftt _06361_ (
    .a(\DFF_1016.Q ),
    .b(\DFF_440.Q ),
    .c(\DFF_1399.Q ),
    .y(_01525_)
  );
  al_nand3 _06362_ (
    .a(g35),
    .b(_01524_),
    .c(_01525_),
    .y(\DFF_1399.D )
  );
  al_and3 _06363_ (
    .a(\DFF_43.Q ),
    .b(\DFF_1412.Q ),
    .c(\DFF_331.Q ),
    .y(_01526_)
  );
  al_oa21ttf _06364_ (
    .a(\DFF_674.Q ),
    .b(_01526_),
    .c(_00066_),
    .y(_01527_)
  );
  al_aoi21ttf _06365_ (
    .a(\DFF_674.Q ),
    .b(_01526_),
    .c(_01527_),
    .y(_01528_)
  );
  al_nand3 _06366_ (
    .a(_01406_),
    .b(_00606_),
    .c(_01528_),
    .y(_01529_)
  );
  al_ao21ftf _06367_ (
    .a(g35),
    .b(\DFF_1412.Q ),
    .c(_01529_),
    .y(\DFF_674.D )
  );
  al_and2 _06368_ (
    .a(\DFF_759.Q ),
    .b(_01125_),
    .y(_01530_)
  );
  al_nand3 _06369_ (
    .a(\DFF_1181.Q ),
    .b(_00604_),
    .c(_00326_),
    .y(_01531_)
  );
  al_oai21ftf _06370_ (
    .a(\DFF_620.Q ),
    .b(_01125_),
    .c(_00066_),
    .y(_01532_)
  );
  al_ao21 _06371_ (
    .a(_01530_),
    .b(_01531_),
    .c(_01532_),
    .y(_01533_)
  );
  al_aoi21ftf _06372_ (
    .a(\DFF_759.Q ),
    .b(_00066_),
    .c(_01533_),
    .y(\DFF_620.D )
  );
  al_inv _06373_ (
    .a(\DFF_1143.Q ),
    .y(_01534_)
  );
  al_inv _06374_ (
    .a(\DFF_886.Q ),
    .y(_01535_)
  );
  al_nand3fft _06375_ (
    .a(_01534_),
    .b(_01535_),
    .c(_00974_),
    .y(_01536_)
  );
  al_aoi21ftf _06376_ (
    .a(\DFF_1171.Q ),
    .b(_01536_),
    .c(g35),
    .y(_01537_)
  );
  al_oai21 _06377_ (
    .a(_00977_),
    .b(_01536_),
    .c(_01537_),
    .y(_01538_)
  );
  al_ao21ftf _06378_ (
    .a(g35),
    .b(\DFF_1025.Q ),
    .c(_01538_),
    .y(\DFF_1171.D )
  );
  al_aoi21ttf _06379_ (
    .a(\DFF_606.Q ),
    .b(\DFF_675.Q ),
    .c(g35),
    .y(_01539_)
  );
  al_ao21ftf _06380_ (
    .a(\DFF_675.Q ),
    .b(\DFF_133.Q ),
    .c(_01539_),
    .y(_01540_)
  );
  al_aoi21ftf _06381_ (
    .a(\DFF_563.Q ),
    .b(_00066_),
    .c(_01540_),
    .y(\DFF_133.D )
  );
  al_nor2 _06382_ (
    .a(_00066_),
    .b(_00546_),
    .y(_01541_)
  );
  al_inv _06383_ (
    .a(\DFF_1037.Q ),
    .y(_01542_)
  );
  al_and3 _06384_ (
    .a(_00433_),
    .b(_00604_),
    .c(_00422_),
    .y(_01543_)
  );
  al_aoi21ttf _06385_ (
    .a(\DFF_379.Q ),
    .b(_01543_),
    .c(_00546_),
    .y(_01544_)
  );
  al_nand2 _06386_ (
    .a(_01542_),
    .b(_01544_),
    .y(_01545_)
  );
  al_mux2h _06387_ (
    .a(\DFF_153.Q ),
    .b(_01545_),
    .s(g35),
    .y(_01546_)
  );
  al_aoi21ftf _06388_ (
    .a(\DFF_1375.Q ),
    .b(_01541_),
    .c(_01546_),
    .y(\DFF_1375.D )
  );
  al_or3 _06389_ (
    .a(\DFF_1273.Q ),
    .b(\DFF_410.Q ),
    .c(\DFF_584.Q ),
    .y(_01547_)
  );
  al_nand3ftt _06390_ (
    .a(_01547_),
    .b(_00499_),
    .c(_01105_),
    .y(_01548_)
  );
  al_ao21ftt _06391_ (
    .a(_01547_),
    .b(_01105_),
    .c(\DFF_1032.Q ),
    .y(_01549_)
  );
  al_nand3 _06392_ (
    .a(g35),
    .b(_01548_),
    .c(_01549_),
    .y(_01550_)
  );
  al_ao21ftf _06393_ (
    .a(g35),
    .b(\DFF_967.Q ),
    .c(_01550_),
    .y(\DFF_1032.D )
  );
  al_nand3 _06394_ (
    .a(_00499_),
    .b(_00691_),
    .c(_01266_),
    .y(_01551_)
  );
  al_ao21 _06395_ (
    .a(_01266_),
    .b(_00691_),
    .c(\DFF_257.Q ),
    .y(_01552_)
  );
  al_nand3 _06396_ (
    .a(g35),
    .b(_01552_),
    .c(_01551_),
    .y(_01553_)
  );
  al_ao21ftf _06397_ (
    .a(g35),
    .b(\DFF_479.Q ),
    .c(_01553_),
    .y(\DFF_257.D )
  );
  al_and2 _06398_ (
    .a(\DFF_188.Q ),
    .b(\DFF_554.Q ),
    .y(_01554_)
  );
  al_and3 _06399_ (
    .a(\DFF_474.Q ),
    .b(\DFF_315.Q ),
    .c(_01554_),
    .y(_01555_)
  );
  al_and2 _06400_ (
    .a(\DFF_1005.Q ),
    .b(g35),
    .y(_01556_)
  );
  al_aoi21ttf _06401_ (
    .a(_01556_),
    .b(_01555_),
    .c(\DFF_251.Q ),
    .y(\DFF_1188.D )
  );
  al_nand3fft _06402_ (
    .a(\DFF_669.Q ),
    .b(\DFF_799.Q ),
    .c(\DFF_736.Q ),
    .y(_01557_)
  );
  al_mux2l _06403_ (
    .a(\DFF_382.Q ),
    .b(\DFF_585.Q ),
    .s(_01557_),
    .y(_01558_)
  );
  al_mux2h _06404_ (
    .a(\DFF_1003.Q ),
    .b(_01558_),
    .s(g35),
    .y(\DFF_382.D )
  );
  al_and3ftt _06405_ (
    .a(g113),
    .b(\DFF_1111.Q ),
    .c(_00342_),
    .y(_01559_)
  );
  al_oa21ftf _06406_ (
    .a(\DFF_811.Q ),
    .b(_00604_),
    .c(_01559_),
    .y(_01560_)
  );
  al_mux2l _06407_ (
    .a(\DFF_931.Q ),
    .b(_01560_),
    .s(_00697_),
    .y(_01561_)
  );
  al_mux2h _06408_ (
    .a(\DFF_811.Q ),
    .b(_01561_),
    .s(g35),
    .y(\DFF_931.D )
  );
  al_and2 _06409_ (
    .a(\DFF_812.Q ),
    .b(_01236_),
    .y(_01562_)
  );
  al_ao21 _06410_ (
    .a(\DFF_812.Q ),
    .b(_01183_),
    .c(_01236_),
    .y(_01563_)
  );
  al_or3fft _06411_ (
    .a(g35),
    .b(_01563_),
    .c(_01562_),
    .y(_01564_)
  );
  al_ao21ftf _06412_ (
    .a(g35),
    .b(\DFF_89.Q ),
    .c(_01564_),
    .y(\DFF_812.D )
  );
  al_mux2l _06413_ (
    .a(\DFF_489.Q ),
    .b(\DFF_770.Q ),
    .s(g35),
    .y(\DFF_489.D )
  );
  al_and2 _06414_ (
    .a(g35),
    .b(g125),
    .y(\DFF_126.D )
  );
  al_and3fft _06415_ (
    .a(\DFF_325.Q ),
    .b(\DFF_739.Q ),
    .c(g35),
    .y(_01565_)
  );
  al_ao21ftt _06416_ (
    .a(g35),
    .b(\DFF_1387.Q ),
    .c(_01565_),
    .y(\DFF_739.D )
  );
  al_nand3 _06417_ (
    .a(_00499_),
    .b(_01169_),
    .c(_01354_),
    .y(_01566_)
  );
  al_ao21 _06418_ (
    .a(_01169_),
    .b(_01354_),
    .c(\DFF_904.Q ),
    .y(_01567_)
  );
  al_nand3 _06419_ (
    .a(g35),
    .b(_01567_),
    .c(_01566_),
    .y(_01568_)
  );
  al_ao21ftf _06420_ (
    .a(g35),
    .b(\DFF_179.Q ),
    .c(_01568_),
    .y(\DFF_904.D )
  );
  al_mux2h _06421_ (
    .a(\DFF_250.Q ),
    .b(_00604_),
    .s(g35),
    .y(\DFF_1272.D )
  );
  al_nand2 _06422_ (
    .a(g35),
    .b(_00722_),
    .y(_01569_)
  );
  al_mux2l _06423_ (
    .a(\DFF_293.Q ),
    .b(\DFF_1266.Q ),
    .s(_01569_),
    .y(\DFF_1266.D )
  );
  al_nand3 _06424_ (
    .a(g35),
    .b(\DFF_1164.Q ),
    .c(_01050_),
    .y(_01570_)
  );
  al_ao21ftf _06425_ (
    .a(_01174_),
    .b(\DFF_237.Q ),
    .c(_01570_),
    .y(\DFF_237.D )
  );
  al_mux2l _06426_ (
    .a(g6748),
    .b(\DFF_38.Q ),
    .s(g35),
    .y(\DFF_121.D )
  );
  al_nand3ftt _06427_ (
    .a(\DFF_1068.Q ),
    .b(\DFF_1150.Q ),
    .c(\DFF_1273.Q ),
    .y(_01571_)
  );
  al_aoi21ftf _06428_ (
    .a(\DFF_1175.Q ),
    .b(_01571_),
    .c(g35),
    .y(_01572_)
  );
  al_ao21ftf _06429_ (
    .a(_01571_),
    .b(_00499_),
    .c(_01572_),
    .y(_01573_)
  );
  al_ao21ftf _06430_ (
    .a(g35),
    .b(\DFF_464.Q ),
    .c(_01573_),
    .y(\DFF_1175.D )
  );
  al_nand3fft _06431_ (
    .a(_01542_),
    .b(\DFF_1375.Q ),
    .c(_00546_),
    .y(_01574_)
  );
  al_and2ft _06432_ (
    .a(\DFF_272.Q ),
    .b(\DFF_500.Q ),
    .y(_01575_)
  );
  al_inv _06433_ (
    .a(\DFF_984.Q ),
    .y(_01576_)
  );
  al_aoi21 _06434_ (
    .a(_01576_),
    .b(_01574_),
    .c(_00066_),
    .y(_01577_)
  );
  al_ao21ftf _06435_ (
    .a(_01574_),
    .b(_01575_),
    .c(_01577_),
    .y(_01578_)
  );
  al_ao21ftf _06436_ (
    .a(g35),
    .b(\DFF_306.Q ),
    .c(_01578_),
    .y(\DFF_984.D )
  );
  al_and3 _06437_ (
    .a(\DFF_1161.Q ),
    .b(g35),
    .c(_00477_),
    .y(_01579_)
  );
  al_or2 _06438_ (
    .a(\DFF_1108.Q ),
    .b(g35),
    .y(_01580_)
  );
  al_aoi21ftf _06439_ (
    .a(\DFF_346.Q ),
    .b(_01579_),
    .c(_01580_),
    .y(_01581_)
  );
  al_oa21 _06440_ (
    .a(\DFF_510.Q ),
    .b(_01174_),
    .c(_01581_),
    .y(\DFF_510.D )
  );
  al_and3 _06441_ (
    .a(\DFF_1393.Q ),
    .b(\DFF_1232.Q ),
    .c(\DFF_269.Q ),
    .y(_01582_)
  );
  al_ao21ftt _06442_ (
    .a(g35),
    .b(\DFF_1393.Q ),
    .c(_01582_),
    .y(\DFF_96.D )
  );
  al_oa21ftt _06443_ (
    .a(g35),
    .b(\DFF_798.Q ),
    .c(\DFF_1232.Q ),
    .y(_01583_)
  );
  al_or3fft _06444_ (
    .a(\DFF_1393.Q ),
    .b(g35),
    .c(_01583_),
    .y(_01584_)
  );
  al_aoi21ttf _06445_ (
    .a(\DFF_1393.Q ),
    .b(g35),
    .c(_01583_),
    .y(_01585_)
  );
  al_nand2ft _06446_ (
    .a(_01585_),
    .b(_01584_),
    .y(\DFF_1393.D )
  );
  al_nor2 _06447_ (
    .a(\DFF_1054.Q ),
    .b(g35),
    .y(_01586_)
  );
  al_and3ftt _06448_ (
    .a(_00348_),
    .b(_00604_),
    .c(_00339_),
    .y(_01587_)
  );
  al_oai21ftf _06449_ (
    .a(\DFF_646.Q ),
    .b(\DFF_1127.Q ),
    .c(\DFF_1181.Q ),
    .y(_01588_)
  );
  al_nand3ftt _06450_ (
    .a(\DFF_1127.Q ),
    .b(\DFF_646.Q ),
    .c(\DFF_1181.Q ),
    .y(_01589_)
  );
  al_nand3 _06451_ (
    .a(_01588_),
    .b(_01589_),
    .c(_01587_),
    .y(_01590_)
  );
  al_oa21ftf _06452_ (
    .a(\DFF_1089.Q ),
    .b(_01587_),
    .c(_00066_),
    .y(_01591_)
  );
  al_aoi21 _06453_ (
    .a(_01590_),
    .b(_01591_),
    .c(_01586_),
    .y(\DFF_1089.D )
  );
  al_nand2 _06454_ (
    .a(g35),
    .b(_01195_),
    .y(_01592_)
  );
  al_mux2l _06455_ (
    .a(\DFF_888.Q ),
    .b(\DFF_1086.Q ),
    .s(_01592_),
    .y(\DFF_1086.D )
  );
  al_and2 _06456_ (
    .a(\DFF_303.Q ),
    .b(_01462_),
    .y(_01593_)
  );
  al_nand2 _06457_ (
    .a(\DFF_280.Q ),
    .b(\DFF_339.Q ),
    .y(_01594_)
  );
  al_oa21ftf _06458_ (
    .a(_01594_),
    .b(_01593_),
    .c(_01463_),
    .y(_01595_)
  );
  al_mux2h _06459_ (
    .a(\DFF_303.Q ),
    .b(_01595_),
    .s(g35),
    .y(\DFF_280.D )
  );
  al_and2ft _06460_ (
    .a(g35),
    .b(\DFF_112.Q ),
    .y(_01596_)
  );
  al_nor3fft _06461_ (
    .a(\DFF_902.Q ),
    .b(_01050_),
    .c(_00871_),
    .y(_01597_)
  );
  al_nand3 _06462_ (
    .a(\DFF_112.Q ),
    .b(\DFF_1019.Q ),
    .c(_01597_),
    .y(_01598_)
  );
  al_and3 _06463_ (
    .a(\DFF_112.Q ),
    .b(\DFF_902.Q ),
    .c(_00872_),
    .y(_01599_)
  );
  al_nor2 _06464_ (
    .a(\DFF_135.Q ),
    .b(\DFF_656.Q ),
    .y(_01600_)
  );
  al_and3fft _06465_ (
    .a(\DFF_1126.Q ),
    .b(\DFF_1042.Q ),
    .c(\DFF_1250.Q ),
    .y(_01601_)
  );
  al_and2 _06466_ (
    .a(\DFF_238.Q ),
    .b(_01601_),
    .y(_01602_)
  );
  al_nand2 _06467_ (
    .a(\DFF_1365.Q ),
    .b(\DFF_573.Q ),
    .y(_01603_)
  );
  al_aoi21ftf _06468_ (
    .a(_00873_),
    .b(_01603_),
    .c(_01602_),
    .y(_01604_)
  );
  al_aoi21ftf _06469_ (
    .a(_01600_),
    .b(_00483_),
    .c(_01604_),
    .y(_01605_)
  );
  al_nand2 _06470_ (
    .a(\DFF_667.Q ),
    .b(g35),
    .y(_01606_)
  );
  al_aoi21 _06471_ (
    .a(_00872_),
    .b(_01605_),
    .c(_01606_),
    .y(_01607_)
  );
  al_oa21 _06472_ (
    .a(\DFF_1019.Q ),
    .b(_01599_),
    .c(_01607_),
    .y(_01608_)
  );
  al_ao21 _06473_ (
    .a(_01598_),
    .b(_01608_),
    .c(_01596_),
    .y(\DFF_1019.D )
  );
  al_mux2h _06474_ (
    .a(\DFF_879.Q ),
    .b(_00894_),
    .s(g35),
    .y(\DFF_821.D )
  );
  al_mux2l _06475_ (
    .a(\DFF_974.Q ),
    .b(\DFF_1340.Q ),
    .s(g35),
    .y(\DFF_974.D )
  );
  al_and2ft _06476_ (
    .a(g35),
    .b(\DFF_1129.Q ),
    .y(_01609_)
  );
  al_nand2ft _06477_ (
    .a(\DFF_77.Q ),
    .b(\DFF_1129.Q ),
    .y(_01610_)
  );
  al_nand2ft _06478_ (
    .a(\DFF_1129.Q ),
    .b(\DFF_77.Q ),
    .y(_01611_)
  );
  al_or3fft _06479_ (
    .a(_01610_),
    .b(_01611_),
    .c(_01372_),
    .y(_01612_)
  );
  al_aoi21ftf _06480_ (
    .a(\DFF_964.Q ),
    .b(_01372_),
    .c(g35),
    .y(_01613_)
  );
  al_ao21 _06481_ (
    .a(_01612_),
    .b(_01613_),
    .c(_01609_),
    .y(\DFF_964.D )
  );
  al_inv _06482_ (
    .a(\DFF_713.Q ),
    .y(_01614_)
  );
  al_inv _06483_ (
    .a(\DFF_505.Q ),
    .y(_01615_)
  );
  al_nand3fft _06484_ (
    .a(_01614_),
    .b(_01615_),
    .c(_00641_),
    .y(_01616_)
  );
  al_aoi21ftf _06485_ (
    .a(_00638_),
    .b(_00528_),
    .c(_00637_),
    .y(_01617_)
  );
  al_aoi21ftf _06486_ (
    .a(\DFF_481.Q ),
    .b(_00638_),
    .c(_01617_),
    .y(_01618_)
  );
  al_aoi21ftf _06487_ (
    .a(\DFF_960.Q ),
    .b(_01616_),
    .c(g35),
    .y(_01619_)
  );
  al_ao21ftf _06488_ (
    .a(_01616_),
    .b(_01618_),
    .c(_01619_),
    .y(_01620_)
  );
  al_ao21ftf _06489_ (
    .a(g35),
    .b(\DFF_890.Q ),
    .c(_01620_),
    .y(\DFF_960.D )
  );
  al_and3 _06490_ (
    .a(\DFF_1420.Q ),
    .b(\DFF_468.Q ),
    .c(\DFF_220.Q ),
    .y(_01621_)
  );
  al_and2 _06491_ (
    .a(\DFF_942.Q ),
    .b(_01621_),
    .y(_01622_)
  );
  al_and2 _06492_ (
    .a(\DFF_664.Q ),
    .b(g35),
    .y(_01623_)
  );
  al_aoi21ttf _06493_ (
    .a(_01623_),
    .b(_01622_),
    .c(\DFF_1214.Q ),
    .y(\DFF_39.D )
  );
  al_aoi21 _06494_ (
    .a(\DFF_1320.Q ),
    .b(_01502_),
    .c(_00066_),
    .y(_01624_)
  );
  al_nand2ft _06495_ (
    .a(g35),
    .b(\DFF_1320.Q ),
    .y(_01625_)
  );
  al_ao21ftf _06496_ (
    .a(\DFF_731.Q ),
    .b(_01624_),
    .c(_01625_),
    .y(\DFF_543.D )
  );
  al_or2ft _06497_ (
    .a(g35),
    .b(_00365_),
    .y(_01626_)
  );
  al_mux2l _06498_ (
    .a(\DFF_839.Q ),
    .b(\DFF_124.Q ),
    .s(_01626_),
    .y(\DFF_124.D )
  );
  al_nor2 _06499_ (
    .a(\DFF_1309.Q ),
    .b(g35),
    .y(_01627_)
  );
  al_and3 _06500_ (
    .a(\DFF_475.Q ),
    .b(\DFF_516.Q ),
    .c(\DFF_478.Q ),
    .y(_01628_)
  );
  al_nand3 _06501_ (
    .a(\DFF_1309.Q ),
    .b(\DFF_741.Q ),
    .c(_01628_),
    .y(_01629_)
  );
  al_nand2 _06502_ (
    .a(\DFF_1077.Q ),
    .b(_01629_),
    .y(_01630_)
  );
  al_and3fft _06503_ (
    .a(\DFF_475.Q ),
    .b(\DFF_516.Q ),
    .c(\DFF_405.Q ),
    .y(_01631_)
  );
  al_and3fft _06504_ (
    .a(\DFF_1309.Q ),
    .b(\DFF_741.Q ),
    .c(_01631_),
    .y(_01632_)
  );
  al_inv _06505_ (
    .a(\DFF_1334.Q ),
    .y(_01633_)
  );
  al_nand2 _06506_ (
    .a(\DFF_335.Q ),
    .b(\DFF_381.Q ),
    .y(_01634_)
  );
  al_nand2 _06507_ (
    .a(\DFF_1077.Q ),
    .b(\DFF_335.Q ),
    .y(_01635_)
  );
  al_mux2l _06508_ (
    .a(_01634_),
    .b(_01635_),
    .s(_00890_),
    .y(_01636_)
  );
  al_or3fft _06509_ (
    .a(_01633_),
    .b(\DFF_478.Q ),
    .c(_01636_),
    .y(_01637_)
  );
  al_nor2 _06510_ (
    .a(\DFF_335.Q ),
    .b(\DFF_381.Q ),
    .y(_01638_)
  );
  al_nor2 _06511_ (
    .a(\DFF_1077.Q ),
    .b(\DFF_335.Q ),
    .y(_01639_)
  );
  al_mux2l _06512_ (
    .a(_01638_),
    .b(_01639_),
    .s(_00890_),
    .y(_01640_)
  );
  al_nand3 _06513_ (
    .a(\DFF_405.Q ),
    .b(\DFF_1334.Q ),
    .c(_01640_),
    .y(_01641_)
  );
  al_and2 _06514_ (
    .a(_01641_),
    .b(_01637_),
    .y(_01642_)
  );
  al_nand3fft _06515_ (
    .a(_01630_),
    .b(_01632_),
    .c(_01642_),
    .y(_01643_)
  );
  al_oai21ftf _06516_ (
    .a(_01629_),
    .b(_01632_),
    .c(\DFF_1077.Q ),
    .y(_01644_)
  );
  al_and2 _06517_ (
    .a(g35),
    .b(_01644_),
    .y(_01645_)
  );
  al_aoi21 _06518_ (
    .a(_01645_),
    .b(_01643_),
    .c(_01627_),
    .y(\DFF_1077.D )
  );
  al_inv _06519_ (
    .a(\DFF_111.Q ),
    .y(_01646_)
  );
  al_nand3fft _06520_ (
    .a(\DFF_759.Q ),
    .b(_01646_),
    .c(_01125_),
    .y(_01647_)
  );
  al_aoi21ftf _06521_ (
    .a(\DFF_973.Q ),
    .b(_01647_),
    .c(g35),
    .y(_01648_)
  );
  al_oai21 _06522_ (
    .a(_01131_),
    .b(_01647_),
    .c(_01648_),
    .y(_01649_)
  );
  al_ao21ftf _06523_ (
    .a(g35),
    .b(\DFF_1172.Q ),
    .c(_01649_),
    .y(\DFF_973.D )
  );
  al_nand2ft _06524_ (
    .a(g35),
    .b(\DFF_210.Q ),
    .y(_01650_)
  );
  al_ao21ftf _06525_ (
    .a(\DFF_1387.Q ),
    .b(g35),
    .c(_01650_),
    .y(\DFF_1387.D )
  );
  al_oa21ftt _06526_ (
    .a(g35),
    .b(\DFF_548.Q ),
    .c(\DFF_1385.Q ),
    .y(\DFF_631.D )
  );
  al_nand3 _06527_ (
    .a(\DFF_792.Q ),
    .b(_00673_),
    .c(_00009_),
    .y(_01651_)
  );
  al_and2ft _06528_ (
    .a(\DFF_1346.Q ),
    .b(\DFF_926.Q ),
    .y(_01652_)
  );
  al_nand2ft _06529_ (
    .a(\DFF_926.Q ),
    .b(\DFF_1346.Q ),
    .y(_01653_)
  );
  al_nand2ft _06530_ (
    .a(_01652_),
    .b(_01653_),
    .y(_01654_)
  );
  al_mux2l _06531_ (
    .a(\DFF_1121.Q ),
    .b(_01654_),
    .s(_01651_),
    .y(_01655_)
  );
  al_mux2h _06532_ (
    .a(\DFF_1346.Q ),
    .b(_01655_),
    .s(g35),
    .y(\DFF_1121.D )
  );
  al_nor2 _06533_ (
    .a(\DFF_741.Q ),
    .b(g35),
    .y(_01656_)
  );
  al_mux2h _06534_ (
    .a(_01631_),
    .b(_01628_),
    .s(\DFF_741.Q ),
    .y(_01657_)
  );
  al_nand3ftt _06535_ (
    .a(_01657_),
    .b(\DFF_1309.Q ),
    .c(_01642_),
    .y(_01658_)
  );
  al_aoi21ftf _06536_ (
    .a(\DFF_1309.Q ),
    .b(_01657_),
    .c(g35),
    .y(_01659_)
  );
  al_aoi21 _06537_ (
    .a(_01659_),
    .b(_01658_),
    .c(_01656_),
    .y(\DFF_1309.D )
  );
  al_inv _06538_ (
    .a(\DFF_635.Q ),
    .y(_01660_)
  );
  al_or2 _06539_ (
    .a(\DFF_412.Q ),
    .b(\DFF_452.Q ),
    .y(_01661_)
  );
  al_nor3ftt _06540_ (
    .a(\DFF_62.Q ),
    .b(_01661_),
    .c(_00008_),
    .y(_01662_)
  );
  al_aoi21 _06541_ (
    .a(_00456_),
    .b(_01662_),
    .c(_01660_),
    .y(_01663_)
  );
  al_and3 _06542_ (
    .a(\DFF_123.Q ),
    .b(\DFF_1005.Q ),
    .c(_00394_),
    .y(_01664_)
  );
  al_nand2 _06543_ (
    .a(_01664_),
    .b(_01663_),
    .y(_01665_)
  );
  al_nand2 _06544_ (
    .a(\DFF_897.Q ),
    .b(\DFF_400.Q ),
    .y(_01666_)
  );
  al_nor2 _06545_ (
    .a(\DFF_897.Q ),
    .b(\DFF_400.Q ),
    .y(_01667_)
  );
  al_nand2ft _06546_ (
    .a(_01667_),
    .b(_01666_),
    .y(_01668_)
  );
  al_mux2l _06547_ (
    .a(\DFF_52.Q ),
    .b(_01668_),
    .s(_01665_),
    .y(_01669_)
  );
  al_mux2h _06548_ (
    .a(\DFF_897.Q ),
    .b(_01669_),
    .s(g35),
    .y(\DFF_52.D )
  );
  al_or3 _06549_ (
    .a(g73),
    .b(g72),
    .c(\DFF_706.Q ),
    .y(_01670_)
  );
  al_aoi21 _06550_ (
    .a(g35),
    .b(_01670_),
    .c(\DFF_491.Q ),
    .y(_01671_)
  );
  al_or3 _06551_ (
    .a(\DFF_724.Q ),
    .b(\DFF_1349.Q ),
    .c(_00605_),
    .y(_01672_)
  );
  al_nand3 _06552_ (
    .a(\DFF_808.Q ),
    .b(\DFF_121.Q ),
    .c(\DFF_38.Q ),
    .y(_01673_)
  );
  al_ao21ftf _06553_ (
    .a(_01670_),
    .b(_01673_),
    .c(_01672_),
    .y(_01674_)
  );
  al_aoi21 _06554_ (
    .a(g35),
    .b(_01674_),
    .c(_01671_),
    .y(\DFF_228.D )
  );
  al_and3fft _06555_ (
    .a(_00066_),
    .b(_01424_),
    .c(_00503_),
    .y(_01675_)
  );
  al_nand2ft _06556_ (
    .a(g35),
    .b(\DFF_687.Q ),
    .y(_01676_)
  );
  al_nand3ftt _06557_ (
    .a(\DFF_250.Q ),
    .b(\DFF_929.Q ),
    .c(g35),
    .y(_01677_)
  );
  al_or3fft _06558_ (
    .a(_01676_),
    .b(_01677_),
    .c(_01675_),
    .y(\DFF_1225.D )
  );
  al_inv _06559_ (
    .a(\DFF_1147.Q ),
    .y(_01678_)
  );
  al_and3 _06560_ (
    .a(\DFF_850.Q ),
    .b(\DFF_915.Q ),
    .c(_01034_),
    .y(_01679_)
  );
  al_and3 _06561_ (
    .a(\DFF_1105.Q ),
    .b(\DFF_940.Q ),
    .c(_01679_),
    .y(_01680_)
  );
  al_inv _06562_ (
    .a(\DFF_1105.Q ),
    .y(_01681_)
  );
  al_nand3fft _06563_ (
    .a(\DFF_850.Q ),
    .b(\DFF_915.Q ),
    .c(_01035_),
    .y(_01682_)
  );
  al_and3fft _06564_ (
    .a(\DFF_940.Q ),
    .b(_01682_),
    .c(_01681_),
    .y(_01683_)
  );
  al_oai21ttf _06565_ (
    .a(_01683_),
    .b(_01680_),
    .c(_01678_),
    .y(_01684_)
  );
  al_nand3 _06566_ (
    .a(\DFF_1147.Q ),
    .b(_01039_),
    .c(_01041_),
    .y(_01685_)
  );
  al_nand3fft _06567_ (
    .a(_01683_),
    .b(_01680_),
    .c(_01685_),
    .y(_01686_)
  );
  al_nand3 _06568_ (
    .a(g35),
    .b(_01686_),
    .c(_01684_),
    .y(_01687_)
  );
  al_ao21ftf _06569_ (
    .a(g35),
    .b(\DFF_940.Q ),
    .c(_01687_),
    .y(\DFF_1147.D )
  );
  al_and3ftt _06570_ (
    .a(\DFF_849.Q ),
    .b(\DFF_894.Q ),
    .c(\DFF_609.Q ),
    .y(_01688_)
  );
  al_aoi21ttf _06571_ (
    .a(_01688_),
    .b(_01662_),
    .c(\DFF_107.Q ),
    .y(_01689_)
  );
  al_nor3fft _06572_ (
    .a(\DFF_599.Q ),
    .b(\DFF_101.Q ),
    .c(_00407_),
    .y(_01690_)
  );
  al_nand2 _06573_ (
    .a(_01690_),
    .b(_01689_),
    .y(_01691_)
  );
  al_or3fft _06574_ (
    .a(\DFF_1018.Q ),
    .b(g35),
    .c(_01691_),
    .y(_01692_)
  );
  al_or2 _06575_ (
    .a(\DFF_1079.Q ),
    .b(g35),
    .y(_01693_)
  );
  al_and2ft _06576_ (
    .a(\DFF_1018.Q ),
    .b(g35),
    .y(_01694_)
  );
  al_ao21ttf _06577_ (
    .a(_01690_),
    .b(_01689_),
    .c(_01694_),
    .y(_01695_)
  );
  al_and3 _06578_ (
    .a(_01693_),
    .b(_01695_),
    .c(_01692_),
    .y(\DFF_1018.D )
  );
  al_ao21ttf _06579_ (
    .a(_00821_),
    .b(_00822_),
    .c(_00829_),
    .y(_01696_)
  );
  al_and3 _06580_ (
    .a(\DFF_1039.Q ),
    .b(g35),
    .c(_01696_),
    .y(_01697_)
  );
  al_nand2ft _06581_ (
    .a(_00824_),
    .b(_00826_),
    .y(_01698_)
  );
  al_ao21ftf _06582_ (
    .a(\DFF_1343.Q ),
    .b(_00962_),
    .c(_01698_),
    .y(_01699_)
  );
  al_oa21 _06583_ (
    .a(\DFF_408.Q ),
    .b(\DFF_990.Q ),
    .c(g35),
    .y(_01700_)
  );
  al_ao21 _06584_ (
    .a(_01700_),
    .b(_01699_),
    .c(_01697_),
    .y(\DFF_1039.D )
  );
  al_and2ft _06585_ (
    .a(\DFF_910.Q ),
    .b(\DFF_575.Q ),
    .y(_01701_)
  );
  al_and2 _06586_ (
    .a(\DFF_244.Q ),
    .b(\DFF_958.Q ),
    .y(_01702_)
  );
  al_nand3 _06587_ (
    .a(_00499_),
    .b(_01701_),
    .c(_01702_),
    .y(_01703_)
  );
  al_ao21 _06588_ (
    .a(_01701_),
    .b(_01702_),
    .c(\DFF_219.Q ),
    .y(_01704_)
  );
  al_nand3 _06589_ (
    .a(g35),
    .b(_01704_),
    .c(_01703_),
    .y(_01705_)
  );
  al_ao21ftf _06590_ (
    .a(g35),
    .b(\DFF_1355.Q ),
    .c(_01705_),
    .y(\DFF_219.D )
  );
  al_nor2 _06591_ (
    .a(\DFF_1127.Q ),
    .b(g35),
    .y(_01706_)
  );
  al_nand3 _06592_ (
    .a(\DFF_1181.Q ),
    .b(_00604_),
    .c(_00339_),
    .y(_01707_)
  );
  al_nand3 _06593_ (
    .a(\DFF_1127.Q ),
    .b(_00721_),
    .c(_01707_),
    .y(_01708_)
  );
  al_oa21ftf _06594_ (
    .a(\DFF_646.Q ),
    .b(_00721_),
    .c(_00066_),
    .y(_01709_)
  );
  al_aoi21 _06595_ (
    .a(_01709_),
    .b(_01708_),
    .c(_01706_),
    .y(\DFF_646.D )
  );
  al_and2ft _06596_ (
    .a(g35),
    .b(\DFF_804.Q ),
    .y(_01710_)
  );
  al_nand2ft _06597_ (
    .a(\DFF_637.Q ),
    .b(\DFF_804.Q ),
    .y(_01711_)
  );
  al_nand2ft _06598_ (
    .a(\DFF_804.Q ),
    .b(\DFF_637.Q ),
    .y(_01712_)
  );
  al_or3fft _06599_ (
    .a(_01711_),
    .b(_01712_),
    .c(_01397_),
    .y(_01713_)
  );
  al_aoi21 _06600_ (
    .a(_01435_),
    .b(_01397_),
    .c(_00066_),
    .y(_01714_)
  );
  al_ao21 _06601_ (
    .a(_01713_),
    .b(_01714_),
    .c(_01710_),
    .y(\DFF_928.D )
  );
  al_and2ft _06602_ (
    .a(g35),
    .b(\DFF_522.Q ),
    .y(_01715_)
  );
  al_ao21 _06603_ (
    .a(\DFF_522.Q ),
    .b(\DFF_54.Q ),
    .c(\DFF_271.Q ),
    .y(_01716_)
  );
  al_nor3fft _06604_ (
    .a(g35),
    .b(_01716_),
    .c(_00365_),
    .y(_01717_)
  );
  al_ao21 _06605_ (
    .a(_01717_),
    .b(_01359_),
    .c(_01715_),
    .y(\DFF_271.D )
  );
  al_and2 _06606_ (
    .a(\DFF_190.Q ),
    .b(g35),
    .y(\DFF_190.D )
  );
  al_and2 _06607_ (
    .a(\DFF_383.Q ),
    .b(\DFF_129.Q ),
    .y(_01718_)
  );
  al_and3 _06608_ (
    .a(\DFF_911.Q ),
    .b(\DFF_1209.Q ),
    .c(_01718_),
    .y(_01719_)
  );
  al_or2 _06609_ (
    .a(\DFF_813.Q ),
    .b(_01719_),
    .y(_01720_)
  );
  al_nand2 _06610_ (
    .a(\DFF_813.Q ),
    .b(_01719_),
    .y(_01721_)
  );
  al_aoi21 _06611_ (
    .a(_01721_),
    .b(_01720_),
    .c(_00066_),
    .y(_01722_)
  );
  al_nand3fft _06612_ (
    .a(\DFF_79.Q ),
    .b(_00066_),
    .c(_00998_),
    .y(_01723_)
  );
  al_ao21ftf _06613_ (
    .a(_01722_),
    .b(\DFF_79.Q ),
    .c(_01723_),
    .y(\DFF_813.D )
  );
  al_or2 _06614_ (
    .a(\DFF_294.Q ),
    .b(\DFF_532.Q ),
    .y(_01724_)
  );
  al_nand3 _06615_ (
    .a(\DFF_240.Q ),
    .b(g35),
    .c(_01724_),
    .y(_01725_)
  );
  al_oai21ftt _06616_ (
    .a(\DFF_654.Q ),
    .b(\DFF_240.Q ),
    .c(g35),
    .y(_01726_)
  );
  al_nor2 _06617_ (
    .a(g35),
    .b(\DFF_294.Q ),
    .y(_01727_)
  );
  al_ao21ftf _06618_ (
    .a(_01727_),
    .b(_01726_),
    .c(_01725_),
    .y(\DFF_654.D )
  );
  al_ao21 _06619_ (
    .a(\DFF_902.Q ),
    .b(_00872_),
    .c(\DFF_112.Q ),
    .y(_01728_)
  );
  al_nand3ftt _06620_ (
    .a(_01599_),
    .b(_01728_),
    .c(_01607_),
    .y(_01729_)
  );
  al_ao21ftf _06621_ (
    .a(g35),
    .b(\DFF_902.Q ),
    .c(_01729_),
    .y(\DFF_112.D )
  );
  al_or3 _06622_ (
    .a(\DFF_792.Q ),
    .b(\DFF_107.Q ),
    .c(\DFF_699.Q ),
    .y(_01730_)
  );
  al_and2ft _06623_ (
    .a(_00460_),
    .b(_00745_),
    .y(_01731_)
  );
  al_and3ftt _06624_ (
    .a(_01730_),
    .b(g35),
    .c(_01731_),
    .y(\DFF_792.D )
  );
  al_and3fft _06625_ (
    .a(\DFF_1364.Q ),
    .b(_00451_),
    .c(_00542_),
    .y(_01732_)
  );
  al_and3ftt _06626_ (
    .a(\DFF_893.Q ),
    .b(\DFF_284.Q ),
    .c(\DFF_962.Q ),
    .y(_01733_)
  );
  al_aoi21 _06627_ (
    .a(\DFF_302.Q ),
    .b(_00561_),
    .c(_01733_),
    .y(_01734_)
  );
  al_and3 _06628_ (
    .a(\DFF_233.Q ),
    .b(\DFF_893.Q ),
    .c(\DFF_962.Q ),
    .y(_01735_)
  );
  al_aoi21 _06629_ (
    .a(\DFF_1112.Q ),
    .b(_00575_),
    .c(_01735_),
    .y(_01736_)
  );
  al_ao21ttf _06630_ (
    .a(_01734_),
    .b(_01736_),
    .c(_01732_),
    .y(_01737_)
  );
  al_nand3ftt _06631_ (
    .a(\DFF_1082.Q ),
    .b(\DFF_893.Q ),
    .c(\DFF_962.Q ),
    .y(_01738_)
  );
  al_aoi21ftf _06632_ (
    .a(\DFF_989.Q ),
    .b(_00561_),
    .c(_01738_),
    .y(_01739_)
  );
  al_or3ftt _06633_ (
    .a(\DFF_962.Q ),
    .b(\DFF_893.Q ),
    .c(\DFF_406.Q ),
    .y(_01740_)
  );
  al_aoi21ftf _06634_ (
    .a(\DFF_37.Q ),
    .b(_00575_),
    .c(_01740_),
    .y(_01741_)
  );
  al_ao21 _06635_ (
    .a(_01739_),
    .b(_01741_),
    .c(_01732_),
    .y(_01742_)
  );
  al_nand3 _06636_ (
    .a(g35),
    .b(_01737_),
    .c(_01742_),
    .y(_01743_)
  );
  al_ao21ftf _06637_ (
    .a(g35),
    .b(\DFF_1112.Q ),
    .c(_01743_),
    .y(\DFF_576.D )
  );
  al_and2ft _06638_ (
    .a(\DFF_244.Q ),
    .b(\DFF_958.Q ),
    .y(_01744_)
  );
  al_nor2 _06639_ (
    .a(\DFF_575.Q ),
    .b(\DFF_910.Q ),
    .y(_01745_)
  );
  al_nand3 _06640_ (
    .a(_00499_),
    .b(_01744_),
    .c(_01745_),
    .y(_01746_)
  );
  al_ao21 _06641_ (
    .a(_01744_),
    .b(_01745_),
    .c(\DFF_51.Q ),
    .y(_01747_)
  );
  al_nand3 _06642_ (
    .a(g35),
    .b(_01747_),
    .c(_01746_),
    .y(_01748_)
  );
  al_ao21ftf _06643_ (
    .a(g35),
    .b(\DFF_627.Q ),
    .c(_01748_),
    .y(\DFF_51.D )
  );
  al_and2ft _06644_ (
    .a(g35),
    .b(\DFF_139.Q ),
    .y(_01749_)
  );
  al_and3 _06645_ (
    .a(_00391_),
    .b(_00393_),
    .c(_00386_),
    .y(_01750_)
  );
  al_nand3 _06646_ (
    .a(_00587_),
    .b(_01663_),
    .c(_01750_),
    .y(_01751_)
  );
  al_ao21 _06647_ (
    .a(\DFF_139.Q ),
    .b(_01663_),
    .c(\DFF_118.Q ),
    .y(_01752_)
  );
  al_nand3 _06648_ (
    .a(\DFF_118.Q ),
    .b(\DFF_139.Q ),
    .c(_01663_),
    .y(_01753_)
  );
  al_and3 _06649_ (
    .a(g35),
    .b(_01753_),
    .c(_01752_),
    .y(_01754_)
  );
  al_ao21 _06650_ (
    .a(_01751_),
    .b(_01754_),
    .c(_01749_),
    .y(\DFF_118.D )
  );
  al_inv _06651_ (
    .a(\DFF_1413.Q ),
    .y(_01755_)
  );
  al_nand3fft _06652_ (
    .a(_01755_),
    .b(\DFF_671.Q ),
    .c(_01150_),
    .y(_01756_)
  );
  al_aoi21 _06653_ (
    .a(_01518_),
    .b(_01756_),
    .c(_00066_),
    .y(_01757_)
  );
  al_oai21 _06654_ (
    .a(_01153_),
    .b(_01756_),
    .c(_01757_),
    .y(_01758_)
  );
  al_ao21ftf _06655_ (
    .a(g35),
    .b(\DFF_255.Q ),
    .c(_01758_),
    .y(\DFF_1394.D )
  );
  al_ao21 _06656_ (
    .a(\DFF_1324.Q ),
    .b(\DFF_891.Q ),
    .c(\DFF_1361.Q ),
    .y(_01759_)
  );
  al_and2 _06657_ (
    .a(\DFF_434.Q ),
    .b(g35),
    .y(_01760_)
  );
  al_and3 _06658_ (
    .a(\DFF_1361.Q ),
    .b(\DFF_1324.Q ),
    .c(\DFF_891.Q ),
    .y(_01761_)
  );
  al_or3fft _06659_ (
    .a(_01759_),
    .b(_01760_),
    .c(_01761_),
    .y(_01762_)
  );
  al_ao21ftf _06660_ (
    .a(g35),
    .b(\DFF_1324.Q ),
    .c(_01762_),
    .y(\DFF_1361.D )
  );
  al_and2 _06661_ (
    .a(\DFF_1150.Q ),
    .b(\DFF_1068.Q ),
    .y(_01763_)
  );
  al_and2 _06662_ (
    .a(\DFF_410.Q ),
    .b(\DFF_584.Q ),
    .y(_01764_)
  );
  al_nand3 _06663_ (
    .a(_00499_),
    .b(_01763_),
    .c(_01764_),
    .y(_01765_)
  );
  al_ao21 _06664_ (
    .a(_01763_),
    .b(_01764_),
    .c(\DFF_779.Q ),
    .y(_01766_)
  );
  al_nand3 _06665_ (
    .a(g35),
    .b(_01765_),
    .c(_01766_),
    .y(_01767_)
  );
  al_ao21ftf _06666_ (
    .a(g35),
    .b(\DFF_291.Q ),
    .c(_01767_),
    .y(\DFF_779.D )
  );
  al_or3 _06667_ (
    .a(\DFF_925.Q ),
    .b(\DFF_653.Q ),
    .c(\DFF_104.Q ),
    .y(_01768_)
  );
  al_nand3ftt _06668_ (
    .a(_01768_),
    .b(_00499_),
    .c(_01170_),
    .y(_01769_)
  );
  al_ao21ftt _06669_ (
    .a(_01768_),
    .b(_01170_),
    .c(\DFF_945.Q ),
    .y(_01770_)
  );
  al_nand3 _06670_ (
    .a(g35),
    .b(_01769_),
    .c(_01770_),
    .y(_01771_)
  );
  al_ao21ftf _06671_ (
    .a(g35),
    .b(\DFF_314.Q ),
    .c(_01771_),
    .y(\DFF_945.D )
  );
  al_and2 _06672_ (
    .a(\DFF_575.Q ),
    .b(\DFF_910.Q ),
    .y(_01772_)
  );
  al_and2ft _06673_ (
    .a(\DFF_958.Q ),
    .b(\DFF_244.Q ),
    .y(_01773_)
  );
  al_nand3 _06674_ (
    .a(_00499_),
    .b(_01772_),
    .c(_01773_),
    .y(_01774_)
  );
  al_ao21 _06675_ (
    .a(_01773_),
    .b(_01772_),
    .c(\DFF_895.Q ),
    .y(_01775_)
  );
  al_nand3 _06676_ (
    .a(g35),
    .b(_01775_),
    .c(_01774_),
    .y(_01776_)
  );
  al_ao21ftf _06677_ (
    .a(g35),
    .b(\DFF_1007.Q ),
    .c(_01776_),
    .y(\DFF_895.D )
  );
  al_nand3 _06678_ (
    .a(_00499_),
    .b(_01070_),
    .c(_01497_),
    .y(_01777_)
  );
  al_ao21 _06679_ (
    .a(_01070_),
    .b(_01497_),
    .c(\DFF_105.Q ),
    .y(_01778_)
  );
  al_nand3 _06680_ (
    .a(g35),
    .b(_01778_),
    .c(_01777_),
    .y(_01779_)
  );
  al_ao21ftf _06681_ (
    .a(g35),
    .b(\DFF_108.Q ),
    .c(_01779_),
    .y(\DFF_105.D )
  );
  al_oa21ftt _06682_ (
    .a(g35),
    .b(\DFF_969.Q ),
    .c(\DFF_3.Q ),
    .y(_01780_)
  );
  al_nand2ft _06683_ (
    .a(\DFF_975.Q ),
    .b(\DFF_907.Q ),
    .y(_01781_)
  );
  al_oa21ftf _06684_ (
    .a(\DFF_907.Q ),
    .b(\DFF_1113.Q ),
    .c(\DFF_969.Q ),
    .y(_01782_)
  );
  al_ao21ftf _06685_ (
    .a(\DFF_3.Q ),
    .b(_01782_),
    .c(_01781_),
    .y(_01783_)
  );
  al_ao21 _06686_ (
    .a(g35),
    .b(_01783_),
    .c(_01780_),
    .y(\DFF_969.D )
  );
  al_nand3 _06687_ (
    .a(\DFF_402.Q ),
    .b(_01615_),
    .c(_00641_),
    .y(_01784_)
  );
  al_aoi21ftf _06688_ (
    .a(\DFF_1097.Q ),
    .b(_01784_),
    .c(g35),
    .y(_01785_)
  );
  al_ao21ftf _06689_ (
    .a(_01784_),
    .b(_01618_),
    .c(_01785_),
    .y(_01786_)
  );
  al_ao21ftf _06690_ (
    .a(g35),
    .b(\DFF_61.Q ),
    .c(_01786_),
    .y(\DFF_1097.D )
  );
  al_and2ft _06691_ (
    .a(\DFF_1150.Q ),
    .b(\DFF_1068.Q ),
    .y(_01787_)
  );
  al_nand3 _06692_ (
    .a(_00499_),
    .b(_01764_),
    .c(_01787_),
    .y(_01788_)
  );
  al_ao21 _06693_ (
    .a(_01787_),
    .b(_01764_),
    .c(\DFF_378.Q ),
    .y(_01789_)
  );
  al_nand3 _06694_ (
    .a(g35),
    .b(_01789_),
    .c(_01788_),
    .y(_01790_)
  );
  al_ao21ftf _06695_ (
    .a(g35),
    .b(\DFF_1120.Q ),
    .c(_01790_),
    .y(\DFF_378.D )
  );
  al_oa21ftt _06696_ (
    .a(\DFF_827.Q ),
    .b(\DFF_57.Q ),
    .c(g35),
    .y(_01791_)
  );
  al_nand3fft _06697_ (
    .a(\DFF_1377.Q ),
    .b(\DFF_827.Q ),
    .c(g35),
    .y(_01792_)
  );
  al_aoi21ttf _06698_ (
    .a(_01792_),
    .b(_01791_),
    .c(\DFF_1249.Q ),
    .y(\DFF_1318.D )
  );
  al_nand3ftt _06699_ (
    .a(_01547_),
    .b(_00499_),
    .c(_00509_),
    .y(_01793_)
  );
  al_ao21ftt _06700_ (
    .a(_01547_),
    .b(_00509_),
    .c(\DFF_1174.Q ),
    .y(_01794_)
  );
  al_nand3 _06701_ (
    .a(g35),
    .b(_01793_),
    .c(_01794_),
    .y(_01795_)
  );
  al_ao21ftf _06702_ (
    .a(g35),
    .b(\DFF_1068.Q ),
    .c(_01795_),
    .y(\DFF_1174.D )
  );
  al_nand2ft _06703_ (
    .a(\DFF_1054.Q ),
    .b(\DFF_1127.Q ),
    .y(_01796_)
  );
  al_and3fft _06704_ (
    .a(_01796_),
    .b(_00725_),
    .c(_00721_),
    .y(_01797_)
  );
  al_ao21ftt _06705_ (
    .a(_01796_),
    .b(_00721_),
    .c(\DFF_735.Q ),
    .y(_01798_)
  );
  al_or3fft _06706_ (
    .a(g35),
    .b(_01798_),
    .c(_01797_),
    .y(_01799_)
  );
  al_ao21ftf _06707_ (
    .a(g35),
    .b(\DFF_864.Q ),
    .c(_01799_),
    .y(\DFF_735.D )
  );
  al_or2ft _06708_ (
    .a(\DFF_243.Q ),
    .b(_00378_),
    .y(_01800_)
  );
  al_inv _06709_ (
    .a(\DFF_29.Q ),
    .y(_01801_)
  );
  al_and2ft _06710_ (
    .a(\DFF_955.Q ),
    .b(g35),
    .y(_01802_)
  );
  al_ao21ftf _06711_ (
    .a(_01801_),
    .b(_01802_),
    .c(_01016_),
    .y(_01803_)
  );
  al_and3ftt _06712_ (
    .a(_01802_),
    .b(_01801_),
    .c(_01016_),
    .y(_01804_)
  );
  al_aoi21 _06713_ (
    .a(_01800_),
    .b(_01803_),
    .c(_01804_),
    .y(\DFF_243.D )
  );
  al_nor3ftt _06714_ (
    .a(\DFF_1138.Q ),
    .b(_00499_),
    .c(_00358_),
    .y(_01805_)
  );
  al_oa21ftt _06715_ (
    .a(\DFF_1138.Q ),
    .b(_00358_),
    .c(_00499_),
    .y(_01806_)
  );
  al_nor3ftt _06716_ (
    .a(g35),
    .b(_01805_),
    .c(_01806_),
    .y(\DFF_1138.D )
  );
  al_ao21 _06717_ (
    .a(\DFF_385.Q ),
    .b(\DFF_393.Q ),
    .c(\DFF_519.Q ),
    .y(_01807_)
  );
  al_nand3ftt _06718_ (
    .a(_01393_),
    .b(_01807_),
    .c(_01442_),
    .y(_01808_)
  );
  al_ao21ftf _06719_ (
    .a(g35),
    .b(\DFF_385.Q ),
    .c(_01808_),
    .y(\DFF_519.D )
  );
  al_inv _06720_ (
    .a(\DFF_646.Q ),
    .y(_01809_)
  );
  al_inv _06721_ (
    .a(\DFF_1054.Q ),
    .y(_01810_)
  );
  al_nand3fft _06722_ (
    .a(_01809_),
    .b(_01810_),
    .c(_00721_),
    .y(_01811_)
  );
  al_aoi21ftf _06723_ (
    .a(\DFF_1180.Q ),
    .b(_01811_),
    .c(g35),
    .y(_01812_)
  );
  al_oai21 _06724_ (
    .a(_00725_),
    .b(_01811_),
    .c(_01812_),
    .y(_01813_)
  );
  al_ao21ftf _06725_ (
    .a(g35),
    .b(\DFF_735.Q ),
    .c(_01813_),
    .y(\DFF_1180.D )
  );
  al_mux2l _06726_ (
    .a(g124),
    .b(g120),
    .s(\DFF_673.Q ),
    .y(_01814_)
  );
  al_mux2h _06727_ (
    .a(\DFF_201.Q ),
    .b(_01814_),
    .s(g35),
    .y(\DFF_1230.D )
  );
  al_mux2l _06728_ (
    .a(\DFF_955.Q ),
    .b(\DFF_29.Q ),
    .s(_01016_),
    .y(\DFF_29.D )
  );
  al_and2 _06729_ (
    .a(\DFF_860.Q ),
    .b(_01761_),
    .y(_01815_)
  );
  al_or2 _06730_ (
    .a(\DFF_860.Q ),
    .b(_01761_),
    .y(_01816_)
  );
  al_oai21ftt _06731_ (
    .a(_01816_),
    .b(_01815_),
    .c(_01760_),
    .y(_01817_)
  );
  al_aoi21ftf _06732_ (
    .a(\DFF_1361.Q ),
    .b(_00066_),
    .c(_01817_),
    .y(\DFF_860.D )
  );
  al_inv _06733_ (
    .a(\DFF_454.Q ),
    .y(_01818_)
  );
  al_and2 _06734_ (
    .a(\DFF_1275.Q ),
    .b(\DFF_454.Q ),
    .y(_01819_)
  );
  al_mux2l _06735_ (
    .a(_01818_),
    .b(_01819_),
    .s(_01317_),
    .y(_01820_)
  );
  al_mux2h _06736_ (
    .a(\DFF_954.Q ),
    .b(_01820_),
    .s(g35),
    .y(\DFF_454.D )
  );
  al_mux2l _06737_ (
    .a(\DFF_236.Q ),
    .b(\DFF_69.Q ),
    .s(g35),
    .y(\DFF_236.D )
  );
  al_mux2l _06738_ (
    .a(\DFF_1126.Q ),
    .b(\DFF_238.Q ),
    .s(_01053_),
    .y(_01821_)
  );
  al_mux2h _06739_ (
    .a(\DFF_1250.Q ),
    .b(_01821_),
    .s(g35),
    .y(\DFF_1126.D )
  );
  al_inv _06740_ (
    .a(\DFF_1016.Q ),
    .y(_01822_)
  );
  al_ao21ftf _06741_ (
    .a(\DFF_1399.Q ),
    .b(_00342_),
    .c(_00605_),
    .y(_01823_)
  );
  al_nand3ftt _06742_ (
    .a(\DFF_184.Q ),
    .b(\DFF_615.Q ),
    .c(_01823_),
    .y(_01824_)
  );
  al_ao21ftf _06743_ (
    .a(_01822_),
    .b(\DFF_549.Q ),
    .c(_01824_),
    .y(_01825_)
  );
  al_or3ftt _06744_ (
    .a(g35),
    .b(\DFF_965.Q ),
    .c(_01825_),
    .y(\DFF_549.D )
  );
  al_inv _06745_ (
    .a(\DFF_667.Q ),
    .y(_01826_)
  );
  al_nand3fft _06746_ (
    .a(_01826_),
    .b(\DFF_1390.Q ),
    .c(_01605_),
    .y(_01827_)
  );
  al_ao21ftf _06747_ (
    .a(\DFF_1019.Q ),
    .b(\DFF_667.Q ),
    .c(_01348_),
    .y(_01828_)
  );
  al_ao21 _06748_ (
    .a(\DFF_1390.Q ),
    .b(_01828_),
    .c(_00066_),
    .y(_01829_)
  );
  al_oai21ftf _06749_ (
    .a(_01348_),
    .b(_01827_),
    .c(_01829_),
    .y(_01830_)
  );
  al_aoi21ftf _06750_ (
    .a(\DFF_1044.Q ),
    .b(_00066_),
    .c(_01830_),
    .y(\DFF_1390.D )
  );
  al_or3fft _06751_ (
    .a(g35),
    .b(_01490_),
    .c(_01488_),
    .y(g26875)
  );
  al_inv _06752_ (
    .a(_01760_),
    .y(_01831_)
  );
  al_and2 _06753_ (
    .a(\DFF_154.Q ),
    .b(\DFF_411.Q ),
    .y(_01832_)
  );
  al_and3 _06754_ (
    .a(\DFF_860.Q ),
    .b(_01761_),
    .c(_01832_),
    .y(_01833_)
  );
  al_and3 _06755_ (
    .a(\DFF_551.Q ),
    .b(\DFF_351.Q ),
    .c(_01833_),
    .y(_01834_)
  );
  al_ao21 _06756_ (
    .a(\DFF_551.Q ),
    .b(_01833_),
    .c(\DFF_351.Q ),
    .y(_01835_)
  );
  al_ao21ftt _06757_ (
    .a(_01834_),
    .b(_01835_),
    .c(_01831_),
    .y(_01836_)
  );
  al_aoi21ftf _06758_ (
    .a(\DFF_551.Q ),
    .b(_00066_),
    .c(_01836_),
    .y(\DFF_351.D )
  );
  al_inv _06759_ (
    .a(_01175_),
    .y(_01837_)
  );
  al_ao21 _06760_ (
    .a(\DFF_175.Q ),
    .b(_01178_),
    .c(\DFF_28.Q ),
    .y(_01838_)
  );
  al_nand3fft _06761_ (
    .a(_01837_),
    .b(_01179_),
    .c(_01838_),
    .y(_01839_)
  );
  al_ao21ftf _06762_ (
    .a(g35),
    .b(\DFF_175.Q ),
    .c(_01839_),
    .y(\DFF_28.D )
  );
  al_nor2 _06763_ (
    .a(\DFF_598.Q ),
    .b(\DFF_68.Q ),
    .y(_01840_)
  );
  al_nand3ftt _06764_ (
    .a(_01311_),
    .b(_00499_),
    .c(_01840_),
    .y(_01841_)
  );
  al_ao21ftt _06765_ (
    .a(_01311_),
    .b(_01840_),
    .c(\DFF_638.Q ),
    .y(_01842_)
  );
  al_nand3 _06766_ (
    .a(g35),
    .b(_01841_),
    .c(_01842_),
    .y(_01843_)
  );
  al_ao21ftf _06767_ (
    .a(g35),
    .b(\DFF_598.Q ),
    .c(_01843_),
    .y(\DFF_638.D )
  );
  al_and2ft _06768_ (
    .a(\DFF_713.Q ),
    .b(\DFF_402.Q ),
    .y(_01844_)
  );
  al_nand3 _06769_ (
    .a(_00444_),
    .b(_01844_),
    .c(_00758_),
    .y(_01845_)
  );
  al_ao21 _06770_ (
    .a(_00444_),
    .b(_00758_),
    .c(\DFF_487.Q ),
    .y(_01846_)
  );
  al_nand3 _06771_ (
    .a(g35),
    .b(_01845_),
    .c(_01846_),
    .y(_01847_)
  );
  al_ao21ftf _06772_ (
    .a(g35),
    .b(\DFF_960.Q ),
    .c(_01847_),
    .y(\DFF_487.D )
  );
  al_and2 _06773_ (
    .a(_01406_),
    .b(_00606_),
    .y(_01848_)
  );
  al_ao21ftf _06774_ (
    .a(\DFF_43.Q ),
    .b(_01848_),
    .c(g35),
    .y(_01849_)
  );
  al_and3 _06775_ (
    .a(g35),
    .b(_00999_),
    .c(_01848_),
    .y(_01850_)
  );
  al_ao21 _06776_ (
    .a(\DFF_331.Q ),
    .b(_01849_),
    .c(_01850_),
    .y(\DFF_43.D )
  );
  al_and2ft _06777_ (
    .a(g35),
    .b(\DFF_452.Q ),
    .y(_01851_)
  );
  al_nor2 _06778_ (
    .a(\DFF_412.Q ),
    .b(_01323_),
    .y(_01852_)
  );
  al_nor2ft _06779_ (
    .a(_01322_),
    .b(_01852_),
    .y(_01853_)
  );
  al_ao21 _06780_ (
    .a(_01853_),
    .b(_01325_),
    .c(_01851_),
    .y(\DFF_412.D )
  );
  al_ao21ttf _06781_ (
    .a(\DFF_354.Q ),
    .b(\DFF_605.Q ),
    .c(g35),
    .y(_01854_)
  );
  al_and2 _06782_ (
    .a(\DFF_691.Q ),
    .b(_01854_),
    .y(_01855_)
  );
  al_or3fft _06783_ (
    .a(\DFF_556.Q ),
    .b(g35),
    .c(_01855_),
    .y(_01856_)
  );
  al_aoi21ftf _06784_ (
    .a(_00066_),
    .b(\DFF_556.Q ),
    .c(_01855_),
    .y(_01857_)
  );
  al_nand2ft _06785_ (
    .a(_01857_),
    .b(_01856_),
    .y(\DFF_556.D )
  );
  al_and3 _06786_ (
    .a(_01413_),
    .b(_01414_),
    .c(_01282_),
    .y(_01858_)
  );
  al_nand2 _06787_ (
    .a(\DFF_903.Q ),
    .b(\DFF_232.Q ),
    .y(_01859_)
  );
  al_nor2 _06788_ (
    .a(\DFF_903.Q ),
    .b(\DFF_232.Q ),
    .y(_01860_)
  );
  al_nand2ft _06789_ (
    .a(_01860_),
    .b(_01859_),
    .y(_01861_)
  );
  al_mux2l _06790_ (
    .a(_01861_),
    .b(\DFF_841.Q ),
    .s(_01858_),
    .y(_01862_)
  );
  al_mux2h _06791_ (
    .a(\DFF_903.Q ),
    .b(_01862_),
    .s(g35),
    .y(\DFF_841.D )
  );
  al_nand3fft _06792_ (
    .a(\DFF_1199.Q ),
    .b(\DFF_892.Q ),
    .c(_00464_),
    .y(_01863_)
  );
  al_nand3fft _06793_ (
    .a(\DFF_1176.Q ),
    .b(\DFF_672.Q ),
    .c(_00342_),
    .y(_01864_)
  );
  al_or2ft _06794_ (
    .a(\DFF_1424.Q ),
    .b(_01864_),
    .y(_01865_)
  );
  al_ao21ftf _06795_ (
    .a(_01863_),
    .b(_01865_),
    .c(g35),
    .y(_01866_)
  );
  al_ao21ftf _06796_ (
    .a(\DFF_78.Q ),
    .b(_01863_),
    .c(_01864_),
    .y(_01867_)
  );
  al_nand3 _06797_ (
    .a(g35),
    .b(_01865_),
    .c(_01867_),
    .y(_01868_)
  );
  al_aoi21ftf _06798_ (
    .a(\DFF_1206.Q ),
    .b(_01866_),
    .c(_01868_),
    .y(\DFF_78.D )
  );
  al_inv _06799_ (
    .a(\DFF_639.Q ),
    .y(_01869_)
  );
  al_and3 _06800_ (
    .a(\DFF_1132.Q ),
    .b(\DFF_665.Q ),
    .c(_01338_),
    .y(_01870_)
  );
  al_and3 _06801_ (
    .a(\DFF_823.Q ),
    .b(\DFF_518.Q ),
    .c(_01870_),
    .y(_01871_)
  );
  al_inv _06802_ (
    .a(\DFF_823.Q ),
    .y(_01872_)
  );
  al_nand3fft _06803_ (
    .a(\DFF_1132.Q ),
    .b(\DFF_665.Q ),
    .c(_01339_),
    .y(_01873_)
  );
  al_and3fft _06804_ (
    .a(\DFF_518.Q ),
    .b(_01873_),
    .c(_01872_),
    .y(_01874_)
  );
  al_oai21ttf _06805_ (
    .a(_01874_),
    .b(_01871_),
    .c(_01869_),
    .y(_01875_)
  );
  al_nand3 _06806_ (
    .a(\DFF_639.Q ),
    .b(_01335_),
    .c(_01337_),
    .y(_01876_)
  );
  al_nand3fft _06807_ (
    .a(_01874_),
    .b(_01871_),
    .c(_01876_),
    .y(_01877_)
  );
  al_nand3 _06808_ (
    .a(g35),
    .b(_01877_),
    .c(_01875_),
    .y(_01878_)
  );
  al_ao21ftf _06809_ (
    .a(g35),
    .b(\DFF_823.Q ),
    .c(_01878_),
    .y(\DFF_639.D )
  );
  al_inv _06810_ (
    .a(\DFF_786.Q ),
    .y(_01879_)
  );
  al_ao21ftt _06811_ (
    .a(_01348_),
    .b(_00322_),
    .c(_01351_),
    .y(_01880_)
  );
  al_ao21ftf _06812_ (
    .a(_01879_),
    .b(_01349_),
    .c(_01880_),
    .y(\DFF_622.D )
  );
  al_or2ft _06813_ (
    .a(\DFF_1370.Q ),
    .b(g26801),
    .y(_01881_)
  );
  al_nand2ft _06814_ (
    .a(\DFF_1370.Q ),
    .b(g26801),
    .y(_01882_)
  );
  al_nand3 _06815_ (
    .a(g35),
    .b(_01882_),
    .c(_01881_),
    .y(_01883_)
  );
  al_aoi21ftf _06816_ (
    .a(\DFF_1121.Q ),
    .b(_00066_),
    .c(_01883_),
    .y(\DFF_1370.D )
  );
  al_inv _06817_ (
    .a(\DFF_18.Q ),
    .y(_01884_)
  );
  al_inv _06818_ (
    .a(\DFF_272.Q ),
    .y(_01885_)
  );
  al_aoi21ftf _06819_ (
    .a(\DFF_1242.Q ),
    .b(\DFF_296.Q ),
    .c(_00719_),
    .y(_01886_)
  );
  al_nand3ftt _06820_ (
    .a(\DFF_941.Q ),
    .b(\DFF_445.Q ),
    .c(\DFF_507.Q ),
    .y(_01887_)
  );
  al_ao21ttf _06821_ (
    .a(_01480_),
    .b(_00346_),
    .c(\DFF_643.Q ),
    .y(_01888_)
  );
  al_nand3 _06822_ (
    .a(_01887_),
    .b(_01886_),
    .c(_01888_),
    .y(_01889_)
  );
  al_and3 _06823_ (
    .a(_01884_),
    .b(_01885_),
    .c(_01889_),
    .y(_01890_)
  );
  al_aoi21ftf _06824_ (
    .a(_01887_),
    .b(_00528_),
    .c(_01886_),
    .y(_01891_)
  );
  al_ao21ftf _06825_ (
    .a(\DFF_828.Q ),
    .b(_01887_),
    .c(_01891_),
    .y(_01892_)
  );
  al_mux2l _06826_ (
    .a(_01892_),
    .b(\DFF_1258.Q ),
    .s(_01890_),
    .y(_01893_)
  );
  al_mux2h _06827_ (
    .a(\DFF_1114.Q ),
    .b(_01893_),
    .s(g35),
    .y(\DFF_1258.D )
  );
  al_nand3 _06828_ (
    .a(_00367_),
    .b(_00556_),
    .c(_00363_),
    .y(_01894_)
  );
  al_ao21 _06829_ (
    .a(\DFF_289.Q ),
    .b(\DFF_910.Q ),
    .c(\DFF_575.Q ),
    .y(_01895_)
  );
  al_nand3ftt _06830_ (
    .a(_01353_),
    .b(_01895_),
    .c(_01894_),
    .y(_01896_)
  );
  al_ao21ftf _06831_ (
    .a(g35),
    .b(\DFF_910.Q ),
    .c(_01896_),
    .y(\DFF_575.D )
  );
  al_oai21ftf _06832_ (
    .a(\DFF_460.Q ),
    .b(\DFF_450.Q ),
    .c(\DFF_405.Q ),
    .y(_01897_)
  );
  al_nand3ftt _06833_ (
    .a(\DFF_147.Q ),
    .b(g35),
    .c(_01897_),
    .y(_01898_)
  );
  al_ao21ftf _06834_ (
    .a(g35),
    .b(\DFF_450.Q ),
    .c(_01898_),
    .y(\DFF_405.D )
  );
  al_and2ft _06835_ (
    .a(g35),
    .b(\DFF_1150.Q ),
    .y(_01899_)
  );
  al_nand2 _06836_ (
    .a(_00556_),
    .b(_00372_),
    .y(_01900_)
  );
  al_ao21 _06837_ (
    .a(\DFF_1150.Q ),
    .b(\DFF_1273.Q ),
    .c(\DFF_1068.Q ),
    .y(_01901_)
  );
  al_nor3fft _06838_ (
    .a(g35),
    .b(_01901_),
    .c(_00373_),
    .y(_01902_)
  );
  al_ao21 _06839_ (
    .a(_01902_),
    .b(_01900_),
    .c(_01899_),
    .y(\DFF_1068.D )
  );
  al_nand2ft _06840_ (
    .a(\DFF_343.Q ),
    .b(_01887_),
    .y(_01903_)
  );
  al_aoi21ttf _06841_ (
    .a(_01903_),
    .b(_01891_),
    .c(_01889_),
    .y(_01904_)
  );
  al_or3fft _06842_ (
    .a(\DFF_435.Q ),
    .b(_01904_),
    .c(_01890_),
    .y(_01905_)
  );
  al_oai21ftf _06843_ (
    .a(\DFF_435.Q ),
    .b(_01890_),
    .c(_01904_),
    .y(_01906_)
  );
  al_ao21 _06844_ (
    .a(_01905_),
    .b(_01906_),
    .c(_00066_),
    .y(_01907_)
  );
  al_aoi21ftf _06845_ (
    .a(\DFF_18.Q ),
    .b(_00066_),
    .c(_01907_),
    .y(\DFF_435.D )
  );
  al_oai21ftf _06846_ (
    .a(\DFF_147.Q ),
    .b(\DFF_299.Q ),
    .c(\DFF_478.Q ),
    .y(_01908_)
  );
  al_nand3ftt _06847_ (
    .a(\DFF_460.Q ),
    .b(g35),
    .c(_01908_),
    .y(_01909_)
  );
  al_ao21ftf _06848_ (
    .a(g35),
    .b(\DFF_299.Q ),
    .c(_01909_),
    .y(\DFF_478.D )
  );
  al_and3 _06849_ (
    .a(\DFF_1290.Q ),
    .b(_01001_),
    .c(_01211_),
    .y(_01910_)
  );
  al_or2 _06850_ (
    .a(_00291_),
    .b(_01910_),
    .y(_01911_)
  );
  al_nand2 _06851_ (
    .a(_00291_),
    .b(_01910_),
    .y(_01912_)
  );
  al_nand3 _06852_ (
    .a(g35),
    .b(_01912_),
    .c(_01911_),
    .y(_01913_)
  );
  al_aoi21ftf _06853_ (
    .a(\DFF_1290.Q ),
    .b(_00066_),
    .c(_01913_),
    .y(\DFF_296.D )
  );
  al_and3 _06854_ (
    .a(_00513_),
    .b(_00514_),
    .c(_00526_),
    .y(_01914_)
  );
  al_oa21ttf _06855_ (
    .a(\DFF_1034.Q ),
    .b(_01914_),
    .c(_00066_),
    .y(_01915_)
  );
  al_ao21ttf _06856_ (
    .a(\DFF_1034.Q ),
    .b(_01914_),
    .c(_01915_),
    .y(_01916_)
  );
  al_ao21ftf _06857_ (
    .a(g35),
    .b(\DFF_444.Q ),
    .c(_01916_),
    .y(\DFF_1034.D )
  );
  al_mux2l _06858_ (
    .a(\DFF_1172.Q ),
    .b(_01131_),
    .s(_01126_),
    .y(_01917_)
  );
  al_mux2h _06859_ (
    .a(\DFF_832.Q ),
    .b(_01917_),
    .s(g35),
    .y(\DFF_1172.D )
  );
  al_aoi21ttf _06860_ (
    .a(\DFF_67.Q ),
    .b(\DFF_60.Q ),
    .c(g35),
    .y(_01918_)
  );
  al_ao21ftf _06861_ (
    .a(\DFF_60.Q ),
    .b(\DFF_1407.Q ),
    .c(_01918_),
    .y(_01919_)
  );
  al_aoi21ftf _06862_ (
    .a(\DFF_717.Q ),
    .b(_00066_),
    .c(_01919_),
    .y(\DFF_1407.D )
  );
  al_nand2ft _06863_ (
    .a(\DFF_891.Q ),
    .b(\DFF_1324.Q ),
    .y(_01920_)
  );
  al_nand2ft _06864_ (
    .a(\DFF_1324.Q ),
    .b(\DFF_891.Q ),
    .y(_01921_)
  );
  al_ao21ttf _06865_ (
    .a(_01920_),
    .b(_01921_),
    .c(_01760_),
    .y(_01922_)
  );
  al_ao21ftf _06866_ (
    .a(g35),
    .b(\DFF_891.Q ),
    .c(_01922_),
    .y(\DFF_1324.D )
  );
  al_aoi21 _06867_ (
    .a(_00556_),
    .b(_00372_),
    .c(_00066_),
    .y(_01923_)
  );
  al_oai21 _06868_ (
    .a(_00508_),
    .b(_01104_),
    .c(_01923_),
    .y(_01924_)
  );
  al_ao21ftf _06869_ (
    .a(g35),
    .b(\DFF_410.Q ),
    .c(_01924_),
    .y(\DFF_584.D )
  );
  al_and3fft _06870_ (
    .a(\DFF_387.Q ),
    .b(\DFF_681.Q ),
    .c(\DFF_457.Q ),
    .y(_01925_)
  );
  al_ao21 _06871_ (
    .a(\DFF_4.Q ),
    .b(_01436_),
    .c(_01925_),
    .y(_01926_)
  );
  al_and3ftt _06872_ (
    .a(\DFF_297.Q ),
    .b(\DFF_681.Q ),
    .c(\DFF_1247.Q ),
    .y(_01927_)
  );
  al_ao21 _06873_ (
    .a(\DFF_65.Q ),
    .b(_01396_),
    .c(_01927_),
    .y(_01928_)
  );
  al_and3ftt _06874_ (
    .a(\DFF_297.Q ),
    .b(\DFF_625.Q ),
    .c(\DFF_387.Q ),
    .y(_01929_)
  );
  al_aoi21 _06875_ (
    .a(\DFF_469.Q ),
    .b(_00426_),
    .c(_01929_),
    .y(_01930_)
  );
  al_nand3fft _06876_ (
    .a(_01928_),
    .b(_01926_),
    .c(_01930_),
    .y(_01931_)
  );
  al_mux2l _06877_ (
    .a(_01931_),
    .b(\DFF_406.Q ),
    .s(_01394_),
    .y(_01932_)
  );
  al_mux2h _06878_ (
    .a(\DFF_681.Q ),
    .b(_01932_),
    .s(g35),
    .y(\DFF_406.D )
  );
  al_oai21ftf _06879_ (
    .a(g35),
    .b(_01544_),
    .c(\DFF_552.Q ),
    .y(_01933_)
  );
  al_aoi21ftf _06880_ (
    .a(\DFF_1037.Q ),
    .b(_01541_),
    .c(_01933_),
    .y(\DFF_1037.D )
  );
  al_inv _06881_ (
    .a(_00499_),
    .y(_01934_)
  );
  al_mux2h _06882_ (
    .a(\DFF_253.Q ),
    .b(_01934_),
    .s(_00361_),
    .y(_01935_)
  );
  al_mux2h _06883_ (
    .a(\DFF_414.Q ),
    .b(_01935_),
    .s(g35),
    .y(\DFF_253.D )
  );
  al_nand2 _06884_ (
    .a(\DFF_1084.Q ),
    .b(_00609_),
    .y(_01936_)
  );
  al_ao21ftf _06885_ (
    .a(\DFF_115.Q ),
    .b(_01936_),
    .c(_00607_),
    .y(_01937_)
  );
  al_ao21ftf _06886_ (
    .a(g35),
    .b(\DFF_1084.Q ),
    .c(_01937_),
    .y(\DFF_115.D )
  );
  al_nor2 _06887_ (
    .a(\DFF_976.Q ),
    .b(g35),
    .y(_01938_)
  );
  al_inv _06888_ (
    .a(\DFF_618.Q ),
    .y(_01939_)
  );
  al_nand2 _06889_ (
    .a(\DFF_834.Q ),
    .b(\DFF_176.Q ),
    .y(_01940_)
  );
  al_nand2 _06890_ (
    .a(\DFF_521.Q ),
    .b(\DFF_834.Q ),
    .y(_01941_)
  );
  al_mux2l _06891_ (
    .a(_01940_),
    .b(_01941_),
    .s(_00890_),
    .y(_01942_)
  );
  al_or3fft _06892_ (
    .a(\DFF_259.Q ),
    .b(_01939_),
    .c(_01942_),
    .y(_01943_)
  );
  al_nor2 _06893_ (
    .a(\DFF_834.Q ),
    .b(\DFF_176.Q ),
    .y(_01944_)
  );
  al_nor2 _06894_ (
    .a(\DFF_521.Q ),
    .b(\DFF_834.Q ),
    .y(_01945_)
  );
  al_mux2l _06895_ (
    .a(_01944_),
    .b(_01945_),
    .s(_00890_),
    .y(_01946_)
  );
  al_nand3 _06896_ (
    .a(\DFF_618.Q ),
    .b(\DFF_205.Q ),
    .c(_01946_),
    .y(_01947_)
  );
  al_and2 _06897_ (
    .a(_01947_),
    .b(_01943_),
    .y(_01948_)
  );
  al_mux2l _06898_ (
    .a(\DFF_259.Q ),
    .b(\DFF_205.Q ),
    .s(\DFF_976.Q ),
    .y(_01949_)
  );
  al_nand3ftt _06899_ (
    .a(_01949_),
    .b(\DFF_8.Q ),
    .c(_01948_),
    .y(_01950_)
  );
  al_aoi21ftf _06900_ (
    .a(\DFF_8.Q ),
    .b(_01949_),
    .c(g35),
    .y(_01951_)
  );
  al_aoi21 _06901_ (
    .a(_01951_),
    .b(_01950_),
    .c(_01938_),
    .y(\DFF_8.D )
  );
  al_and2ft _06902_ (
    .a(\DFF_68.Q ),
    .b(\DFF_598.Q ),
    .y(_01952_)
  );
  al_nand3 _06903_ (
    .a(_00499_),
    .b(_01409_),
    .c(_01952_),
    .y(_01953_)
  );
  al_ao21 _06904_ (
    .a(_01409_),
    .b(_01952_),
    .c(\DFF_1212.Q ),
    .y(_01954_)
  );
  al_nand3 _06905_ (
    .a(g35),
    .b(_01954_),
    .c(_01953_),
    .y(_01955_)
  );
  al_ao21ftf _06906_ (
    .a(g35),
    .b(\DFF_13.Q ),
    .c(_01955_),
    .y(\DFF_1212.D )
  );
  al_mux2l _06907_ (
    .a(\DFF_15.Q ),
    .b(\DFF_413.Q ),
    .s(g35),
    .y(\DFF_15.D )
  );
  al_aoi21ttf _06908_ (
    .a(_00454_),
    .b(_01662_),
    .c(\DFF_699.Q ),
    .y(_01956_)
  );
  al_and3 _06909_ (
    .a(\DFF_737.Q ),
    .b(\DFF_1320.Q ),
    .c(_00399_),
    .y(_01957_)
  );
  al_nand2 _06910_ (
    .a(_01957_),
    .b(_01956_),
    .y(_01958_)
  );
  al_or3fft _06911_ (
    .a(\DFF_213.Q ),
    .b(g35),
    .c(_01958_),
    .y(_01959_)
  );
  al_or2 _06912_ (
    .a(\DFF_361.Q ),
    .b(g35),
    .y(_01960_)
  );
  al_and2ft _06913_ (
    .a(\DFF_213.Q ),
    .b(g35),
    .y(_01961_)
  );
  al_ao21ttf _06914_ (
    .a(_01957_),
    .b(_01956_),
    .c(_01961_),
    .y(_01962_)
  );
  al_and3 _06915_ (
    .a(_01960_),
    .b(_01962_),
    .c(_01959_),
    .y(\DFF_213.D )
  );
  al_nand2 _06916_ (
    .a(\DFF_448.Q ),
    .b(g35),
    .y(_01963_)
  );
  al_and3 _06917_ (
    .a(\DFF_893.Q ),
    .b(\DFF_746.Q ),
    .c(\DFF_962.Q ),
    .y(_01964_)
  );
  al_and3 _06918_ (
    .a(\DFF_845.Q ),
    .b(\DFF_1364.Q ),
    .c(_01964_),
    .y(_01965_)
  );
  al_aoi21 _06919_ (
    .a(_00442_),
    .b(_01965_),
    .c(_01963_),
    .y(_01966_)
  );
  al_or2 _06920_ (
    .a(\DFF_1020.Q ),
    .b(g35),
    .y(_01967_)
  );
  al_and3 _06921_ (
    .a(\DFF_845.Q ),
    .b(_01964_),
    .c(_00549_),
    .y(_01968_)
  );
  al_aoi21ftf _06922_ (
    .a(_01963_),
    .b(_01968_),
    .c(_01967_),
    .y(_01969_)
  );
  al_aoi21ftf _06923_ (
    .a(\DFF_428.Q ),
    .b(_01966_),
    .c(_01969_),
    .y(\DFF_428.D )
  );
  al_nor2 _06924_ (
    .a(\DFF_189.Q ),
    .b(g35),
    .y(_01970_)
  );
  al_and3 _06925_ (
    .a(_00604_),
    .b(_00758_),
    .c(_00443_),
    .y(_01971_)
  );
  al_nand3ftt _06926_ (
    .a(\DFF_189.Q ),
    .b(\DFF_562.Q ),
    .c(\DFF_379.Q ),
    .y(_01972_)
  );
  al_oai21ftf _06927_ (
    .a(\DFF_562.Q ),
    .b(\DFF_189.Q ),
    .c(\DFF_379.Q ),
    .y(_01973_)
  );
  al_nand3 _06928_ (
    .a(_01972_),
    .b(_01973_),
    .c(_01971_),
    .y(_01974_)
  );
  al_oa21ftf _06929_ (
    .a(\DFF_581.Q ),
    .b(_01971_),
    .c(_00066_),
    .y(_01975_)
  );
  al_aoi21 _06930_ (
    .a(_01974_),
    .b(_01975_),
    .c(_01970_),
    .y(\DFF_581.D )
  );
  al_and2ft _06931_ (
    .a(\DFF_1304.Q ),
    .b(\DFF_407.Q ),
    .y(_01976_)
  );
  al_nand3 _06932_ (
    .a(_00499_),
    .b(_01408_),
    .c(_01976_),
    .y(_01977_)
  );
  al_ao21 _06933_ (
    .a(_01976_),
    .b(_01408_),
    .c(\DFF_983.Q ),
    .y(_01978_)
  );
  al_nand3 _06934_ (
    .a(g35),
    .b(_01978_),
    .c(_01977_),
    .y(_01979_)
  );
  al_ao21ftf _06935_ (
    .a(g35),
    .b(\DFF_602.Q ),
    .c(_01979_),
    .y(\DFF_983.D )
  );
  al_nand3 _06936_ (
    .a(_00498_),
    .b(_00499_),
    .c(_01702_),
    .y(_01980_)
  );
  al_ao21 _06937_ (
    .a(_00498_),
    .b(_01702_),
    .c(\DFF_44.Q ),
    .y(_01981_)
  );
  al_nand3 _06938_ (
    .a(g35),
    .b(_01981_),
    .c(_01980_),
    .y(_01982_)
  );
  al_ao21ftf _06939_ (
    .a(g35),
    .b(\DFF_71.Q ),
    .c(_01982_),
    .y(\DFF_44.D )
  );
  al_and2 _06940_ (
    .a(\DFF_1107.Q ),
    .b(_00466_),
    .y(_01983_)
  );
  al_aoi21 _06941_ (
    .a(_00744_),
    .b(_00388_),
    .c(_00066_),
    .y(_01984_)
  );
  al_and2ft _06942_ (
    .a(_01983_),
    .b(_01984_),
    .y(_01985_)
  );
  al_nand2 _06943_ (
    .a(\DFF_985.Q ),
    .b(_00466_),
    .y(_01986_)
  );
  al_or2 _06944_ (
    .a(\DFF_985.Q ),
    .b(_00466_),
    .y(_01987_)
  );
  al_nand3 _06945_ (
    .a(_01986_),
    .b(_01987_),
    .c(_01985_),
    .y(_01988_)
  );
  al_ao21ftf _06946_ (
    .a(g35),
    .b(\DFF_1029.Q ),
    .c(_01988_),
    .y(\DFF_985.D )
  );
  al_mux2l _06947_ (
    .a(\DFF_1403.Q ),
    .b(\DFF_311.Q ),
    .s(g35),
    .y(\DFF_1403.D )
  );
  al_and3 _06948_ (
    .a(\DFF_218.Q ),
    .b(\DFF_1107.Q ),
    .c(_00466_),
    .y(_01989_)
  );
  al_nand3 _06949_ (
    .a(\DFF_1199.Q ),
    .b(\DFF_914.Q ),
    .c(_01989_),
    .y(_01990_)
  );
  al_ao21 _06950_ (
    .a(\DFF_914.Q ),
    .b(_01989_),
    .c(\DFF_1199.Q ),
    .y(_01991_)
  );
  al_nand3 _06951_ (
    .a(_01990_),
    .b(_01991_),
    .c(_01984_),
    .y(_01992_)
  );
  al_ao21ftf _06952_ (
    .a(g35),
    .b(\DFF_914.Q ),
    .c(_01992_),
    .y(\DFF_1199.D )
  );
  al_inv _06953_ (
    .a(\DFF_308.Q ),
    .y(_01993_)
  );
  al_and3 _06954_ (
    .a(\DFF_426.Q ),
    .b(\DFF_394.Q ),
    .c(\DFF_396.Q ),
    .y(_01994_)
  );
  al_and3 _06955_ (
    .a(\DFF_1246.Q ),
    .b(\DFF_676.Q ),
    .c(_01994_),
    .y(_01995_)
  );
  al_and3 _06956_ (
    .a(\DFF_1015.Q ),
    .b(\DFF_260.Q ),
    .c(_01995_),
    .y(_01996_)
  );
  al_inv _06957_ (
    .a(\DFF_1015.Q ),
    .y(_01997_)
  );
  al_and3fft _06958_ (
    .a(\DFF_426.Q ),
    .b(\DFF_394.Q ),
    .c(\DFF_329.Q ),
    .y(_01998_)
  );
  al_nand3fft _06959_ (
    .a(\DFF_1246.Q ),
    .b(\DFF_676.Q ),
    .c(_01998_),
    .y(_01999_)
  );
  al_and3fft _06960_ (
    .a(\DFF_260.Q ),
    .b(_01999_),
    .c(_01997_),
    .y(_02000_)
  );
  al_oai21ttf _06961_ (
    .a(_02000_),
    .b(_01996_),
    .c(_01993_),
    .y(_02001_)
  );
  al_mux2l _06962_ (
    .a(\DFF_1015.Q ),
    .b(\DFF_308.Q ),
    .s(g84),
    .y(_02002_)
  );
  al_and2ft _06963_ (
    .a(\DFF_1271.Q ),
    .b(\DFF_260.Q ),
    .y(_02003_)
  );
  al_nand3 _06964_ (
    .a(\DFF_396.Q ),
    .b(_02002_),
    .c(_02003_),
    .y(_02004_)
  );
  al_and2 _06965_ (
    .a(\DFF_329.Q ),
    .b(\DFF_1271.Q ),
    .y(_02005_)
  );
  al_nand3fft _06966_ (
    .a(\DFF_260.Q ),
    .b(_02002_),
    .c(_02005_),
    .y(_02006_)
  );
  al_nand3 _06967_ (
    .a(\DFF_308.Q ),
    .b(_02004_),
    .c(_02006_),
    .y(_02007_)
  );
  al_nand3fft _06968_ (
    .a(_02000_),
    .b(_01996_),
    .c(_02007_),
    .y(_02008_)
  );
  al_nand3 _06969_ (
    .a(g35),
    .b(_02008_),
    .c(_02001_),
    .y(_02009_)
  );
  al_ao21ftf _06970_ (
    .a(g35),
    .b(\DFF_260.Q ),
    .c(_02009_),
    .y(\DFF_308.D )
  );
  al_and2ft _06971_ (
    .a(\DFF_27.Q ),
    .b(\DFF_120.Q ),
    .y(_02010_)
  );
  al_nor2 _06972_ (
    .a(\DFF_1408.Q ),
    .b(\DFF_199.Q ),
    .y(_02011_)
  );
  al_nand3 _06973_ (
    .a(_00499_),
    .b(_02010_),
    .c(_02011_),
    .y(_02012_)
  );
  al_ao21 _06974_ (
    .a(_02010_),
    .b(_02011_),
    .c(\DFF_227.Q ),
    .y(_02013_)
  );
  al_nand3 _06975_ (
    .a(g35),
    .b(_02013_),
    .c(_02012_),
    .y(_02014_)
  );
  al_ao21ftf _06976_ (
    .a(g35),
    .b(\DFF_707.Q ),
    .c(_02014_),
    .y(\DFF_227.D )
  );
  al_oa21ftt _06977_ (
    .a(\DFF_109.Q ),
    .b(\DFF_7.Q ),
    .c(\DFF_1235.Q ),
    .y(_02015_)
  );
  al_oai21ftf _06978_ (
    .a(_01187_),
    .b(_01186_),
    .c(_02015_),
    .y(_02016_)
  );
  al_nand3fft _06979_ (
    .a(_00066_),
    .b(_01188_),
    .c(_02016_),
    .y(_02017_)
  );
  al_ao21ftf _06980_ (
    .a(g35),
    .b(\DFF_863.Q ),
    .c(_02017_),
    .y(\DFF_1235.D )
  );
  al_inv _06981_ (
    .a(\DFF_794.Q ),
    .y(_02018_)
  );
  al_nand3fft _06982_ (
    .a(_02018_),
    .b(_01061_),
    .c(_01056_),
    .y(_02019_)
  );
  al_nand2 _06983_ (
    .a(\DFF_1226.Q ),
    .b(\DFF_33.Q ),
    .y(_02020_)
  );
  al_nor2 _06984_ (
    .a(\DFF_1226.Q ),
    .b(\DFF_33.Q ),
    .y(_02021_)
  );
  al_nand2ft _06985_ (
    .a(_02021_),
    .b(_02020_),
    .y(_02022_)
  );
  al_mux2l _06986_ (
    .a(\DFF_1418.Q ),
    .b(_02022_),
    .s(_02019_),
    .y(_02023_)
  );
  al_mux2h _06987_ (
    .a(\DFF_1226.Q ),
    .b(_02023_),
    .s(g35),
    .y(\DFF_1418.D )
  );
  al_nand3 _06988_ (
    .a(\DFF_870.Q ),
    .b(\DFF_1161.Q ),
    .c(_00477_),
    .y(_02024_)
  );
  al_ao21 _06989_ (
    .a(\DFF_1161.Q ),
    .b(_00477_),
    .c(\DFF_870.Q ),
    .y(_02025_)
  );
  al_nand2ft _06990_ (
    .a(\DFF_524.Q ),
    .b(\DFF_872.Q ),
    .y(_02026_)
  );
  al_aoi21 _06991_ (
    .a(\DFF_23.Q ),
    .b(_02026_),
    .c(_00066_),
    .y(_02027_)
  );
  al_nand3 _06992_ (
    .a(_02024_),
    .b(_02025_),
    .c(_02027_),
    .y(_02028_)
  );
  al_ao21ftf _06993_ (
    .a(g35),
    .b(\DFF_524.Q ),
    .c(_02028_),
    .y(\DFF_870.D )
  );
  al_mux2l _06994_ (
    .a(g64),
    .b(\DFF_194.Q ),
    .s(g35),
    .y(\DFF_515.D )
  );
  al_and2 _06995_ (
    .a(\DFF_1408.Q ),
    .b(\DFF_199.Q ),
    .y(_02029_)
  );
  al_or3 _06996_ (
    .a(\DFF_245.Q ),
    .b(\DFF_120.Q ),
    .c(\DFF_27.Q ),
    .y(_02030_)
  );
  al_nand3ftt _06997_ (
    .a(_02030_),
    .b(_02029_),
    .c(_00499_),
    .y(_02031_)
  );
  al_ao21ftt _06998_ (
    .a(_02030_),
    .b(_02029_),
    .c(\DFF_309.Q ),
    .y(_02032_)
  );
  al_nand3 _06999_ (
    .a(g35),
    .b(_02031_),
    .c(_02032_),
    .y(_02033_)
  );
  al_ao21ftf _07000_ (
    .a(g35),
    .b(\DFF_738.Q ),
    .c(_02033_),
    .y(\DFF_309.D )
  );
  al_ao21 _07001_ (
    .a(_00465_),
    .b(_01865_),
    .c(_00066_),
    .y(_02034_)
  );
  al_oa21ftf _07002_ (
    .a(\DFF_1424.Q ),
    .b(_01864_),
    .c(_00066_),
    .y(_02035_)
  );
  al_and2 _07003_ (
    .a(\DFF_1199.Q ),
    .b(\DFF_892.Q ),
    .y(_02036_)
  );
  al_aoi21 _07004_ (
    .a(_00464_),
    .b(_02036_),
    .c(\DFF_313.Q ),
    .y(_02037_)
  );
  al_ao21ftf _07005_ (
    .a(_02037_),
    .b(_01864_),
    .c(_02035_),
    .y(_02038_)
  );
  al_aoi21ftf _07006_ (
    .a(\DFF_782.Q ),
    .b(_02034_),
    .c(_02038_),
    .y(\DFF_313.D )
  );
  al_inv _07007_ (
    .a(\DFF_1236.Q ),
    .y(_02039_)
  );
  al_aoi21ttf _07008_ (
    .a(_00577_),
    .b(_00438_),
    .c(_01363_),
    .y(_02040_)
  );
  al_oa21ftf _07009_ (
    .a(_01362_),
    .b(_01363_),
    .c(_00066_),
    .y(_02041_)
  );
  al_ao21ttf _07010_ (
    .a(_02039_),
    .b(_02040_),
    .c(_02041_),
    .y(_02042_)
  );
  al_ao21ftf _07011_ (
    .a(g35),
    .b(\DFF_1093.Q ),
    .c(_02042_),
    .y(\DFF_1295.D )
  );
  al_or2 _07012_ (
    .a(g35),
    .b(\DFF_239.Q ),
    .y(_02043_)
  );
  al_aoi21ftf _07013_ (
    .a(\DFF_541.Q ),
    .b(_01579_),
    .c(_02043_),
    .y(_02044_)
  );
  al_oa21 _07014_ (
    .a(\DFF_324.Q ),
    .b(_01174_),
    .c(_02044_),
    .y(\DFF_324.D )
  );
  al_and3 _07015_ (
    .a(_01534_),
    .b(_01535_),
    .c(_00974_),
    .y(_02045_)
  );
  al_nand2 _07016_ (
    .a(\DFF_1395.Q ),
    .b(\DFF_1268.Q ),
    .y(_02046_)
  );
  al_nor2 _07017_ (
    .a(\DFF_1395.Q ),
    .b(\DFF_1268.Q ),
    .y(_02047_)
  );
  al_nand2ft _07018_ (
    .a(_02047_),
    .b(_02046_),
    .y(_02048_)
  );
  al_mux2l _07019_ (
    .a(_02048_),
    .b(\DFF_488.Q ),
    .s(_02045_),
    .y(_02049_)
  );
  al_mux2h _07020_ (
    .a(\DFF_1268.Q ),
    .b(_02049_),
    .s(g35),
    .y(\DFF_488.D )
  );
  al_and3fft _07021_ (
    .a(\DFF_798.Q ),
    .b(\DFF_269.Q ),
    .c(g35),
    .y(\DFF_269.D )
  );
  al_nor2 _07022_ (
    .a(\DFF_851.Q ),
    .b(g35),
    .y(_02050_)
  );
  al_mux2l _07023_ (
    .a(\DFF_838.Q ),
    .b(\DFF_1048.Q ),
    .s(\DFF_851.Q ),
    .y(_02051_)
  );
  al_nand3ftt _07024_ (
    .a(_02051_),
    .b(\DFF_122.Q ),
    .c(_00899_),
    .y(_02052_)
  );
  al_aoi21ftf _07025_ (
    .a(\DFF_122.Q ),
    .b(_02051_),
    .c(g35),
    .y(_02053_)
  );
  al_aoi21 _07026_ (
    .a(_02053_),
    .b(_02052_),
    .c(_02050_),
    .y(\DFF_122.D )
  );
  al_nand2ft _07027_ (
    .a(\DFF_368.Q ),
    .b(_00847_),
    .y(_02054_)
  );
  al_nand3 _07028_ (
    .a(g35),
    .b(_02054_),
    .c(_00848_),
    .y(_02055_)
  );
  al_ao21ftf _07029_ (
    .a(g35),
    .b(\DFF_70.Q ),
    .c(_02055_),
    .y(\DFF_368.D )
  );
  al_ao21ttf _07030_ (
    .a(_00836_),
    .b(_00837_),
    .c(_00844_),
    .y(_02056_)
  );
  al_ao21 _07031_ (
    .a(g35),
    .b(_02056_),
    .c(_00835_),
    .y(_02057_)
  );
  al_nand2 _07032_ (
    .a(\DFF_368.Q ),
    .b(\DFF_421.Q ),
    .y(_02058_)
  );
  al_ao21ttf _07033_ (
    .a(_02058_),
    .b(_00838_),
    .c(_00844_),
    .y(_02059_)
  );
  al_and2 _07034_ (
    .a(\DFF_979.Q ),
    .b(g35),
    .y(_02060_)
  );
  al_ao21ttf _07035_ (
    .a(_02060_),
    .b(_02059_),
    .c(_02057_),
    .y(\DFF_979.D )
  );
  al_and2ft _07036_ (
    .a(g35),
    .b(\DFF_1188.Q ),
    .y(_02061_)
  );
  al_ao21 _07037_ (
    .a(_01663_),
    .b(_01751_),
    .c(\DFF_139.Q ),
    .y(_02062_)
  );
  al_aoi21 _07038_ (
    .a(\DFF_139.Q ),
    .b(_01663_),
    .c(_00066_),
    .y(_02063_)
  );
  al_ao21 _07039_ (
    .a(_02063_),
    .b(_02062_),
    .c(_02061_),
    .y(\DFF_139.D )
  );
  al_aoi21ttf _07040_ (
    .a(_00468_),
    .b(_00584_),
    .c(\DFF_130.Q ),
    .y(_02064_)
  );
  al_nand3 _07041_ (
    .a(\DFF_670.Q ),
    .b(\DFF_1359.Q ),
    .c(_00390_),
    .y(_02065_)
  );
  al_and2ft _07042_ (
    .a(\DFF_1347.Q ),
    .b(\DFF_443.Q ),
    .y(_02066_)
  );
  al_nand3 _07043_ (
    .a(\DFF_370.Q ),
    .b(\DFF_76.Q ),
    .c(_02066_),
    .y(_02067_)
  );
  al_and3 _07044_ (
    .a(\DFF_538.Q ),
    .b(_02067_),
    .c(_02065_),
    .y(_02068_)
  );
  al_or2 _07045_ (
    .a(\DFF_1347.Q ),
    .b(\DFF_443.Q ),
    .y(_02069_)
  );
  al_nand2 _07046_ (
    .a(\DFF_1378.Q ),
    .b(\DFF_1155.Q ),
    .y(_02070_)
  );
  al_nand2 _07047_ (
    .a(\DFF_1263.Q ),
    .b(\DFF_1303.Q ),
    .y(_02071_)
  );
  al_ao21 _07048_ (
    .a(_02070_),
    .b(_02071_),
    .c(_02069_),
    .y(_02072_)
  );
  al_nand2ft _07049_ (
    .a(\DFF_443.Q ),
    .b(\DFF_1347.Q ),
    .y(_02073_)
  );
  al_nand2 _07050_ (
    .a(\DFF_1218.Q ),
    .b(\DFF_856.Q ),
    .y(_02074_)
  );
  al_nand2 _07051_ (
    .a(\DFF_819.Q ),
    .b(\DFF_1386.Q ),
    .y(_02075_)
  );
  al_ao21 _07052_ (
    .a(_02074_),
    .b(_02075_),
    .c(_02073_),
    .y(_02076_)
  );
  al_nand3 _07053_ (
    .a(_02072_),
    .b(_02076_),
    .c(_02068_),
    .y(_02077_)
  );
  al_nand2 _07054_ (
    .a(\DFF_1351.Q ),
    .b(\DFF_1303.Q ),
    .y(_02078_)
  );
  al_nand2 _07055_ (
    .a(\DFF_1197.Q ),
    .b(\DFF_1155.Q ),
    .y(_02079_)
  );
  al_ao21ttf _07056_ (
    .a(_02078_),
    .b(_02079_),
    .c(_02066_),
    .y(_02080_)
  );
  al_or3fft _07057_ (
    .a(\DFF_134.Q ),
    .b(\DFF_76.Q ),
    .c(_02069_),
    .y(_02081_)
  );
  al_and3 _07058_ (
    .a(_00736_),
    .b(_02081_),
    .c(_02080_),
    .y(_02082_)
  );
  al_nand2 _07059_ (
    .a(\DFF_1354.Q ),
    .b(\DFF_645.Q ),
    .y(_02083_)
  );
  al_nand2 _07060_ (
    .a(\DFF_1280.Q ),
    .b(\DFF_1359.Q ),
    .y(_02084_)
  );
  al_ao21 _07061_ (
    .a(_02083_),
    .b(_02084_),
    .c(_02073_),
    .y(_02085_)
  );
  al_nand2 _07062_ (
    .a(\DFF_819.Q ),
    .b(\DFF_1208.Q ),
    .y(_02086_)
  );
  al_aoi21ttf _07063_ (
    .a(\DFF_1401.Q ),
    .b(\DFF_856.Q ),
    .c(_02086_),
    .y(_02087_)
  );
  al_oai21ftt _07064_ (
    .a(_00390_),
    .b(_02087_),
    .c(_02085_),
    .y(_02088_)
  );
  al_ao21ftf _07065_ (
    .a(_02088_),
    .b(_02082_),
    .c(_02077_),
    .y(_02089_)
  );
  al_and3 _07066_ (
    .a(\DFF_538.Q ),
    .b(\DFF_1354.Q ),
    .c(_00390_),
    .y(_02090_)
  );
  al_and3 _07067_ (
    .a(\DFF_1038.Q ),
    .b(\DFF_225.Q ),
    .c(_00390_),
    .y(_02091_)
  );
  al_or3fft _07068_ (
    .a(\DFF_1293.Q ),
    .b(\DFF_1410.Q ),
    .c(_02069_),
    .y(_02092_)
  );
  al_nor2 _07069_ (
    .a(\DFF_819.Q ),
    .b(\DFF_538.Q ),
    .y(_02093_)
  );
  al_nand2 _07070_ (
    .a(\DFF_819.Q ),
    .b(\DFF_538.Q ),
    .y(_02094_)
  );
  al_nand2ft _07071_ (
    .a(_02093_),
    .b(_02094_),
    .y(_02095_)
  );
  al_and3 _07072_ (
    .a(\DFF_529.Q ),
    .b(\DFF_1166.Q ),
    .c(_02066_),
    .y(_02096_)
  );
  al_and3ftt _07073_ (
    .a(_02096_),
    .b(_02092_),
    .c(_02095_),
    .y(_02097_)
  );
  al_nand3 _07074_ (
    .a(\DFF_1293.Q ),
    .b(\DFF_1210.Q ),
    .c(_02066_),
    .y(_02098_)
  );
  al_and3ftt _07075_ (
    .a(_02093_),
    .b(_02094_),
    .c(_02098_),
    .y(_02099_)
  );
  al_or3fft _07076_ (
    .a(\DFF_1038.Q ),
    .b(\DFF_9.Q ),
    .c(_02073_),
    .y(_02100_)
  );
  al_or3fft _07077_ (
    .a(\DFF_529.Q ),
    .b(\DFF_640.Q ),
    .c(_02069_),
    .y(_02101_)
  );
  al_nand3 _07078_ (
    .a(_02100_),
    .b(_02101_),
    .c(_02099_),
    .y(_02102_)
  );
  al_ao21ftf _07079_ (
    .a(_02091_),
    .b(_02097_),
    .c(_02102_),
    .y(_02103_)
  );
  al_aoi21ttf _07080_ (
    .a(\DFF_729.Q ),
    .b(_02090_),
    .c(_02103_),
    .y(_02104_)
  );
  al_ao21ttf _07081_ (
    .a(_02089_),
    .b(_02104_),
    .c(_02064_),
    .y(_02105_)
  );
  al_nand2 _07082_ (
    .a(_02090_),
    .b(_02064_),
    .y(_02106_)
  );
  al_nand3 _07083_ (
    .a(\DFF_1372.Q ),
    .b(_02106_),
    .c(_02105_),
    .y(_02107_)
  );
  al_ao21 _07084_ (
    .a(\DFF_1372.Q ),
    .b(_02106_),
    .c(_02105_),
    .y(_02108_)
  );
  al_nand3 _07085_ (
    .a(g35),
    .b(_02107_),
    .c(_02108_),
    .y(_02109_)
  );
  al_aoi21ftf _07086_ (
    .a(\DFF_124.Q ),
    .b(_00066_),
    .c(_02109_),
    .y(\DFF_1372.D )
  );
  al_nand3ftt _07087_ (
    .a(_01768_),
    .b(_00499_),
    .c(_01354_),
    .y(_02110_)
  );
  al_ao21ftt _07088_ (
    .a(_01768_),
    .b(_01354_),
    .c(\DFF_494.Q ),
    .y(_02111_)
  );
  al_nand3 _07089_ (
    .a(g35),
    .b(_02110_),
    .c(_02111_),
    .y(_02112_)
  );
  al_ao21ftf _07090_ (
    .a(g35),
    .b(\DFF_337.Q ),
    .c(_02112_),
    .y(\DFF_494.D )
  );
  al_and2 _07091_ (
    .a(\DFF_271.Q ),
    .b(\DFF_522.Q ),
    .y(_02113_)
  );
  al_and2ft _07092_ (
    .a(\DFF_803.Q ),
    .b(\DFF_35.Q ),
    .y(_02114_)
  );
  al_nand3 _07093_ (
    .a(_00499_),
    .b(_02113_),
    .c(_02114_),
    .y(_02115_)
  );
  al_ao21 _07094_ (
    .a(_02114_),
    .b(_02113_),
    .c(\DFF_640.Q ),
    .y(_02116_)
  );
  al_nand3 _07095_ (
    .a(g35),
    .b(_02116_),
    .c(_02115_),
    .y(_02117_)
  );
  al_ao21ftf _07096_ (
    .a(g35),
    .b(\DFF_1208.Q ),
    .c(_02117_),
    .y(\DFF_640.D )
  );
  al_nand3ftt _07097_ (
    .a(\DFF_598.Q ),
    .b(\DFF_68.Q ),
    .c(\DFF_1098.Q ),
    .y(_02118_)
  );
  al_aoi21ftf _07098_ (
    .a(\DFF_1040.Q ),
    .b(_02118_),
    .c(g35),
    .y(_02119_)
  );
  al_ao21ftf _07099_ (
    .a(_02118_),
    .b(_00499_),
    .c(_02119_),
    .y(_02120_)
  );
  al_ao21ftf _07100_ (
    .a(g35),
    .b(\DFF_1406.Q ),
    .c(_02120_),
    .y(\DFF_1040.D )
  );
  al_aoi21 _07101_ (
    .a(\DFF_1005.Q ),
    .b(_01555_),
    .c(_00066_),
    .y(_02121_)
  );
  al_nand2ft _07102_ (
    .a(g35),
    .b(\DFF_1005.Q ),
    .y(_02122_)
  );
  al_ao21ftf _07103_ (
    .a(\DFF_1188.Q ),
    .b(_02121_),
    .c(_02122_),
    .y(\DFF_251.D )
  );
  al_nor2 _07104_ (
    .a(\DFF_1147.Q ),
    .b(g35),
    .y(_02123_)
  );
  al_mux2l _07105_ (
    .a(_01683_),
    .b(_01680_),
    .s(_01678_),
    .y(_02124_)
  );
  al_or3fft _07106_ (
    .a(\DFF_1257.Q ),
    .b(_01042_),
    .c(_02124_),
    .y(_02125_)
  );
  al_aoi21ftf _07107_ (
    .a(\DFF_1257.Q ),
    .b(_02124_),
    .c(g35),
    .y(_02126_)
  );
  al_aoi21 _07108_ (
    .a(_02125_),
    .b(_02126_),
    .c(_02123_),
    .y(\DFF_1257.D )
  );
  al_and2 _07109_ (
    .a(g35),
    .b(\DFF_1059.Q ),
    .y(\DFF_585.D )
  );
  al_nor2 _07110_ (
    .a(\DFF_951.Q ),
    .b(g35),
    .y(_02127_)
  );
  al_nand3ftt _07111_ (
    .a(\DFF_451.Q ),
    .b(\DFF_951.Q ),
    .c(_01968_),
    .y(_02128_)
  );
  al_nand2 _07112_ (
    .a(\DFF_951.Q ),
    .b(_01968_),
    .y(_02129_)
  );
  al_aoi21 _07113_ (
    .a(\DFF_451.Q ),
    .b(_02129_),
    .c(_01963_),
    .y(_02130_)
  );
  al_aoi21 _07114_ (
    .a(_02128_),
    .b(_02130_),
    .c(_02127_),
    .y(\DFF_451.D )
  );
  al_inv _07115_ (
    .a(\DFF_521.Q ),
    .y(_02131_)
  );
  al_and3fft _07116_ (
    .a(\DFF_8.Q ),
    .b(\DFF_976.Q ),
    .c(\DFF_205.Q ),
    .y(_02132_)
  );
  al_nand3fft _07117_ (
    .a(\DFF_725.Q ),
    .b(\DFF_592.Q ),
    .c(_02132_),
    .y(_02133_)
  );
  al_and3 _07118_ (
    .a(\DFF_259.Q ),
    .b(\DFF_8.Q ),
    .c(\DFF_976.Q ),
    .y(_02134_)
  );
  al_nand3 _07119_ (
    .a(\DFF_725.Q ),
    .b(\DFF_592.Q ),
    .c(_02134_),
    .y(_02135_)
  );
  al_mux2l _07120_ (
    .a(_02133_),
    .b(_02135_),
    .s(_02131_),
    .y(_02136_)
  );
  al_nand3 _07121_ (
    .a(\DFF_834.Q ),
    .b(_02136_),
    .c(_01948_),
    .y(_02137_)
  );
  al_oai21 _07122_ (
    .a(\DFF_834.Q ),
    .b(_02136_),
    .c(_02137_),
    .y(_02138_)
  );
  al_mux2h _07123_ (
    .a(\DFF_521.Q ),
    .b(_02138_),
    .s(g35),
    .y(\DFF_834.D )
  );
  al_or3fft _07124_ (
    .a(_01449_),
    .b(_01455_),
    .c(_01453_),
    .y(_02139_)
  );
  al_ao21 _07125_ (
    .a(_01449_),
    .b(_01452_),
    .c(\DFF_1388.Q ),
    .y(_02140_)
  );
  al_nand3 _07126_ (
    .a(g35),
    .b(_02140_),
    .c(_02139_),
    .y(_02141_)
  );
  al_aoi21ftf _07127_ (
    .a(\DFF_586.Q ),
    .b(_00066_),
    .c(_02141_),
    .y(\DFF_1388.D )
  );
  al_mux2l _07128_ (
    .a(\DFF_1035.Q ),
    .b(\DFF_706.Q ),
    .s(g35),
    .y(\DFF_1035.D )
  );
  al_aoi21 _07129_ (
    .a(\DFF_965.Q ),
    .b(_00748_),
    .c(_01822_),
    .y(_02142_)
  );
  al_ao21 _07130_ (
    .a(g35),
    .b(_01825_),
    .c(_02142_),
    .y(\DFF_965.D )
  );
  al_nand3 _07131_ (
    .a(_00499_),
    .b(_01952_),
    .c(_01976_),
    .y(_02143_)
  );
  al_ao21 _07132_ (
    .a(_01952_),
    .b(_01976_),
    .c(\DFF_13.Q ),
    .y(_02144_)
  );
  al_nand3 _07133_ (
    .a(g35),
    .b(_02144_),
    .c(_02143_),
    .y(_02145_)
  );
  al_ao21ftf _07134_ (
    .a(g35),
    .b(\DFF_390.Q ),
    .c(_02145_),
    .y(\DFF_13.D )
  );
  al_nand3 _07135_ (
    .a(g35),
    .b(_00744_),
    .c(_00388_),
    .y(_02146_)
  );
  al_ao21 _07136_ (
    .a(\DFF_1326.Q ),
    .b(g35),
    .c(\DFF_99.Q ),
    .y(_02147_)
  );
  al_nand3 _07137_ (
    .a(\DFF_99.Q ),
    .b(\DFF_1326.Q ),
    .c(g35),
    .y(_02148_)
  );
  al_and3 _07138_ (
    .a(_02147_),
    .b(_02148_),
    .c(_02146_),
    .y(\DFF_1326.D )
  );
  al_nor2 _07139_ (
    .a(\DFF_153.Q ),
    .b(\DFF_1009.Q ),
    .y(_02149_)
  );
  al_nand3fft _07140_ (
    .a(\DFF_1063.Q ),
    .b(\DFF_472.Q ),
    .c(_02149_),
    .y(_02150_)
  );
  al_or3 _07141_ (
    .a(\DFF_342.Q ),
    .b(\DFF_1093.Q ),
    .c(_02150_),
    .y(_02151_)
  );
  al_or3 _07142_ (
    .a(\DFF_567.Q ),
    .b(\DFF_1089.Q ),
    .c(_02151_),
    .y(_02152_)
  );
  al_nor2 _07143_ (
    .a(\DFF_462.Q ),
    .b(\DFF_1028.Q ),
    .y(_02153_)
  );
  al_or2 _07144_ (
    .a(\DFF_1254.Q ),
    .b(\DFF_1337.Q ),
    .y(_02154_)
  );
  al_nor2 _07145_ (
    .a(\DFF_594.Q ),
    .b(\DFF_943.Q ),
    .y(_02155_)
  );
  al_nand3fft _07146_ (
    .a(\DFF_581.Q ),
    .b(\DFF_658.Q ),
    .c(_02155_),
    .y(_02156_)
  );
  al_and3fft _07147_ (
    .a(_02154_),
    .b(_02156_),
    .c(_02153_),
    .y(_02157_)
  );
  al_and3ftt _07148_ (
    .a(\DFF_733.Q ),
    .b(g91),
    .c(g35),
    .y(_02158_)
  );
  al_or3fft _07149_ (
    .a(_02157_),
    .b(_02158_),
    .c(_02152_),
    .y(_02159_)
  );
  al_aoi21ftf _07150_ (
    .a(\DFF_95.Q ),
    .b(_00066_),
    .c(_02159_),
    .y(\DFF_733.D )
  );
  al_and2 _07151_ (
    .a(\DFF_160.Q ),
    .b(_02146_),
    .y(\DFF_99.D )
  );
  al_or3ftt _07152_ (
    .a(\DFF_1273.Q ),
    .b(\DFF_1150.Q ),
    .c(\DFF_1068.Q ),
    .y(_02160_)
  );
  al_aoi21ftf _07153_ (
    .a(\DFF_967.Q ),
    .b(_02160_),
    .c(g35),
    .y(_02161_)
  );
  al_ao21ftf _07154_ (
    .a(_02160_),
    .b(_00499_),
    .c(_02161_),
    .y(_02162_)
  );
  al_ao21ftf _07155_ (
    .a(g35),
    .b(\DFF_617.Q ),
    .c(_02162_),
    .y(\DFF_967.D )
  );
  al_nor2 _07156_ (
    .a(\DFF_426.Q ),
    .b(g35),
    .y(_02163_)
  );
  al_and2 _07157_ (
    .a(_02004_),
    .b(_02006_),
    .y(_02164_)
  );
  al_mux2l _07158_ (
    .a(\DFF_396.Q ),
    .b(\DFF_329.Q ),
    .s(\DFF_426.Q ),
    .y(_02165_)
  );
  al_nand3ftt _07159_ (
    .a(_02165_),
    .b(\DFF_394.Q ),
    .c(_02164_),
    .y(_02166_)
  );
  al_aoi21ftf _07160_ (
    .a(\DFF_394.Q ),
    .b(_02165_),
    .c(g35),
    .y(_02167_)
  );
  al_aoi21 _07161_ (
    .a(_02167_),
    .b(_02166_),
    .c(_02163_),
    .y(\DFF_394.D )
  );
  al_mux2l _07162_ (
    .a(\DFF_231.Q ),
    .b(\DFF_766.Q ),
    .s(g35),
    .y(\DFF_231.D )
  );
  al_or2ft _07163_ (
    .a(\DFF_287.Q ),
    .b(_00376_),
    .y(_02168_)
  );
  al_inv _07164_ (
    .a(\DFF_275.Q ),
    .y(_02169_)
  );
  al_or2ft _07165_ (
    .a(g35),
    .b(_00376_),
    .y(_02170_)
  );
  al_and2ft _07166_ (
    .a(\DFF_1004.Q ),
    .b(g35),
    .y(_02171_)
  );
  al_ao21ftf _07167_ (
    .a(_02169_),
    .b(_02171_),
    .c(_02170_),
    .y(_02172_)
  );
  al_and3ftt _07168_ (
    .a(_02171_),
    .b(_02169_),
    .c(_02170_),
    .y(_02173_)
  );
  al_aoi21 _07169_ (
    .a(_02168_),
    .b(_02172_),
    .c(_02173_),
    .y(\DFF_287.D )
  );
  al_inv _07170_ (
    .a(\DFF_496.Q ),
    .y(_02174_)
  );
  al_and2ft _07171_ (
    .a(\DFF_771.Q ),
    .b(\DFF_382.Q ),
    .y(_02175_)
  );
  al_oa21ttf _07172_ (
    .a(_00926_),
    .b(_02175_),
    .c(_02174_),
    .y(_02176_)
  );
  al_or3 _07173_ (
    .a(\DFF_496.Q ),
    .b(_00926_),
    .c(_02175_),
    .y(_02177_)
  );
  al_nor2ft _07174_ (
    .a(_02177_),
    .b(_02176_),
    .y(_02178_)
  );
  al_nand2ft _07175_ (
    .a(_00931_),
    .b(_00927_),
    .y(_02179_)
  );
  al_oai21ttf _07176_ (
    .a(_00925_),
    .b(_00932_),
    .c(_02179_),
    .y(_02180_)
  );
  al_nand3fft _07177_ (
    .a(_00925_),
    .b(_00932_),
    .c(_02179_),
    .y(_02181_)
  );
  al_aoi21 _07178_ (
    .a(_02181_),
    .b(_02180_),
    .c(_02178_),
    .y(_02182_)
  );
  al_nand3 _07179_ (
    .a(_02181_),
    .b(_02180_),
    .c(_02178_),
    .y(_02183_)
  );
  al_nand2ft _07180_ (
    .a(_02182_),
    .b(_02183_),
    .y(_02184_)
  );
  al_nand3ftt _07181_ (
    .a(_00481_),
    .b(\DFF_988.Q ),
    .c(_02184_),
    .y(_02185_)
  );
  al_ao21ftt _07182_ (
    .a(_00481_),
    .b(\DFF_988.Q ),
    .c(_02184_),
    .y(_02186_)
  );
  al_and3 _07183_ (
    .a(g35),
    .b(_02185_),
    .c(_02186_),
    .y(\DFF_988.D )
  );
  al_aoi21 _07184_ (
    .a(\DFF_33.Q ),
    .b(_00722_),
    .c(_00066_),
    .y(_02187_)
  );
  al_oai21 _07185_ (
    .a(\DFF_33.Q ),
    .b(_00722_),
    .c(_02187_),
    .y(_02188_)
  );
  al_aoi21ftf _07186_ (
    .a(\DFF_1277.Q ),
    .b(_00066_),
    .c(_02188_),
    .y(\DFF_33.D )
  );
  al_mux2l _07187_ (
    .a(\DFF_1004.Q ),
    .b(\DFF_275.Q ),
    .s(_02170_),
    .y(\DFF_275.D )
  );
  al_oa21 _07188_ (
    .a(\DFF_116.Q ),
    .b(\DFF_25.Q ),
    .c(g35),
    .y(\DFF_25.D )
  );
  al_oa21 _07189_ (
    .a(\DFF_294.Q ),
    .b(\DFF_532.Q ),
    .c(g35),
    .y(_02189_)
  );
  al_mux2l _07190_ (
    .a(_00066_),
    .b(_02189_),
    .s(\DFF_240.Q ),
    .y(\DFF_294.D )
  );
  al_oa21ftt _07191_ (
    .a(g35),
    .b(\DFF_1124.Q ),
    .c(\DFF_1116.Q ),
    .y(\DFF_288.D )
  );
  al_or2 _07192_ (
    .a(_00066_),
    .b(_02045_),
    .y(_02190_)
  );
  al_mux2l _07193_ (
    .a(\DFF_1395.Q ),
    .b(\DFF_1268.Q ),
    .s(_02190_),
    .y(\DFF_1268.D )
  );
  al_aoi21 _07194_ (
    .a(\DFF_910.Q ),
    .b(g35),
    .c(\DFF_289.Q ),
    .y(_02191_)
  );
  al_inv _07195_ (
    .a(\DFF_289.Q ),
    .y(_02192_)
  );
  al_ao21ftf _07196_ (
    .a(_02192_),
    .b(\DFF_910.Q ),
    .c(_01894_),
    .y(_02193_)
  );
  al_aoi21 _07197_ (
    .a(g35),
    .b(_02193_),
    .c(_02191_),
    .y(\DFF_910.D )
  );
  al_mux2l _07198_ (
    .a(\DFF_1340.Q ),
    .b(\DFF_1417.Q ),
    .s(g35),
    .y(\DFF_1340.D )
  );
  al_aoi21 _07199_ (
    .a(\DFF_203.Q ),
    .b(g35),
    .c(\DFF_509.Q ),
    .y(_02194_)
  );
  al_nand3 _07200_ (
    .a(\DFF_203.Q ),
    .b(g35),
    .c(\DFF_509.Q ),
    .y(_02195_)
  );
  al_and2ft _07201_ (
    .a(_02194_),
    .b(_02195_),
    .y(\DFF_349.D )
  );
  al_or3 _07202_ (
    .a(\DFF_511.Q ),
    .b(\DFF_1207.Q ),
    .c(\DFF_675.Q ),
    .y(_02196_)
  );
  al_nand3 _07203_ (
    .a(\DFF_339.Q ),
    .b(\DFF_261.Q ),
    .c(_02196_),
    .y(_02197_)
  );
  al_and2ft _07204_ (
    .a(\DFF_698.Q ),
    .b(g35),
    .y(_02198_)
  );
  al_aoi21ftf _07205_ (
    .a(\DFF_1133.Q ),
    .b(_02197_),
    .c(_02198_),
    .y(_02199_)
  );
  al_ao21ftf _07206_ (
    .a(_02197_),
    .b(\DFF_1133.Q ),
    .c(_02199_),
    .y(_02200_)
  );
  al_ao21ftf _07207_ (
    .a(g35),
    .b(\DFF_261.Q ),
    .c(_02200_),
    .y(\DFF_1133.D )
  );
  al_nand3 _07208_ (
    .a(_01535_),
    .b(\DFF_265.Q ),
    .c(_00974_),
    .y(_02201_)
  );
  al_aoi21ftf _07209_ (
    .a(\DFF_887.Q ),
    .b(_02201_),
    .c(g35),
    .y(_02202_)
  );
  al_oai21 _07210_ (
    .a(_00977_),
    .b(_02201_),
    .c(_02202_),
    .y(_02203_)
  );
  al_ao21ftf _07211_ (
    .a(g35),
    .b(\DFF_930.Q ),
    .c(_02203_),
    .y(\DFF_887.D )
  );
  al_mux2l _07212_ (
    .a(\DFF_346.Q ),
    .b(\DFF_764.Q ),
    .s(_01557_),
    .y(_02204_)
  );
  al_mux2h _07213_ (
    .a(\DFF_541.Q ),
    .b(_02204_),
    .s(g35),
    .y(\DFF_346.D )
  );
  al_ao21 _07214_ (
    .a(\DFF_845.Q ),
    .b(_01964_),
    .c(\DFF_1364.Q ),
    .y(_02205_)
  );
  al_ao21ftt _07215_ (
    .a(_01965_),
    .b(_02205_),
    .c(_01963_),
    .y(_02206_)
  );
  al_aoi21ftf _07216_ (
    .a(\DFF_845.Q ),
    .b(_00066_),
    .c(_02206_),
    .y(\DFF_1364.D )
  );
  al_nand3fft _07217_ (
    .a(_01534_),
    .b(\DFF_265.Q ),
    .c(_00974_),
    .y(_02207_)
  );
  al_aoi21ftf _07218_ (
    .a(\DFF_930.Q ),
    .b(_02207_),
    .c(g35),
    .y(_02208_)
  );
  al_oai21 _07219_ (
    .a(_00977_),
    .b(_02207_),
    .c(_02208_),
    .y(_02209_)
  );
  al_ao21ftf _07220_ (
    .a(g35),
    .b(\DFF_273.Q ),
    .c(_02209_),
    .y(\DFF_930.D )
  );
  al_nand3 _07221_ (
    .a(\DFF_1346.Q ),
    .b(_01651_),
    .c(_00689_),
    .y(_02210_)
  );
  al_ao21 _07222_ (
    .a(\DFF_1346.Q ),
    .b(_01651_),
    .c(_00689_),
    .y(_02211_)
  );
  al_nand3 _07223_ (
    .a(g35),
    .b(_02210_),
    .c(_02211_),
    .y(_02212_)
  );
  al_aoi21ftf _07224_ (
    .a(\DFF_926.Q ),
    .b(_00066_),
    .c(_02212_),
    .y(\DFF_1346.D )
  );
  al_nand3fft _07225_ (
    .a(\DFF_598.Q ),
    .b(\DFF_68.Q ),
    .c(\DFF_1098.Q ),
    .y(_02213_)
  );
  al_aoi21ftf _07226_ (
    .a(\DFF_100.Q ),
    .b(_02213_),
    .c(g35),
    .y(_02214_)
  );
  al_ao21ftf _07227_ (
    .a(_02213_),
    .b(_00499_),
    .c(_02214_),
    .y(_02215_)
  );
  al_ao21ftf _07228_ (
    .a(g35),
    .b(\DFF_659.Q ),
    .c(_02215_),
    .y(\DFF_100.D )
  );
  al_nand3 _07229_ (
    .a(_00499_),
    .b(_01745_),
    .c(_01773_),
    .y(_02216_)
  );
  al_ao21 _07230_ (
    .a(_01773_),
    .b(_01745_),
    .c(\DFF_627.Q ),
    .y(_02217_)
  );
  al_nand3 _07231_ (
    .a(g35),
    .b(_02217_),
    .c(_02216_),
    .y(_02218_)
  );
  al_ao21ftf _07232_ (
    .a(g35),
    .b(\DFF_333.Q ),
    .c(_02218_),
    .y(\DFF_627.D )
  );
  al_ao21 _07233_ (
    .a(_01664_),
    .b(_01663_),
    .c(_00066_),
    .y(_02219_)
  );
  al_mux2l _07234_ (
    .a(\DFF_400.Q ),
    .b(\DFF_897.Q ),
    .s(_02219_),
    .y(\DFF_897.D )
  );
  al_nand3 _07235_ (
    .a(_00499_),
    .b(_01763_),
    .c(_00508_),
    .y(_02220_)
  );
  al_ao21 _07236_ (
    .a(_00508_),
    .b(_01763_),
    .c(\DFF_291.Q ),
    .y(_02221_)
  );
  al_nand3 _07237_ (
    .a(g35),
    .b(_02221_),
    .c(_02220_),
    .y(_02222_)
  );
  al_ao21ftf _07238_ (
    .a(g35),
    .b(\DFF_588.Q ),
    .c(_02222_),
    .y(\DFF_291.D )
  );
  al_nand3ftt _07239_ (
    .a(\DFF_467.Q ),
    .b(\DFF_587.Q ),
    .c(\DFF_473.Q ),
    .y(_02223_)
  );
  al_aoi21ftf _07240_ (
    .a(\DFF_1264.Q ),
    .b(_02223_),
    .c(g35),
    .y(_02224_)
  );
  al_ao21ftf _07241_ (
    .a(_02223_),
    .b(_00499_),
    .c(_02224_),
    .y(_02225_)
  );
  al_ao21ftf _07242_ (
    .a(g35),
    .b(\DFF_550.Q ),
    .c(_02225_),
    .y(\DFF_1264.D )
  );
  al_and2 _07243_ (
    .a(\DFF_358.Q ),
    .b(_00603_),
    .y(_02226_)
  );
  al_nand3 _07244_ (
    .a(\DFF_63.Q ),
    .b(\DFF_718.Q ),
    .c(_02226_),
    .y(_02227_)
  );
  al_aoi21ttf _07245_ (
    .a(\DFF_807.Q ),
    .b(_02226_),
    .c(_01505_),
    .y(_02228_)
  );
  al_aoi21ftf _07246_ (
    .a(\DFF_660.Q ),
    .b(_02227_),
    .c(_02228_),
    .y(_02229_)
  );
  al_ao21ftf _07247_ (
    .a(_02227_),
    .b(\DFF_660.Q ),
    .c(_02229_),
    .y(_02230_)
  );
  al_ao21ftf _07248_ (
    .a(g35),
    .b(\DFF_718.Q ),
    .c(_02230_),
    .y(\DFF_660.D )
  );
  al_or2ft _07249_ (
    .a(\DFF_1306.Q ),
    .b(_00358_),
    .y(_02231_)
  );
  al_nand2ft _07250_ (
    .a(\DFF_1306.Q ),
    .b(_00358_),
    .y(_02232_)
  );
  al_nand3 _07251_ (
    .a(g35),
    .b(_02232_),
    .c(_02231_),
    .y(_02233_)
  );
  al_aoi21ftf _07252_ (
    .a(\DFF_679.Q ),
    .b(_00066_),
    .c(_02233_),
    .y(\DFF_1306.D )
  );
  al_nor2 _07253_ (
    .a(\DFF_230.Q ),
    .b(g35),
    .y(_02234_)
  );
  al_mux2l _07254_ (
    .a(\DFF_732.Q ),
    .b(\DFF_1279.Q ),
    .s(\DFF_230.Q ),
    .y(_02235_)
  );
  al_nand3ftt _07255_ (
    .a(_02235_),
    .b(\DFF_1056.Q ),
    .c(_01042_),
    .y(_02236_)
  );
  al_aoi21ftf _07256_ (
    .a(\DFF_1056.Q ),
    .b(_02235_),
    .c(g35),
    .y(_02237_)
  );
  al_aoi21 _07257_ (
    .a(_02237_),
    .b(_02236_),
    .c(_02234_),
    .y(\DFF_1056.D )
  );
  al_mux2l _07258_ (
    .a(\DFF_255.Q ),
    .b(_01153_),
    .s(_01195_),
    .y(_02238_)
  );
  al_mux2h _07259_ (
    .a(\DFF_77.Q ),
    .b(_02238_),
    .s(g35),
    .y(\DFF_255.D )
  );
  al_and2ft _07260_ (
    .a(\DFF_1275.Q ),
    .b(g35),
    .y(_02239_)
  );
  al_nand3ftt _07261_ (
    .a(\DFF_871.Q ),
    .b(\DFF_1017.Q ),
    .c(g35),
    .y(_02240_)
  );
  al_ao21ttf _07262_ (
    .a(\DFF_1017.Q ),
    .b(g35),
    .c(\DFF_871.Q ),
    .y(_02241_)
  );
  al_aoi21 _07263_ (
    .a(_02240_),
    .b(_02241_),
    .c(_02239_),
    .y(\DFF_1017.D )
  );
  al_and2 _07264_ (
    .a(g113),
    .b(g35),
    .y(\DFF_178.D )
  );
  al_and3ftt _07265_ (
    .a(\DFF_563.Q ),
    .b(\DFF_214.Q ),
    .c(\DFF_600.Q ),
    .y(_02242_)
  );
  al_nand3fft _07266_ (
    .a(\DFF_24.Q ),
    .b(\DFF_137.Q ),
    .c(_00718_),
    .y(_02243_)
  );
  al_ao21ftf _07267_ (
    .a(\DFF_24.Q ),
    .b(_00718_),
    .c(\DFF_137.Q ),
    .y(_02244_)
  );
  al_nand3 _07268_ (
    .a(_02242_),
    .b(_02243_),
    .c(_02244_),
    .y(_02245_)
  );
  al_ao21 _07269_ (
    .a(_02242_),
    .b(_01005_),
    .c(\DFF_1382.Q ),
    .y(_02246_)
  );
  al_nand3 _07270_ (
    .a(g35),
    .b(_02246_),
    .c(_02245_),
    .y(_02247_)
  );
  al_ao21ftf _07271_ (
    .a(g35),
    .b(\DFF_98.Q ),
    .c(_02247_),
    .y(\DFF_1382.D )
  );
  al_and2 _07272_ (
    .a(\DFF_328.Q ),
    .b(_01179_),
    .y(_02248_)
  );
  al_nand3 _07273_ (
    .a(\DFF_74.Q ),
    .b(\DFF_157.Q ),
    .c(_02248_),
    .y(_02249_)
  );
  al_nand3 _07274_ (
    .a(\DFF_157.Q ),
    .b(\DFF_328.Q ),
    .c(_01179_),
    .y(_02250_)
  );
  al_ao21ttf _07275_ (
    .a(\DFF_74.Q ),
    .b(_00941_),
    .c(_02250_),
    .y(_02251_)
  );
  al_nand3 _07276_ (
    .a(g35),
    .b(_02251_),
    .c(_02249_),
    .y(_02252_)
  );
  al_ao21ftf _07277_ (
    .a(g35),
    .b(\DFF_157.Q ),
    .c(_02252_),
    .y(\DFF_74.D )
  );
  al_oai21ftf _07278_ (
    .a(\DFF_1414.Q ),
    .b(\DFF_492.Q ),
    .c(\DFF_805.Q ),
    .y(_02253_)
  );
  al_nand3ftt _07279_ (
    .a(\DFF_830.Q ),
    .b(g35),
    .c(_02253_),
    .y(_02254_)
  );
  al_ao21ftf _07280_ (
    .a(g35),
    .b(\DFF_492.Q ),
    .c(_02254_),
    .y(\DFF_805.D )
  );
  al_mux2l _07281_ (
    .a(\DFF_760.Q ),
    .b(\DFF_48.Q ),
    .s(\DFF_1269.Q ),
    .y(_02255_)
  );
  al_mux2h _07282_ (
    .a(\DFF_1269.Q ),
    .b(_02255_),
    .s(g35),
    .y(\DFF_753.D )
  );
  al_and2ft _07283_ (
    .a(g35),
    .b(\DFF_846.Q ),
    .y(_02256_)
  );
  al_and3 _07284_ (
    .a(\DFF_792.Q ),
    .b(_00587_),
    .c(_00009_),
    .y(_02257_)
  );
  al_aoi21 _07285_ (
    .a(_02257_),
    .b(_00414_),
    .c(_00066_),
    .y(_02258_)
  );
  al_and3 _07286_ (
    .a(\DFF_792.Q ),
    .b(g25114),
    .c(_00009_),
    .y(_02259_)
  );
  al_nand3 _07287_ (
    .a(\DFF_792.Q ),
    .b(\DFF_846.Q ),
    .c(_00009_),
    .y(_02260_)
  );
  al_aoi21 _07288_ (
    .a(_01327_),
    .b(_02260_),
    .c(_02259_),
    .y(_02261_)
  );
  al_ao21 _07289_ (
    .a(_02261_),
    .b(_02258_),
    .c(_02256_),
    .y(\DFF_449.D )
  );
  al_nand2 _07290_ (
    .a(\DFF_1243.Q ),
    .b(\DFF_649.Q ),
    .y(_02262_)
  );
  al_nor2 _07291_ (
    .a(\DFF_1243.Q ),
    .b(\DFF_649.Q ),
    .y(_02263_)
  );
  al_nand2ft _07292_ (
    .a(_02263_),
    .b(_02262_),
    .y(_02264_)
  );
  al_mux2l _07293_ (
    .a(_02264_),
    .b(\DFF_814.Q ),
    .s(_01890_),
    .y(_02265_)
  );
  al_mux2h _07294_ (
    .a(\DFF_649.Q ),
    .b(_02265_),
    .s(g35),
    .y(\DFF_814.D )
  );
  al_nand2 _07295_ (
    .a(\DFF_768.Q ),
    .b(\DFF_6.Q ),
    .y(_02266_)
  );
  al_nor2 _07296_ (
    .a(\DFF_768.Q ),
    .b(\DFF_6.Q ),
    .y(_02267_)
  );
  al_nand2ft _07297_ (
    .a(_02267_),
    .b(_02266_),
    .y(_02268_)
  );
  al_mux2l _07298_ (
    .a(\DFF_825.Q ),
    .b(_02268_),
    .s(_00564_),
    .y(_02269_)
  );
  al_mux2h _07299_ (
    .a(\DFF_6.Q ),
    .b(_02269_),
    .s(g35),
    .y(\DFF_825.D )
  );
  al_nand3ftt _07300_ (
    .a(\DFF_519.Q ),
    .b(\DFF_385.Q ),
    .c(\DFF_393.Q ),
    .y(_02270_)
  );
  al_aoi21ftf _07301_ (
    .a(\DFF_93.Q ),
    .b(_02270_),
    .c(g35),
    .y(_02271_)
  );
  al_ao21ftf _07302_ (
    .a(_02270_),
    .b(_00499_),
    .c(_02271_),
    .y(_02272_)
  );
  al_ao21ftf _07303_ (
    .a(g35),
    .b(\DFF_1255.Q ),
    .c(_02272_),
    .y(\DFF_93.D )
  );
  al_ao21 _07304_ (
    .a(\DFF_792.Q ),
    .b(_00009_),
    .c(\DFF_846.Q ),
    .y(_02273_)
  );
  al_nand3 _07305_ (
    .a(_02260_),
    .b(_02273_),
    .c(_02258_),
    .y(_02274_)
  );
  al_ao21ftf _07306_ (
    .a(g35),
    .b(\DFF_1285.Q ),
    .c(_02274_),
    .y(\DFF_846.D )
  );
  al_nand2ft _07307_ (
    .a(g35),
    .b(\DFF_728.Q ),
    .y(_02275_)
  );
  al_oa21ftt _07308_ (
    .a(\DFF_109.Q ),
    .b(\DFF_7.Q ),
    .c(g35),
    .y(_02276_)
  );
  al_oa21 _07309_ (
    .a(\DFF_506.Q ),
    .b(_01185_),
    .c(_02276_),
    .y(_02277_)
  );
  al_ao21ftf _07310_ (
    .a(_01231_),
    .b(_02277_),
    .c(_02275_),
    .y(\DFF_506.D )
  );
  al_and3fft _07311_ (
    .a(\DFF_1148.Q ),
    .b(\DFF_717.Q ),
    .c(\DFF_327.Q ),
    .y(_02278_)
  );
  al_ao21ttf _07312_ (
    .a(\DFF_167.Q ),
    .b(_02278_),
    .c(\DFF_822.Q ),
    .y(_02279_)
  );
  al_nand2ft _07313_ (
    .a(\DFF_182.Q ),
    .b(_02278_),
    .y(_02280_)
  );
  al_aoi21 _07314_ (
    .a(_02280_),
    .b(_02279_),
    .c(_00066_),
    .y(\DFF_822.D )
  );
  al_oai21ftt _07315_ (
    .a(g35),
    .b(\DFF_605.Q ),
    .c(\DFF_354.Q ),
    .y(_02281_)
  );
  al_ao21ttf _07316_ (
    .a(\DFF_691.Q ),
    .b(g35),
    .c(_02281_),
    .y(_02282_)
  );
  al_and3 _07317_ (
    .a(\DFF_354.Q ),
    .b(\DFF_605.Q ),
    .c(g35),
    .y(_02283_)
  );
  al_aoi21ttf _07318_ (
    .a(\DFF_691.Q ),
    .b(_02283_),
    .c(_02282_),
    .y(\DFF_691.D )
  );
  al_nor2 _07319_ (
    .a(g35),
    .b(\DFF_183.Q ),
    .y(_02284_)
  );
  al_nand2 _07320_ (
    .a(\DFF_920.Q ),
    .b(\DFF_848.Q ),
    .y(_02285_)
  );
  al_nand2 _07321_ (
    .a(\DFF_30.Q ),
    .b(\DFF_17.Q ),
    .y(_02286_)
  );
  al_ao21ttf _07322_ (
    .a(_02285_),
    .b(_02286_),
    .c(_00399_),
    .y(_02287_)
  );
  al_nand2ft _07323_ (
    .a(\DFF_833.Q ),
    .b(\DFF_429.Q ),
    .y(_02288_)
  );
  al_nand2 _07324_ (
    .a(\DFF_1201.Q ),
    .b(\DFF_22.Q ),
    .y(_02289_)
  );
  al_ao21ttf _07325_ (
    .a(\DFF_241.Q ),
    .b(\DFF_1087.Q ),
    .c(_02289_),
    .y(_02290_)
  );
  al_aoi21ftf _07326_ (
    .a(_02288_),
    .b(_02290_),
    .c(_02287_),
    .y(_02291_)
  );
  al_nor2 _07327_ (
    .a(\DFF_429.Q ),
    .b(\DFF_833.Q ),
    .y(_02292_)
  );
  al_and3 _07328_ (
    .a(\DFF_1085.Q ),
    .b(\DFF_1102.Q ),
    .c(_02292_),
    .y(_02293_)
  );
  al_nand2ft _07329_ (
    .a(\DFF_429.Q ),
    .b(\DFF_833.Q ),
    .y(_02294_)
  );
  al_nand2 _07330_ (
    .a(\DFF_737.Q ),
    .b(\DFF_93.Q ),
    .y(_02295_)
  );
  al_nand2 _07331_ (
    .a(\DFF_471.Q ),
    .b(\DFF_279.Q ),
    .y(_02296_)
  );
  al_ao21 _07332_ (
    .a(_02295_),
    .b(_02296_),
    .c(_02294_),
    .y(_02297_)
  );
  al_nand3fft _07333_ (
    .a(\DFF_1320.Q ),
    .b(_02293_),
    .c(_02297_),
    .y(_02298_)
  );
  al_or3fft _07334_ (
    .a(\DFF_192.Q ),
    .b(\DFF_1102.Q ),
    .c(_02288_),
    .y(_02299_)
  );
  al_nand3 _07335_ (
    .a(\DFF_877.Q ),
    .b(\DFF_279.Q ),
    .c(_00399_),
    .y(_02300_)
  );
  al_and3 _07336_ (
    .a(\DFF_1320.Q ),
    .b(_02299_),
    .c(_02300_),
    .y(_02301_)
  );
  al_nand2 _07337_ (
    .a(\DFF_398.Q ),
    .b(\DFF_848.Q ),
    .y(_02302_)
  );
  al_nand2 _07338_ (
    .a(\DFF_30.Q ),
    .b(\DFF_1291.Q ),
    .y(_02303_)
  );
  al_ao21 _07339_ (
    .a(_02302_),
    .b(_02303_),
    .c(_02294_),
    .y(_02304_)
  );
  al_nand2 _07340_ (
    .a(\DFF_267.Q ),
    .b(\DFF_1087.Q ),
    .y(_02305_)
  );
  al_nand2 _07341_ (
    .a(\DFF_526.Q ),
    .b(\DFF_22.Q ),
    .y(_02306_)
  );
  al_ao21ttf _07342_ (
    .a(_02305_),
    .b(_02306_),
    .c(_02292_),
    .y(_02307_)
  );
  al_nand3 _07343_ (
    .a(_02304_),
    .b(_02307_),
    .c(_02301_),
    .y(_02308_)
  );
  al_ao21ftf _07344_ (
    .a(_02298_),
    .b(_02291_),
    .c(_02308_),
    .y(_02309_)
  );
  al_nand2 _07345_ (
    .a(\DFF_183.Q ),
    .b(_01957_),
    .y(_02310_)
  );
  al_and3 _07346_ (
    .a(\DFF_797.Q ),
    .b(\DFF_815.Q ),
    .c(_00399_),
    .y(_02311_)
  );
  al_nor2 _07347_ (
    .a(\DFF_30.Q ),
    .b(\DFF_1320.Q ),
    .y(_02312_)
  );
  al_nand2 _07348_ (
    .a(\DFF_30.Q ),
    .b(\DFF_1320.Q ),
    .y(_02313_)
  );
  al_nand2ft _07349_ (
    .a(_02312_),
    .b(_02313_),
    .y(_02314_)
  );
  al_or3fft _07350_ (
    .a(\DFF_326.Q ),
    .b(\DFF_1058.Q ),
    .c(_02288_),
    .y(_02315_)
  );
  al_and3 _07351_ (
    .a(\DFF_110.Q ),
    .b(\DFF_1255.Q ),
    .c(_02292_),
    .y(_02316_)
  );
  al_and3ftt _07352_ (
    .a(_02316_),
    .b(_02315_),
    .c(_02314_),
    .y(_02317_)
  );
  al_nor3fft _07353_ (
    .a(\DFF_110.Q ),
    .b(\DFF_336.Q ),
    .c(_02288_),
    .y(_02318_)
  );
  al_nor3fft _07354_ (
    .a(\DFF_797.Q ),
    .b(\DFF_949.Q ),
    .c(_02294_),
    .y(_02319_)
  );
  al_nand3 _07355_ (
    .a(\DFF_326.Q ),
    .b(\DFF_854.Q ),
    .c(_02292_),
    .y(_02320_)
  );
  al_and3ftt _07356_ (
    .a(_02312_),
    .b(_02313_),
    .c(_02320_),
    .y(_02321_)
  );
  al_nand3fft _07357_ (
    .a(_02318_),
    .b(_02319_),
    .c(_02321_),
    .y(_02322_)
  );
  al_ao21ftf _07358_ (
    .a(_02311_),
    .b(_02317_),
    .c(_02322_),
    .y(_02323_)
  );
  al_nand3 _07359_ (
    .a(_02310_),
    .b(_02323_),
    .c(_02309_),
    .y(_02324_)
  );
  al_nand2 _07360_ (
    .a(_01956_),
    .b(_02324_),
    .y(_02325_)
  );
  al_oa21ftf _07361_ (
    .a(\DFF_249.Q ),
    .b(_01956_),
    .c(_00066_),
    .y(_02326_)
  );
  al_aoi21 _07362_ (
    .a(_02326_),
    .b(_02325_),
    .c(_02284_),
    .y(\DFF_249.D )
  );
  al_nand3fft _07363_ (
    .a(\DFF_519.Q ),
    .b(\DFF_385.Q ),
    .c(\DFF_393.Q ),
    .y(_02327_)
  );
  al_aoi21ftf _07364_ (
    .a(\DFF_526.Q ),
    .b(_02327_),
    .c(g35),
    .y(_02328_)
  );
  al_ao21ftf _07365_ (
    .a(_02327_),
    .b(_00499_),
    .c(_02328_),
    .y(_02329_)
  );
  al_ao21ftf _07366_ (
    .a(g35),
    .b(\DFF_877.Q ),
    .c(_02329_),
    .y(\DFF_526.D )
  );
  al_oai21ftf _07367_ (
    .a(\DFF_1275.Q ),
    .b(\DFF_1008.Q ),
    .c(\DFF_740.Q ),
    .y(_02330_)
  );
  al_ao21 _07368_ (
    .a(\DFF_937.Q ),
    .b(_02330_),
    .c(_00066_),
    .y(_02331_)
  );
  al_ao21ftf _07369_ (
    .a(_02239_),
    .b(\DFF_740.Q ),
    .c(_02331_),
    .y(\DFF_1092.D )
  );
  al_mux2h _07370_ (
    .a(\DFF_1271.Q ),
    .b(_02006_),
    .s(g35),
    .y(\DFF_466.D )
  );
  al_mux2l _07371_ (
    .a(\DFF_177.Q ),
    .b(\DFF_161.Q ),
    .s(g35),
    .y(\DFF_177.D )
  );
  al_mux2l _07372_ (
    .a(\DFF_324.Q ),
    .b(\DFF_972.Q ),
    .s(_01174_),
    .y(\DFF_972.D )
  );
  al_nand3fft _07373_ (
    .a(g73),
    .b(\DFF_1425.Q ),
    .c(g72),
    .y(_02332_)
  );
  al_mux2l _07374_ (
    .a(_02332_),
    .b(\DFF_744.Q ),
    .s(_01208_),
    .y(\DFF_384.D )
  );
  al_and3 _07375_ (
    .a(g35),
    .b(_00933_),
    .c(_00929_),
    .y(\DFF_128.D )
  );
  al_nand3fft _07376_ (
    .a(\DFF_221.Q ),
    .b(g73),
    .c(g72),
    .y(_02333_)
  );
  al_mux2l _07377_ (
    .a(_02333_),
    .b(\DFF_352.Q ),
    .s(_01208_),
    .y(\DFF_744.D )
  );
  al_and2ft _07378_ (
    .a(\DFF_1066.Q ),
    .b(\DFF_651.Q ),
    .y(_02334_)
  );
  al_nand2ft _07379_ (
    .a(\DFF_651.Q ),
    .b(\DFF_1066.Q ),
    .y(_02335_)
  );
  al_nand2ft _07380_ (
    .a(_02334_),
    .b(_02335_),
    .y(_02336_)
  );
  al_mux2l _07381_ (
    .a(\DFF_1021.Q ),
    .b(_02336_),
    .s(_01691_),
    .y(_02337_)
  );
  al_mux2h _07382_ (
    .a(\DFF_1066.Q ),
    .b(_02337_),
    .s(g35),
    .y(\DFF_1021.D )
  );
  al_aoi21ttf _07383_ (
    .a(_00469_),
    .b(_00584_),
    .c(\DFF_935.Q ),
    .y(_02338_)
  );
  al_and3 _07384_ (
    .a(\DFF_1185.Q ),
    .b(\DFF_198.Q ),
    .c(_00412_),
    .y(_02339_)
  );
  al_ao21ttf _07385_ (
    .a(_02339_),
    .b(_02338_),
    .c(\DFF_716.Q ),
    .y(_02340_)
  );
  al_ao21 _07386_ (
    .a(_02339_),
    .b(_02338_),
    .c(_00066_),
    .y(_02341_)
  );
  al_nand2ft _07387_ (
    .a(\DFF_755.Q ),
    .b(g35),
    .y(_02342_)
  );
  al_ao21ftf _07388_ (
    .a(_02342_),
    .b(\DFF_433.Q ),
    .c(_02341_),
    .y(_02343_)
  );
  al_and3ftt _07389_ (
    .a(\DFF_433.Q ),
    .b(_02342_),
    .c(_02341_),
    .y(_02344_)
  );
  al_aoi21 _07390_ (
    .a(_02340_),
    .b(_02343_),
    .c(_02344_),
    .y(\DFF_716.D )
  );
  al_inv _07391_ (
    .a(\DFF_594.Q ),
    .y(_02345_)
  );
  al_and2 _07392_ (
    .a(\DFF_713.Q ),
    .b(_00641_),
    .y(_02346_)
  );
  al_and2 _07393_ (
    .a(_00322_),
    .b(_00328_),
    .y(_02347_)
  );
  al_nand3 _07394_ (
    .a(\DFF_1181.Q ),
    .b(_00604_),
    .c(_02347_),
    .y(_02348_)
  );
  al_oa21ftf _07395_ (
    .a(\DFF_402.Q ),
    .b(_00641_),
    .c(_00066_),
    .y(_02349_)
  );
  al_ao21ttf _07396_ (
    .a(_02346_),
    .b(_02348_),
    .c(_02349_),
    .y(_02350_)
  );
  al_aoi21ftf _07397_ (
    .a(g35),
    .b(_02345_),
    .c(_02350_),
    .y(\DFF_402.D )
  );
  al_nand3fft _07398_ (
    .a(_01884_),
    .b(_01885_),
    .c(_01889_),
    .y(_02351_)
  );
  al_aoi21ftf _07399_ (
    .a(\DFF_306.Q ),
    .b(_02351_),
    .c(g35),
    .y(_02352_)
  );
  al_oai21 _07400_ (
    .a(_01892_),
    .b(_02351_),
    .c(_02352_),
    .y(_02353_)
  );
  al_ao21ftf _07401_ (
    .a(g35),
    .b(\DFF_173.Q ),
    .c(_02353_),
    .y(\DFF_306.D )
  );
  al_mux2l _07402_ (
    .a(\DFF_541.Q ),
    .b(\DFF_380.Q ),
    .s(_01557_),
    .y(_02354_)
  );
  al_mux2h _07403_ (
    .a(\DFF_362.Q ),
    .b(_02354_),
    .s(g35),
    .y(\DFF_541.D )
  );
  al_oa21ftt _07404_ (
    .a(g35),
    .b(\DFF_701.Q ),
    .c(\DFF_523.Q ),
    .y(_02355_)
  );
  al_aoi21ftf _07405_ (
    .a(\DFF_939.Q ),
    .b(g35),
    .c(_02355_),
    .y(_02356_)
  );
  al_or3fft _07406_ (
    .a(\DFF_540.Q ),
    .b(g35),
    .c(_02356_),
    .y(_02357_)
  );
  al_aoi21ftf _07407_ (
    .a(_00066_),
    .b(\DFF_540.Q ),
    .c(_02356_),
    .y(_02358_)
  );
  al_nand2ft _07408_ (
    .a(_02358_),
    .b(_02357_),
    .y(\DFF_540.D )
  );
  al_oai21ftt _07409_ (
    .a(g35),
    .b(_00546_),
    .c(\DFF_1167.Q ),
    .y(_02359_)
  );
  al_and2ft _07410_ (
    .a(\DFF_552.Q ),
    .b(\DFF_1037.Q ),
    .y(_02360_)
  );
  al_nand2 _07411_ (
    .a(_02360_),
    .b(_00546_),
    .y(_02361_)
  );
  al_nand3 _07412_ (
    .a(\DFF_977.Q ),
    .b(g35),
    .c(_02361_),
    .y(_02362_)
  );
  al_and2ft _07413_ (
    .a(_02359_),
    .b(_02362_),
    .y(_02363_)
  );
  al_or2ft _07414_ (
    .a(_02359_),
    .b(_02362_),
    .y(_02364_)
  );
  al_nand2ft _07415_ (
    .a(_02363_),
    .b(_02364_),
    .y(\DFF_977.D )
  );
  al_and2 _07416_ (
    .a(g35),
    .b(_01442_),
    .y(_02365_)
  );
  al_and3ftt _07417_ (
    .a(\DFF_734.Q ),
    .b(_01441_),
    .c(_02365_),
    .y(\DFF_734.D )
  );
  al_mux2h _07418_ (
    .a(\DFF_57.Q ),
    .b(_01943_),
    .s(g35),
    .y(\DFF_1377.D )
  );
  al_oai21ftt _07419_ (
    .a(\DFF_1131.Q ),
    .b(\DFF_195.Q ),
    .c(g35),
    .y(_02366_)
  );
  al_ao21ftf _07420_ (
    .a(g35),
    .b(\DFF_948.Q ),
    .c(_02366_),
    .y(\DFF_195.D )
  );
  al_and2 _07421_ (
    .a(\DFF_587.Q ),
    .b(\DFF_467.Q ),
    .y(_02367_)
  );
  al_or3 _07422_ (
    .a(\DFF_784.Q ),
    .b(\DFF_473.Q ),
    .c(\DFF_776.Q ),
    .y(_02368_)
  );
  al_nand3ftt _07423_ (
    .a(_02368_),
    .b(_02367_),
    .c(_00499_),
    .y(_02369_)
  );
  al_ao21ftt _07424_ (
    .a(_02368_),
    .b(_02367_),
    .c(\DFF_91.Q ),
    .y(_02370_)
  );
  al_nand3 _07425_ (
    .a(g35),
    .b(_02369_),
    .c(_02370_),
    .y(_02371_)
  );
  al_ao21ftf _07426_ (
    .a(g35),
    .b(\DFF_1264.Q ),
    .c(_02371_),
    .y(\DFF_91.D )
  );
  al_nand3ftt _07427_ (
    .a(\DFF_1314.Q ),
    .b(g35),
    .c(_00718_),
    .y(_02372_)
  );
  al_aoi21ftf _07428_ (
    .a(\DFF_127.Q ),
    .b(_00066_),
    .c(_02372_),
    .y(\DFF_1314.D )
  );
  al_and2ft _07429_ (
    .a(g35),
    .b(\DFF_50.Q ),
    .y(_02373_)
  );
  al_ao21 _07430_ (
    .a(\DFF_789.Q ),
    .b(_00941_),
    .c(_00952_),
    .y(_02374_)
  );
  al_ao21 _07431_ (
    .a(\DFF_789.Q ),
    .b(_00952_),
    .c(_00066_),
    .y(_02375_)
  );
  al_oai21ftf _07432_ (
    .a(_02374_),
    .b(_02375_),
    .c(_02373_),
    .y(\DFF_789.D )
  );
  al_nand3 _07433_ (
    .a(\DFF_947.Q ),
    .b(\DFF_1219.Q ),
    .c(_00404_),
    .y(_02376_)
  );
  al_and2ft _07434_ (
    .a(\DFF_286.Q ),
    .b(\DFF_517.Q ),
    .y(_02377_)
  );
  al_nand3 _07435_ (
    .a(\DFF_257.Q ),
    .b(\DFF_662.Q ),
    .c(_02377_),
    .y(_02378_)
  );
  al_and3 _07436_ (
    .a(\DFF_5.Q ),
    .b(_02378_),
    .c(_02376_),
    .y(_02379_)
  );
  al_nor2 _07437_ (
    .a(\DFF_286.Q ),
    .b(\DFF_517.Q ),
    .y(_02380_)
  );
  al_nand2 _07438_ (
    .a(\DFF_340.Q ),
    .b(\DFF_642.Q ),
    .y(_02381_)
  );
  al_nand2 _07439_ (
    .a(\DFF_995.Q ),
    .b(\DFF_590.Q ),
    .y(_02382_)
  );
  al_ao21ttf _07440_ (
    .a(_02381_),
    .b(_02382_),
    .c(_02380_),
    .y(_02383_)
  );
  al_nand2ft _07441_ (
    .a(\DFF_517.Q ),
    .b(\DFF_286.Q ),
    .y(_02384_)
  );
  al_nand2 _07442_ (
    .a(\DFF_479.Q ),
    .b(\DFF_367.Q ),
    .y(_02385_)
  );
  al_nand2 _07443_ (
    .a(\DFF_1001.Q ),
    .b(\DFF_1350.Q ),
    .y(_02386_)
  );
  al_ao21 _07444_ (
    .a(_02385_),
    .b(_02386_),
    .c(_02384_),
    .y(_02387_)
  );
  al_nand3 _07445_ (
    .a(_02383_),
    .b(_02387_),
    .c(_02379_),
    .y(_02388_)
  );
  al_nand2 _07446_ (
    .a(\DFF_312.Q ),
    .b(\DFF_642.Q ),
    .y(_02389_)
  );
  al_ao21ttf _07447_ (
    .a(\DFF_1264.Q ),
    .b(\DFF_995.Q ),
    .c(_02389_),
    .y(_02390_)
  );
  al_and3 _07448_ (
    .a(\DFF_1160.Q ),
    .b(\DFF_662.Q ),
    .c(_02380_),
    .y(_02391_)
  );
  al_ao21 _07449_ (
    .a(_02377_),
    .b(_02390_),
    .c(_02391_),
    .y(_02392_)
  );
  al_inv _07450_ (
    .a(\DFF_5.Q ),
    .y(_02393_)
  );
  al_nand2 _07451_ (
    .a(\DFF_785.Q ),
    .b(\DFF_156.Q ),
    .y(_02394_)
  );
  al_nand2 _07452_ (
    .a(\DFF_550.Q ),
    .b(\DFF_1219.Q ),
    .y(_02395_)
  );
  al_ao21 _07453_ (
    .a(_02394_),
    .b(_02395_),
    .c(_02384_),
    .y(_02396_)
  );
  al_nand2 _07454_ (
    .a(\DFF_1001.Q ),
    .b(\DFF_91.Q ),
    .y(_02397_)
  );
  al_nand2 _07455_ (
    .a(\DFF_986.Q ),
    .b(\DFF_367.Q ),
    .y(_02398_)
  );
  al_aoi21ttf _07456_ (
    .a(_02397_),
    .b(_02398_),
    .c(_00404_),
    .y(_02399_)
  );
  al_nor3fft _07457_ (
    .a(_02393_),
    .b(_02396_),
    .c(_02399_),
    .y(_02400_)
  );
  al_ao21ftf _07458_ (
    .a(_02392_),
    .b(_02400_),
    .c(_02388_),
    .y(_02401_)
  );
  al_nand2 _07459_ (
    .a(\DFF_253.Q ),
    .b(_00983_),
    .y(_02402_)
  );
  al_and3 _07460_ (
    .a(\DFF_181.Q ),
    .b(\DFF_1317.Q ),
    .c(_02380_),
    .y(_02403_)
  );
  al_and3 _07461_ (
    .a(\DFF_305.Q ),
    .b(\DFF_868.Q ),
    .c(_00404_),
    .y(_02404_)
  );
  al_nand3 _07462_ (
    .a(\DFF_401.Q ),
    .b(\DFF_1128.Q ),
    .c(_02377_),
    .y(_02405_)
  );
  al_and2ft _07463_ (
    .a(\DFF_5.Q ),
    .b(\DFF_1001.Q ),
    .y(_02406_)
  );
  al_nand2ft _07464_ (
    .a(\DFF_1001.Q ),
    .b(\DFF_5.Q ),
    .y(_02407_)
  );
  al_and3ftt _07465_ (
    .a(_02406_),
    .b(_02407_),
    .c(_02405_),
    .y(_02408_)
  );
  al_nand3fft _07466_ (
    .a(_02403_),
    .b(_02404_),
    .c(_02408_),
    .y(_02409_)
  );
  al_and3 _07467_ (
    .a(\DFF_401.Q ),
    .b(\DFF_917.Q ),
    .c(_02380_),
    .y(_02410_)
  );
  al_nand2ft _07468_ (
    .a(_02406_),
    .b(_02407_),
    .y(_02411_)
  );
  al_and3 _07469_ (
    .a(\DFF_181.Q ),
    .b(\DFF_414.Q ),
    .c(_02377_),
    .y(_02412_)
  );
  al_or3fft _07470_ (
    .a(\DFF_305.Q ),
    .b(\DFF_1013.Q ),
    .c(_02384_),
    .y(_02413_)
  );
  al_and3ftt _07471_ (
    .a(_02412_),
    .b(_02413_),
    .c(_02411_),
    .y(_02414_)
  );
  al_ao21ftf _07472_ (
    .a(_02410_),
    .b(_02414_),
    .c(_02409_),
    .y(_02415_)
  );
  al_nand3 _07473_ (
    .a(_02402_),
    .b(_02415_),
    .c(_02401_),
    .y(_02416_)
  );
  al_nand2 _07474_ (
    .a(_00585_),
    .b(_02416_),
    .y(_02417_)
  );
  al_nand3 _07475_ (
    .a(\DFF_546.Q ),
    .b(_00984_),
    .c(_02417_),
    .y(_02418_)
  );
  al_ao21 _07476_ (
    .a(\DFF_546.Q ),
    .b(_00984_),
    .c(_02417_),
    .y(_02419_)
  );
  al_nand3 _07477_ (
    .a(g35),
    .b(_02418_),
    .c(_02419_),
    .y(_02420_)
  );
  al_aoi21ftf _07478_ (
    .a(\DFF_87.Q ),
    .b(_00066_),
    .c(_02420_),
    .y(\DFF_546.D )
  );
  al_nand3 _07479_ (
    .a(\DFF_1371.Q ),
    .b(\DFF_375.Q ),
    .c(\DFF_372.Q ),
    .y(_02421_)
  );
  al_nand2 _07480_ (
    .a(g35),
    .b(_02421_),
    .y(_02422_)
  );
  al_aoi21ttf _07481_ (
    .a(\DFF_1194.Q ),
    .b(g35),
    .c(\DFF_1313.Q ),
    .y(_02423_)
  );
  al_mux2l _07482_ (
    .a(_02423_),
    .b(\DFF_1194.Q ),
    .s(_02422_),
    .y(\DFF_1194.D )
  );
  al_ao21ttf _07483_ (
    .a(\DFF_1094.Q ),
    .b(_01210_),
    .c(\DFF_580.Q ),
    .y(_02424_)
  );
  al_nand2ft _07484_ (
    .a(\DFF_98.Q ),
    .b(_01210_),
    .y(_02425_)
  );
  al_aoi21 _07485_ (
    .a(_02425_),
    .b(_02424_),
    .c(_00066_),
    .y(\DFF_580.D )
  );
  al_and2ft _07486_ (
    .a(\DFF_467.Q ),
    .b(\DFF_587.Q ),
    .y(_02426_)
  );
  al_nand3ftt _07487_ (
    .a(_02368_),
    .b(_00499_),
    .c(_02426_),
    .y(_02427_)
  );
  al_ao21ftt _07488_ (
    .a(_02368_),
    .b(_02426_),
    .c(\DFF_312.Q ),
    .y(_02428_)
  );
  al_nand3 _07489_ (
    .a(g35),
    .b(_02427_),
    .c(_02428_),
    .y(_02429_)
  );
  al_ao21ftf _07490_ (
    .a(g35),
    .b(\DFF_156.Q ),
    .c(_02429_),
    .y(\DFF_312.D )
  );
  al_and3 _07491_ (
    .a(\DFF_874.Q ),
    .b(\DFF_1090.Q ),
    .c(_01190_),
    .y(_02430_)
  );
  al_ao21 _07492_ (
    .a(\DFF_966.Q ),
    .b(_02430_),
    .c(_01230_),
    .y(_02431_)
  );
  al_or3fft _07493_ (
    .a(g35),
    .b(_02431_),
    .c(_01236_),
    .y(_02432_)
  );
  al_ao21ftf _07494_ (
    .a(g35),
    .b(\DFF_966.Q ),
    .c(_02432_),
    .y(\DFF_89.D )
  );
  al_nor3ftt _07495_ (
    .a(\DFF_559.Q ),
    .b(_00499_),
    .c(_00378_),
    .y(_02433_)
  );
  al_oa21ftt _07496_ (
    .a(\DFF_559.Q ),
    .b(_00378_),
    .c(_00499_),
    .y(_02434_)
  );
  al_nor3ftt _07497_ (
    .a(g35),
    .b(_02433_),
    .c(_02434_),
    .y(\DFF_559.D )
  );
  al_nor2 _07498_ (
    .a(\DFF_36.Q ),
    .b(g35),
    .y(_02435_)
  );
  al_mux2l _07499_ (
    .a(\DFF_1298.Q ),
    .b(\DFF_805.Q ),
    .s(\DFF_36.Q ),
    .y(_02436_)
  );
  al_nand3ftt _07500_ (
    .a(_02436_),
    .b(\DFF_762.Q ),
    .c(_01455_),
    .y(_02437_)
  );
  al_aoi21ftf _07501_ (
    .a(\DFF_762.Q ),
    .b(_02436_),
    .c(g35),
    .y(_02438_)
  );
  al_aoi21 _07502_ (
    .a(_02438_),
    .b(_02437_),
    .c(_02435_),
    .y(\DFF_762.D )
  );
  al_and2ft _07503_ (
    .a(g35),
    .b(\DFF_1281.Q ),
    .y(_02439_)
  );
  al_nand3 _07504_ (
    .a(\DFF_1344.Q ),
    .b(_01061_),
    .c(_01056_),
    .y(_02440_)
  );
  al_nand2ft _07505_ (
    .a(\DFF_1266.Q ),
    .b(\DFF_1281.Q ),
    .y(_02441_)
  );
  al_nand2ft _07506_ (
    .a(\DFF_1281.Q ),
    .b(\DFF_1266.Q ),
    .y(_02442_)
  );
  al_or3fft _07507_ (
    .a(_02441_),
    .b(_02442_),
    .c(_02440_),
    .y(_02443_)
  );
  al_aoi21ftf _07508_ (
    .a(\DFF_583.Q ),
    .b(_02440_),
    .c(g35),
    .y(_02444_)
  );
  al_ao21 _07509_ (
    .a(_02443_),
    .b(_02444_),
    .c(_02439_),
    .y(\DFF_583.D )
  );
  al_nand3ftt _07510_ (
    .a(_01796_),
    .b(g25167),
    .c(_01056_),
    .y(_02445_)
  );
  al_ao21 _07511_ (
    .a(g25167),
    .b(_01056_),
    .c(\DFF_164.Q ),
    .y(_02446_)
  );
  al_nand3 _07512_ (
    .a(g35),
    .b(_02445_),
    .c(_02446_),
    .y(_02447_)
  );
  al_ao21ftf _07513_ (
    .a(g35),
    .b(\DFF_1180.Q ),
    .c(_02447_),
    .y(\DFF_164.D )
  );
  al_and2ft _07514_ (
    .a(g35),
    .b(\DFF_487.Q ),
    .y(_02448_)
  );
  al_nand3 _07515_ (
    .a(_00442_),
    .b(_00577_),
    .c(_00424_),
    .y(_02449_)
  );
  al_oai21ftf _07516_ (
    .a(\DFF_189.Q ),
    .b(\DFF_623.Q ),
    .c(\DFF_562.Q ),
    .y(_02450_)
  );
  al_nand3 _07517_ (
    .a(_00758_),
    .b(_02450_),
    .c(_02449_),
    .y(_02451_)
  );
  al_inv _07518_ (
    .a(\DFF_623.Q ),
    .y(_02452_)
  );
  al_oa21ftf _07519_ (
    .a(_02452_),
    .b(_00758_),
    .c(_00066_),
    .y(_02453_)
  );
  al_ao21 _07520_ (
    .a(_02453_),
    .b(_02451_),
    .c(_02448_),
    .y(\DFF_623.D )
  );
  al_mux2l _07521_ (
    .a(\DFF_311.Q ),
    .b(\DFF_1151.Q ),
    .s(g35),
    .y(\DFF_311.D )
  );
  al_mux2l _07522_ (
    .a(\DFF_1320.Q ),
    .b(\DFF_396.Q ),
    .s(g35),
    .y(\DFF_376.D )
  );
  al_and2 _07523_ (
    .a(\DFF_519.Q ),
    .b(g35),
    .y(\DFF_85.D )
  );
  al_or2 _07524_ (
    .a(_00066_),
    .b(_01890_),
    .y(_02454_)
  );
  al_mux2l _07525_ (
    .a(\DFF_1243.Q ),
    .b(\DFF_649.Q ),
    .s(_02454_),
    .y(\DFF_649.D )
  );
  al_and2 _07526_ (
    .a(g35),
    .b(g64),
    .y(\DFF_752.D )
  );
  al_mux2l _07527_ (
    .a(g6750),
    .b(\DFF_911.Q ),
    .s(g35),
    .y(\DFF_129.D )
  );
  al_or2 _07528_ (
    .a(_00066_),
    .b(_01858_),
    .y(_02455_)
  );
  al_mux2l _07529_ (
    .a(\DFF_232.Q ),
    .b(\DFF_903.Q ),
    .s(_02455_),
    .y(\DFF_903.D )
  );
  al_mux2l _07530_ (
    .a(\DFF_1230.Q ),
    .b(\DFF_1139.Q ),
    .s(_00853_),
    .y(\DFF_1139.D )
  );
  al_nand3ftt _07531_ (
    .a(_02030_),
    .b(_00499_),
    .c(_02011_),
    .y(_02456_)
  );
  al_ao21ftt _07532_ (
    .a(_02030_),
    .b(_02011_),
    .c(\DFF_707.Q ),
    .y(_02457_)
  );
  al_nand3 _07533_ (
    .a(g35),
    .b(_02456_),
    .c(_02457_),
    .y(_02458_)
  );
  al_ao21ftf _07534_ (
    .a(g35),
    .b(\DFF_199.Q ),
    .c(_02458_),
    .y(\DFF_707.D )
  );
  al_or2 _07535_ (
    .a(\DFF_1060.Q ),
    .b(_00475_),
    .y(_02459_)
  );
  al_nand3 _07536_ (
    .a(_00489_),
    .b(_02459_),
    .c(_00495_),
    .y(_02460_)
  );
  al_ao21ftf _07537_ (
    .a(g35),
    .b(\DFF_359.Q ),
    .c(_02460_),
    .y(\DFF_1060.D )
  );
  al_mux2l _07538_ (
    .a(\DFF_161.Q ),
    .b(\DFF_1193.Q ),
    .s(g35),
    .y(\DFF_161.D )
  );
  al_oai21ftf _07539_ (
    .a(\DFF_218.Q ),
    .b(\DFF_1424.D ),
    .c(\DFF_914.Q ),
    .y(_02461_)
  );
  al_nand3 _07540_ (
    .a(\DFF_1199.Q ),
    .b(\DFF_231.Q ),
    .c(\DFF_892.Q ),
    .y(_02462_)
  );
  al_oa21ttf _07541_ (
    .a(\DFF_1199.Q ),
    .b(\DFF_892.Q ),
    .c(\DFF_847.Q ),
    .y(_02463_)
  );
  al_ao21 _07542_ (
    .a(_02462_),
    .b(_02463_),
    .c(\DFF_218.Q ),
    .y(_02464_)
  );
  al_ao21ftf _07543_ (
    .a(_00464_),
    .b(_02461_),
    .c(_02464_),
    .y(_02465_)
  );
  al_or3 _07544_ (
    .a(\DFF_160.Q ),
    .b(\DFF_935.Q ),
    .c(\DFF_130.Q ),
    .y(_02466_)
  );
  al_or2 _07545_ (
    .a(\DFF_99.Q ),
    .b(_02466_),
    .y(_02467_)
  );
  al_and3fft _07546_ (
    .a(\DFF_1199.Q ),
    .b(\DFF_892.Q ),
    .c(\DFF_766.Q ),
    .y(_02468_)
  );
  al_aoi21 _07547_ (
    .a(\DFF_721.Q ),
    .b(_00470_),
    .c(_02468_),
    .y(_02469_)
  );
  al_nand3ftt _07548_ (
    .a(\DFF_892.Q ),
    .b(\DFF_1199.Q ),
    .c(\DFF_855.Q ),
    .y(_02470_)
  );
  al_nand3 _07549_ (
    .a(\DFF_1199.Q ),
    .b(\DFF_892.Q ),
    .c(\DFF_276.Q ),
    .y(_02471_)
  );
  al_and3 _07550_ (
    .a(_02470_),
    .b(_02471_),
    .c(_02469_),
    .y(_02472_)
  );
  al_nand2ft _07551_ (
    .a(\DFF_1424.D ),
    .b(_02472_),
    .y(_02473_)
  );
  al_nand2ft _07552_ (
    .a(_02472_),
    .b(\DFF_1424.D ),
    .y(_02474_)
  );
  al_nand3 _07553_ (
    .a(_00583_),
    .b(_02473_),
    .c(_02474_),
    .y(_02475_)
  );
  al_nand3ftt _07554_ (
    .a(_02467_),
    .b(_02465_),
    .c(_02475_),
    .y(_02476_)
  );
  al_nand2 _07555_ (
    .a(\DFF_714.Q ),
    .b(\DFF_935.Q ),
    .y(_02477_)
  );
  al_aoi21ttf _07556_ (
    .a(\DFF_535.Q ),
    .b(\DFF_160.Q ),
    .c(_02477_),
    .y(_02478_)
  );
  al_nand2ft _07557_ (
    .a(\DFF_857.Q ),
    .b(\DFF_99.Q ),
    .y(_02479_)
  );
  al_ao21ftf _07558_ (
    .a(\DFF_697.Q ),
    .b(\DFF_130.Q ),
    .c(_02479_),
    .y(_02480_)
  );
  al_nand3ftt _07559_ (
    .a(_02480_),
    .b(_02467_),
    .c(_02478_),
    .y(_02481_)
  );
  al_and3 _07560_ (
    .a(g35),
    .b(_02481_),
    .c(_02476_),
    .y(\DFF_221.D )
  );
  al_nand3 _07561_ (
    .a(\DFF_1321.Q ),
    .b(_01297_),
    .c(_00899_),
    .y(_02482_)
  );
  al_oai21 _07562_ (
    .a(\DFF_1321.Q ),
    .b(_01297_),
    .c(_02482_),
    .y(_02483_)
  );
  al_mux2h _07563_ (
    .a(\DFF_712.Q ),
    .b(_02483_),
    .s(g35),
    .y(\DFF_1321.D )
  );
  al_ao21ttf _07564_ (
    .a(g35),
    .b(_00718_),
    .c(\DFF_867.Q ),
    .y(_02484_)
  );
  al_aoi21 _07565_ (
    .a(g35),
    .b(_01464_),
    .c(_02484_),
    .y(\DFF_758.D )
  );
  al_and3 _07566_ (
    .a(\DFF_283.Q ),
    .b(g35),
    .c(_02056_),
    .y(_02485_)
  );
  al_nand2ft _07567_ (
    .a(_00840_),
    .b(_00838_),
    .y(_02486_)
  );
  al_ao21ftf _07568_ (
    .a(\DFF_979.Q ),
    .b(_01476_),
    .c(_02486_),
    .y(_02487_)
  );
  al_oa21 _07569_ (
    .a(\DFF_698.Q ),
    .b(\DFF_511.Q ),
    .c(g35),
    .y(_02488_)
  );
  al_ao21 _07570_ (
    .a(_02488_),
    .b(_02487_),
    .c(_02485_),
    .y(\DFF_283.D )
  );
  al_ao21ftt _07571_ (
    .a(g35),
    .b(\DFF_221.Q ),
    .c(\DFF_221.D ),
    .y(\DFF_439.D )
  );
  al_and2ft _07572_ (
    .a(\DFF_1252.Q ),
    .b(\DFF_1283.Q ),
    .y(_02489_)
  );
  al_nand2 _07573_ (
    .a(\DFF_151.Q ),
    .b(\DFF_1352.Q ),
    .y(_02490_)
  );
  al_nand2 _07574_ (
    .a(\DFF_172.Q ),
    .b(\DFF_666.Q ),
    .y(_02491_)
  );
  al_ao21ttf _07575_ (
    .a(_02490_),
    .b(_02491_),
    .c(_02489_),
    .y(_02492_)
  );
  al_or2 _07576_ (
    .a(\DFF_1252.Q ),
    .b(\DFF_1283.Q ),
    .y(_02493_)
  );
  al_or3fft _07577_ (
    .a(\DFF_1355.Q ),
    .b(\DFF_1262.Q ),
    .c(_02493_),
    .y(_02494_)
  );
  al_and3 _07578_ (
    .a(_00727_),
    .b(_02494_),
    .c(_02492_),
    .y(_02495_)
  );
  al_nand2 _07579_ (
    .a(\DFF_392.Q ),
    .b(\DFF_695.Q ),
    .y(_02496_)
  );
  al_nand2 _07580_ (
    .a(\DFF_46.Q ),
    .b(\DFF_1007.Q ),
    .y(_02497_)
  );
  al_ao21 _07581_ (
    .a(_02496_),
    .b(_02497_),
    .c(_00407_),
    .y(_02498_)
  );
  al_nand2ft _07582_ (
    .a(\DFF_1283.Q ),
    .b(\DFF_1252.Q ),
    .y(_02499_)
  );
  al_nand2 _07583_ (
    .a(\DFF_219.Q ),
    .b(\DFF_783.Q ),
    .y(_02500_)
  );
  al_ao21ttf _07584_ (
    .a(\DFF_101.Q ),
    .b(\DFF_84.Q ),
    .c(_02500_),
    .y(_02501_)
  );
  al_ao21ftf _07585_ (
    .a(_02499_),
    .b(_02501_),
    .c(_02498_),
    .y(_02502_)
  );
  al_or3fft _07586_ (
    .a(\DFF_884.Q ),
    .b(\DFF_783.Q ),
    .c(_00407_),
    .y(_02503_)
  );
  al_nand3 _07587_ (
    .a(\DFF_51.Q ),
    .b(\DFF_1262.Q ),
    .c(_02489_),
    .y(_02504_)
  );
  al_and3 _07588_ (
    .a(\DFF_599.Q ),
    .b(_02504_),
    .c(_02503_),
    .y(_02505_)
  );
  al_nand2 _07589_ (
    .a(\DFF_333.Q ),
    .b(\DFF_1352.Q ),
    .y(_02506_)
  );
  al_nand2 _07590_ (
    .a(\DFF_307.Q ),
    .b(\DFF_666.Q ),
    .y(_02507_)
  );
  al_ao21 _07591_ (
    .a(_02506_),
    .b(_02507_),
    .c(_02493_),
    .y(_02508_)
  );
  al_nand2 _07592_ (
    .a(\DFF_627.Q ),
    .b(\DFF_695.Q ),
    .y(_02509_)
  );
  al_nand2 _07593_ (
    .a(\DFF_46.Q ),
    .b(\DFF_938.Q ),
    .y(_02510_)
  );
  al_ao21 _07594_ (
    .a(_02509_),
    .b(_02510_),
    .c(_02499_),
    .y(_02511_)
  );
  al_nand3 _07595_ (
    .a(_02508_),
    .b(_02511_),
    .c(_02505_),
    .y(_02512_)
  );
  al_ao21ftf _07596_ (
    .a(_02502_),
    .b(_02495_),
    .c(_02512_),
    .y(_02513_)
  );
  al_nor3fft _07597_ (
    .a(\DFF_1335.Q ),
    .b(\DFF_895.Q ),
    .c(_02493_),
    .y(_02514_)
  );
  al_and2ft _07598_ (
    .a(\DFF_599.Q ),
    .b(\DFF_46.Q ),
    .y(_02515_)
  );
  al_nand2ft _07599_ (
    .a(\DFF_46.Q ),
    .b(\DFF_599.Q ),
    .y(_02516_)
  );
  al_nand2ft _07600_ (
    .a(_02515_),
    .b(_02516_),
    .y(_02517_)
  );
  al_or3fft _07601_ (
    .a(\DFF_117.Q ),
    .b(\DFF_1297.Q ),
    .c(_02499_),
    .y(_02518_)
  );
  al_and3 _07602_ (
    .a(\DFF_263.Q ),
    .b(\DFF_55.Q ),
    .c(_02489_),
    .y(_02519_)
  );
  al_and3ftt _07603_ (
    .a(_02519_),
    .b(_02518_),
    .c(_02517_),
    .y(_02520_)
  );
  al_nor3fft _07604_ (
    .a(\DFF_117.Q ),
    .b(\DFF_71.Q ),
    .c(_00407_),
    .y(_02521_)
  );
  al_nor3fft _07605_ (
    .a(\DFF_263.Q ),
    .b(\DFF_44.Q ),
    .c(_02493_),
    .y(_02522_)
  );
  al_nand3 _07606_ (
    .a(\DFF_1335.Q ),
    .b(\DFF_476.Q ),
    .c(_02489_),
    .y(_02523_)
  );
  al_and3ftt _07607_ (
    .a(_02515_),
    .b(_02516_),
    .c(_02523_),
    .y(_02524_)
  );
  al_nand3fft _07608_ (
    .a(_02521_),
    .b(_02522_),
    .c(_02524_),
    .y(_02525_)
  );
  al_ao21ftf _07609_ (
    .a(_02514_),
    .b(_02520_),
    .c(_02525_),
    .y(_02526_)
  );
  al_aoi21ttf _07610_ (
    .a(\DFF_1423.Q ),
    .b(_01690_),
    .c(_02526_),
    .y(_02527_)
  );
  al_ao21ttf _07611_ (
    .a(_02513_),
    .b(_02527_),
    .c(_01689_),
    .y(_02528_)
  );
  al_nand3 _07612_ (
    .a(\DFF_1066.Q ),
    .b(_01691_),
    .c(_02528_),
    .y(_02529_)
  );
  al_ao21 _07613_ (
    .a(\DFF_1066.Q ),
    .b(_01691_),
    .c(_02528_),
    .y(_02530_)
  );
  al_nand3 _07614_ (
    .a(g35),
    .b(_02529_),
    .c(_02530_),
    .y(_02531_)
  );
  al_aoi21ftf _07615_ (
    .a(\DFF_651.Q ),
    .b(_00066_),
    .c(_02531_),
    .y(\DFF_1066.D )
  );
  al_mux2l _07616_ (
    .a(\DFF_755.Q ),
    .b(\DFF_433.Q ),
    .s(_02341_),
    .y(\DFF_433.D )
  );
  al_and2 _07617_ (
    .a(\DFF_599.Q ),
    .b(g35),
    .y(_02532_)
  );
  al_aoi21ttf _07618_ (
    .a(_02532_),
    .b(_00729_),
    .c(\DFF_1162.Q ),
    .y(\DFF_1404.D )
  );
  al_or3 _07619_ (
    .a(\DFF_937.Q ),
    .b(\DFF_408.Q ),
    .c(\DFF_60.Q ),
    .y(_02533_)
  );
  al_nand3 _07620_ (
    .a(\DFF_1008.Q ),
    .b(\DFF_1275.Q ),
    .c(_02533_),
    .y(_02534_)
  );
  al_and2ft _07621_ (
    .a(\DFF_990.Q ),
    .b(g35),
    .y(_02535_)
  );
  al_aoi21ftf _07622_ (
    .a(\DFF_740.Q ),
    .b(_02534_),
    .c(_02535_),
    .y(_02536_)
  );
  al_ao21ftf _07623_ (
    .a(_02534_),
    .b(\DFF_740.Q ),
    .c(_02536_),
    .y(_02537_)
  );
  al_ao21ftf _07624_ (
    .a(g35),
    .b(\DFF_1008.Q ),
    .c(_02537_),
    .y(\DFF_740.D )
  );
  al_nand3 _07625_ (
    .a(\DFF_1342.Q ),
    .b(g35),
    .c(_00365_),
    .y(_02538_)
  );
  al_or2 _07626_ (
    .a(\DFF_1409.Q ),
    .b(g35),
    .y(_02539_)
  );
  al_or3ftt _07627_ (
    .a(g35),
    .b(\DFF_1342.Q ),
    .c(_00365_),
    .y(_02540_)
  );
  al_and3 _07628_ (
    .a(_02539_),
    .b(_02538_),
    .c(_02540_),
    .y(\DFF_1342.D )
  );
  al_nand3ftt _07629_ (
    .a(_00497_),
    .b(_01772_),
    .c(_00499_),
    .y(_02541_)
  );
  al_ao21ftt _07630_ (
    .a(_00497_),
    .b(_01772_),
    .c(\DFF_1007.Q ),
    .y(_02542_)
  );
  al_nand3 _07631_ (
    .a(g35),
    .b(_02541_),
    .c(_02542_),
    .y(_02543_)
  );
  al_ao21ftf _07632_ (
    .a(g35),
    .b(\DFF_172.Q ),
    .c(_02543_),
    .y(\DFF_1007.D )
  );
  al_nand3 _07633_ (
    .a(_00499_),
    .b(_00508_),
    .c(_01787_),
    .y(_02544_)
  );
  al_ao21 _07634_ (
    .a(_00508_),
    .b(_01787_),
    .c(\DFF_1120.Q ),
    .y(_02545_)
  );
  al_nand3 _07635_ (
    .a(g35),
    .b(_02545_),
    .c(_02544_),
    .y(_02546_)
  );
  al_ao21ftf _07636_ (
    .a(g35),
    .b(\DFF_1294.Q ),
    .c(_02546_),
    .y(\DFF_1120.D )
  );
  al_nand3 _07637_ (
    .a(\DFF_1148.Q ),
    .b(\DFF_60.Q ),
    .c(\DFF_717.Q ),
    .y(_02547_)
  );
  al_aoi21 _07638_ (
    .a(\DFF_1131.Q ),
    .b(_02547_),
    .c(_00066_),
    .y(_02548_)
  );
  al_ao21ftf _07639_ (
    .a(_02547_),
    .b(\DFF_67.Q ),
    .c(_02548_),
    .y(_02549_)
  );
  al_aoi21ftf _07640_ (
    .a(\DFF_1407.Q ),
    .b(_00066_),
    .c(_02549_),
    .y(\DFF_1131.D )
  );
  al_mux2l _07641_ (
    .a(\DFF_69.Q ),
    .b(\DFF_1178.Q ),
    .s(g35),
    .y(\DFF_69.D )
  );
  al_mux2l _07642_ (
    .a(\DFF_1319.Q ),
    .b(\DFF_1270.Q ),
    .s(g35),
    .y(\DFF_1319.D )
  );
  al_and2ft _07643_ (
    .a(g35),
    .b(\DFF_1090.Q ),
    .y(_02550_)
  );
  al_and2 _07644_ (
    .a(\DFF_1090.Q ),
    .b(_01234_),
    .y(_02551_)
  );
  al_ao21ftt _07645_ (
    .a(_00189_),
    .b(_01183_),
    .c(_02551_),
    .y(_02552_)
  );
  al_nor2 _07646_ (
    .a(_00066_),
    .b(_02430_),
    .y(_02553_)
  );
  al_ao21 _07647_ (
    .a(_02553_),
    .b(_02552_),
    .c(_02550_),
    .y(\DFF_874.D )
  );
  al_oai21ftf _07648_ (
    .a(\DFF_830.Q ),
    .b(\DFF_810.Q ),
    .c(\DFF_1298.Q ),
    .y(_02554_)
  );
  al_nand3ftt _07649_ (
    .a(\DFF_1414.Q ),
    .b(g35),
    .c(_02554_),
    .y(_02555_)
  );
  al_ao21ftf _07650_ (
    .a(g35),
    .b(\DFF_810.Q ),
    .c(_02555_),
    .y(\DFF_1298.D )
  );
  al_aoi21ftf _07651_ (
    .a(_00829_),
    .b(_00828_),
    .c(_00830_),
    .y(_02556_)
  );
  al_mux2h _07652_ (
    .a(\DFF_1343.Q ),
    .b(_02556_),
    .s(g35),
    .y(\DFF_1153.D )
  );
  al_ao21ftt _07653_ (
    .a(\DFF_487.Q ),
    .b(_00550_),
    .c(\DFF_1104.Q ),
    .y(_02557_)
  );
  al_and2ft _07654_ (
    .a(g35),
    .b(\DFF_534.Q ),
    .y(_02558_)
  );
  al_ao21 _07655_ (
    .a(_00552_),
    .b(_02557_),
    .c(_02558_),
    .y(\DFF_1104.D )
  );
  al_nand2 _07656_ (
    .a(\DFF_901.Q ),
    .b(\DFF_1275.Q ),
    .y(_02559_)
  );
  al_aoi21 _07657_ (
    .a(_02559_),
    .b(_01472_),
    .c(_00534_),
    .y(_02560_)
  );
  al_mux2h _07658_ (
    .a(\DFF_1117.Q ),
    .b(_02560_),
    .s(g35),
    .y(\DFF_901.D )
  );
  al_or2 _07659_ (
    .a(_00066_),
    .b(_01914_),
    .y(_02561_)
  );
  al_mux2l _07660_ (
    .a(\DFF_795.Q ),
    .b(\DFF_637.Q ),
    .s(_02561_),
    .y(\DFF_637.D )
  );
  al_oai21ftt _07661_ (
    .a(g44),
    .b(\DFF_1178.Q ),
    .c(g35),
    .y(_02562_)
  );
  al_ao21ftf _07662_ (
    .a(g35),
    .b(\DFF_881.Q ),
    .c(_02562_),
    .y(\DFF_1178.D )
  );
  al_oai21 _07663_ (
    .a(\DFF_242.Q ),
    .b(\DFF_858.Q ),
    .c(g35),
    .y(_02563_)
  );
  al_ao21ftf _07664_ (
    .a(g35),
    .b(\DFF_749.Q ),
    .c(_02563_),
    .y(\DFF_242.D )
  );
  al_nor2 _07665_ (
    .a(\DFF_191.Q ),
    .b(g35),
    .y(_02564_)
  );
  al_and2 _07666_ (
    .a(_01335_),
    .b(_01337_),
    .y(_02565_)
  );
  al_mux2l _07667_ (
    .a(\DFF_539.Q ),
    .b(\DFF_1392.Q ),
    .s(\DFF_191.Q ),
    .y(_02566_)
  );
  al_nand3ftt _07668_ (
    .a(_02566_),
    .b(\DFF_557.Q ),
    .c(_02565_),
    .y(_02567_)
  );
  al_aoi21ftf _07669_ (
    .a(\DFF_557.Q ),
    .b(_02566_),
    .c(g35),
    .y(_02568_)
  );
  al_aoi21 _07670_ (
    .a(_02568_),
    .b(_02567_),
    .c(_02564_),
    .y(\DFF_557.D )
  );
  al_ao21 _07671_ (
    .a(\DFF_47.Q ),
    .b(\DFF_1145.Q ),
    .c(\DFF_353.Q ),
    .y(_02569_)
  );
  al_and3ftt _07672_ (
    .a(\DFF_447.Q ),
    .b(\DFF_591.Q ),
    .c(_01348_),
    .y(_02570_)
  );
  al_nand3 _07673_ (
    .a(\DFF_1145.Q ),
    .b(_02569_),
    .c(_02570_),
    .y(_02571_)
  );
  al_ao21 _07674_ (
    .a(_02569_),
    .b(_02570_),
    .c(\DFF_1145.Q ),
    .y(_02572_)
  );
  al_oa21ftt _07675_ (
    .a(\DFF_866.Q ),
    .b(\DFF_900.Q ),
    .c(g35),
    .y(_02573_)
  );
  al_inv _07676_ (
    .a(_02573_),
    .y(_02574_)
  );
  al_ao21 _07677_ (
    .a(_02571_),
    .b(_02572_),
    .c(_02574_),
    .y(_02575_)
  );
  al_aoi21ftf _07678_ (
    .a(\DFF_353.Q ),
    .b(_00066_),
    .c(_02575_),
    .y(\DFF_1145.D )
  );
  al_and2ft _07679_ (
    .a(\DFF_1419.Q ),
    .b(_00827_),
    .y(_02576_)
  );
  al_mux2l _07680_ (
    .a(\DFF_1419.Q ),
    .b(_02576_),
    .s(_01206_),
    .y(_02577_)
  );
  al_mux2h _07681_ (
    .a(\DFF_316.Q ),
    .b(_02577_),
    .s(g35),
    .y(\DFF_1419.D )
  );
  al_ao21 _07682_ (
    .a(\DFF_447.Q ),
    .b(_01348_),
    .c(_01879_),
    .y(_02578_)
  );
  al_ao21ttf _07683_ (
    .a(\DFF_591.Q ),
    .b(_01350_),
    .c(_01348_),
    .y(_02579_)
  );
  al_aoi21 _07684_ (
    .a(_02579_),
    .b(_02578_),
    .c(_00066_),
    .y(\DFF_786.D )
  );
  al_oa21 _07685_ (
    .a(\DFF_349.Q ),
    .b(\DFF_1245.Q ),
    .c(g35),
    .y(\DFF_1245.D )
  );
  al_and2ft _07686_ (
    .a(g35),
    .b(\DFF_518.Q ),
    .y(_02580_)
  );
  al_inv _07687_ (
    .a(\DFF_518.Q ),
    .y(_02581_)
  );
  al_inv _07688_ (
    .a(\DFF_665.Q ),
    .y(_02582_)
  );
  al_nand2ft _07689_ (
    .a(\DFF_1132.Q ),
    .b(_01339_),
    .y(_02583_)
  );
  al_or3fft _07690_ (
    .a(_02582_),
    .b(_02581_),
    .c(_02583_),
    .y(_02584_)
  );
  al_aoi21ftf _07691_ (
    .a(_02581_),
    .b(_01870_),
    .c(_02584_),
    .y(_02585_)
  );
  al_ao21ftf _07692_ (
    .a(_01872_),
    .b(_01335_),
    .c(_02585_),
    .y(_02586_)
  );
  al_oa21ftf _07693_ (
    .a(\DFF_823.Q ),
    .b(_02585_),
    .c(_00066_),
    .y(_02587_)
  );
  al_ao21 _07694_ (
    .a(_02586_),
    .b(_02587_),
    .c(_02580_),
    .y(\DFF_823.D )
  );
  al_or2 _07695_ (
    .a(_00066_),
    .b(_02040_),
    .y(_02588_)
  );
  al_and3fft _07696_ (
    .a(_00066_),
    .b(_01363_),
    .c(_02039_),
    .y(_02589_)
  );
  al_aoi21 _07697_ (
    .a(_01361_),
    .b(_02588_),
    .c(_02589_),
    .y(\DFF_1236.D )
  );
  al_mux2l _07698_ (
    .a(\DFF_541.Q ),
    .b(\DFF_430.Q ),
    .s(_00478_),
    .y(_02590_)
  );
  al_mux2h _07699_ (
    .a(\DFF_427.Q ),
    .b(_02590_),
    .s(g35),
    .y(\DFF_430.D )
  );
  al_inv _07700_ (
    .a(\DFF_472.Q ),
    .y(_02591_)
  );
  al_and2 _07701_ (
    .a(\DFF_1413.Q ),
    .b(_01150_),
    .y(_02592_)
  );
  al_nand3 _07702_ (
    .a(\DFF_1181.Q ),
    .b(_00604_),
    .c(_00323_),
    .y(_02593_)
  );
  al_oa21ftf _07703_ (
    .a(\DFF_671.Q ),
    .b(_01150_),
    .c(_00066_),
    .y(_02594_)
  );
  al_ao21ttf _07704_ (
    .a(_02592_),
    .b(_02593_),
    .c(_02594_),
    .y(_02595_)
  );
  al_aoi21ftf _07705_ (
    .a(g35),
    .b(_02591_),
    .c(_02595_),
    .y(\DFF_671.D )
  );
  al_mux2l _07706_ (
    .a(\DFF_1125.Q ),
    .b(\DFF_1245.Q ),
    .s(g35),
    .y(\DFF_1125.D )
  );
  al_or2 _07707_ (
    .a(_01755_),
    .b(_01150_),
    .y(_02596_)
  );
  al_inv _07708_ (
    .a(\DFF_996.Q ),
    .y(_02597_)
  );
  al_and2 _07709_ (
    .a(_02597_),
    .b(_01150_),
    .y(_02598_)
  );
  al_nand3 _07710_ (
    .a(_01151_),
    .b(_02598_),
    .c(_02593_),
    .y(_02599_)
  );
  al_aoi21 _07711_ (
    .a(_02596_),
    .b(_02599_),
    .c(_00066_),
    .y(\DFF_1413.D )
  );
  al_oai21ftf _07712_ (
    .a(\DFF_86.Q ),
    .b(\DFF_553.Q ),
    .c(\DFF_1048.Q ),
    .y(_02600_)
  );
  al_nand3ftt _07713_ (
    .a(\DFF_1316.Q ),
    .b(g35),
    .c(_02600_),
    .y(_02601_)
  );
  al_ao21ftf _07714_ (
    .a(g35),
    .b(\DFF_553.Q ),
    .c(_02601_),
    .y(\DFF_1048.D )
  );
  al_aoi21 _07715_ (
    .a(\DFF_47.Q ),
    .b(_02571_),
    .c(_02574_),
    .y(_02602_)
  );
  al_oai21 _07716_ (
    .a(\DFF_47.Q ),
    .b(_02571_),
    .c(_02602_),
    .y(_02603_)
  );
  al_aoi21ftf _07717_ (
    .a(\DFF_1145.Q ),
    .b(_00066_),
    .c(_02603_),
    .y(\DFF_47.D )
  );
  al_nand3 _07718_ (
    .a(_00499_),
    .b(_00706_),
    .c(_02114_),
    .y(_02604_)
  );
  al_ao21 _07719_ (
    .a(_00706_),
    .b(_02114_),
    .c(\DFF_1401.Q ),
    .y(_02605_)
  );
  al_nand3 _07720_ (
    .a(g35),
    .b(_02605_),
    .c(_02604_),
    .y(_02606_)
  );
  al_ao21ftf _07721_ (
    .a(g35),
    .b(\DFF_1197.Q ),
    .c(_02606_),
    .y(\DFF_1401.D )
  );
  al_nand3 _07722_ (
    .a(_01884_),
    .b(\DFF_500.Q ),
    .c(_01889_),
    .y(_02607_)
  );
  al_aoi21ftf _07723_ (
    .a(\DFF_16.Q ),
    .b(_02607_),
    .c(g35),
    .y(_02608_)
  );
  al_oai21 _07724_ (
    .a(_01892_),
    .b(_02607_),
    .c(_02608_),
    .y(_02609_)
  );
  al_ao21ftf _07725_ (
    .a(g35),
    .b(\DFF_41.Q ),
    .c(_02609_),
    .y(\DFF_16.D )
  );
  al_or2ft _07726_ (
    .a(\DFF_395.Q ),
    .b(_00971_),
    .y(_02610_)
  );
  al_ao21ttf _07727_ (
    .a(_02610_),
    .b(_00976_),
    .c(_00974_),
    .y(_02611_)
  );
  al_or3fft _07728_ (
    .a(\DFF_1115.Q ),
    .b(_02611_),
    .c(_02045_),
    .y(_02612_)
  );
  al_oai21ftf _07729_ (
    .a(\DFF_1115.Q ),
    .b(_02045_),
    .c(_02611_),
    .y(_02613_)
  );
  al_nand3 _07730_ (
    .a(g35),
    .b(_02612_),
    .c(_02613_),
    .y(_02614_)
  );
  al_aoi21ftf _07731_ (
    .a(\DFF_886.Q ),
    .b(_00066_),
    .c(_02614_),
    .y(\DFF_1115.D )
  );
  al_oa21ftt _07732_ (
    .a(g35),
    .b(\DFF_701.Q ),
    .c(\DFF_939.Q ),
    .y(_02615_)
  );
  al_aoi21ttf _07733_ (
    .a(\DFF_523.Q ),
    .b(g35),
    .c(_02615_),
    .y(_02616_)
  );
  al_or3fft _07734_ (
    .a(\DFF_523.Q ),
    .b(g35),
    .c(_02615_),
    .y(_02617_)
  );
  al_nand2ft _07735_ (
    .a(_02616_),
    .b(_02617_),
    .y(\DFF_523.D )
  );
  al_nand3fft _07736_ (
    .a(\DFF_20.Q ),
    .b(\DFF_916.Q ),
    .c(\DFF_104.Q ),
    .y(_02618_)
  );
  al_aoi21ftf _07737_ (
    .a(\DFF_337.Q ),
    .b(_02618_),
    .c(g35),
    .y(_02619_)
  );
  al_ao21ftf _07738_ (
    .a(_02618_),
    .b(_00499_),
    .c(_02619_),
    .y(_02620_)
  );
  al_ao21ftf _07739_ (
    .a(g35),
    .b(\DFF_1366.Q ),
    .c(_02620_),
    .y(\DFF_337.D )
  );
  al_oa21ftt _07740_ (
    .a(g35),
    .b(\DFF_466.Q ),
    .c(\DFF_1333.Q ),
    .y(\DFF_572.D )
  );
  al_nand3 _07741_ (
    .a(_00320_),
    .b(_00526_),
    .c(_00530_),
    .y(_02621_)
  );
  al_ao21 _07742_ (
    .a(_00320_),
    .b(_00526_),
    .c(\DFF_469.Q ),
    .y(_02622_)
  );
  al_nand3 _07743_ (
    .a(g35),
    .b(_02622_),
    .c(_02621_),
    .y(_02623_)
  );
  al_ao21ftf _07744_ (
    .a(g35),
    .b(\DFF_1247.Q ),
    .c(_02623_),
    .y(\DFF_469.D )
  );
  al_and2 _07745_ (
    .a(\DFF_20.Q ),
    .b(\DFF_916.Q ),
    .y(_02624_)
  );
  al_and2 _07746_ (
    .a(\DFF_925.Q ),
    .b(\DFF_653.Q ),
    .y(_02625_)
  );
  al_nand3 _07747_ (
    .a(_00499_),
    .b(_02624_),
    .c(_02625_),
    .y(_02626_)
  );
  al_ao21 _07748_ (
    .a(_02624_),
    .b(_02625_),
    .c(\DFF_298.Q ),
    .y(_02627_)
  );
  al_nand3 _07749_ (
    .a(g35),
    .b(_02626_),
    .c(_02627_),
    .y(_02628_)
  );
  al_ao21ftf _07750_ (
    .a(g35),
    .b(\DFF_82.Q ),
    .c(_02628_),
    .y(\DFF_298.D )
  );
  al_or2 _07751_ (
    .a(\DFF_343.Q ),
    .b(_01147_),
    .y(_02629_)
  );
  al_ao21ttf _07752_ (
    .a(_02629_),
    .b(_01152_),
    .c(_01150_),
    .y(_02630_)
  );
  al_nand3 _07753_ (
    .a(\DFF_1376.Q ),
    .b(_01195_),
    .c(_02630_),
    .y(_02631_)
  );
  al_ao21 _07754_ (
    .a(\DFF_1376.Q ),
    .b(_01195_),
    .c(_02630_),
    .y(_02632_)
  );
  al_nand3 _07755_ (
    .a(g35),
    .b(_02631_),
    .c(_02632_),
    .y(_02633_)
  );
  al_aoi21ftf _07756_ (
    .a(\DFF_996.Q ),
    .b(_00066_),
    .c(_02633_),
    .y(\DFF_1376.D )
  );
  al_nand3 _07757_ (
    .a(\DFF_755.Q ),
    .b(g35),
    .c(_00373_),
    .y(_02634_)
  );
  al_or3ftt _07758_ (
    .a(g35),
    .b(\DFF_755.Q ),
    .c(_00373_),
    .y(_02635_)
  );
  al_or2 _07759_ (
    .a(\DFF_987.Q ),
    .b(g35),
    .y(_02636_)
  );
  al_and3 _07760_ (
    .a(_02636_),
    .b(_02634_),
    .c(_02635_),
    .y(\DFF_755.D )
  );
  al_mux2l _07761_ (
    .a(\DFF_374.Q ),
    .b(\DFF_1050.Q ),
    .s(_02455_),
    .y(\DFF_1050.D )
  );
  al_nor2 _07762_ (
    .a(\DFF_1141.Q ),
    .b(g35),
    .y(_02637_)
  );
  al_and2 _07763_ (
    .a(_00322_),
    .b(_00319_),
    .y(_02638_)
  );
  al_nand3 _07764_ (
    .a(\DFF_1181.Q ),
    .b(_00604_),
    .c(_02638_),
    .y(_02639_)
  );
  al_nand3 _07765_ (
    .a(\DFF_1141.Q ),
    .b(_01282_),
    .c(_02639_),
    .y(_02640_)
  );
  al_oa21ftf _07766_ (
    .a(\DFF_1047.Q ),
    .b(_01282_),
    .c(_00066_),
    .y(_02641_)
  );
  al_aoi21 _07767_ (
    .a(_02641_),
    .b(_02640_),
    .c(_02637_),
    .y(\DFF_1047.D )
  );
  al_nor2 _07768_ (
    .a(\DFF_793.Q ),
    .b(g35),
    .y(_02642_)
  );
  al_and3 _07769_ (
    .a(_00604_),
    .b(_00563_),
    .c(_00440_),
    .y(_02643_)
  );
  al_nand3ftt _07770_ (
    .a(\DFF_793.Q ),
    .b(\DFF_148.Q ),
    .c(\DFF_379.Q ),
    .y(_02644_)
  );
  al_oai21ftf _07771_ (
    .a(\DFF_148.Q ),
    .b(\DFF_793.Q ),
    .c(\DFF_379.Q ),
    .y(_02645_)
  );
  al_nand3 _07772_ (
    .a(_02644_),
    .b(_02645_),
    .c(_02643_),
    .y(_02646_)
  );
  al_oa21ftf _07773_ (
    .a(\DFF_1028.Q ),
    .b(_02643_),
    .c(_00066_),
    .y(_02647_)
  );
  al_aoi21 _07774_ (
    .a(_02646_),
    .b(_02647_),
    .c(_02642_),
    .y(\DFF_1028.D )
  );
  al_nand3fft _07775_ (
    .a(\DFF_48.Q ),
    .b(\DFF_760.Q ),
    .c(g35),
    .y(_02648_)
  );
  al_oa21 _07776_ (
    .a(g35),
    .b(\DFF_753.Q ),
    .c(_02648_),
    .y(\DFF_1329.D )
  );
  al_and2 _07777_ (
    .a(\DFF_1010.Q ),
    .b(_00526_),
    .y(_02649_)
  );
  al_nand3 _07778_ (
    .a(\DFF_1181.Q ),
    .b(_00604_),
    .c(_01377_),
    .y(_02650_)
  );
  al_oa21ftf _07779_ (
    .a(\DFF_1233.Q ),
    .b(_00526_),
    .c(_00066_),
    .y(_02651_)
  );
  al_ao21ttf _07780_ (
    .a(_02649_),
    .b(_02650_),
    .c(_02651_),
    .y(_02652_)
  );
  al_aoi21ftf _07781_ (
    .a(\DFF_1010.Q ),
    .b(_00066_),
    .c(_02652_),
    .y(\DFF_1233.D )
  );
  al_and2ft _07782_ (
    .a(g35),
    .b(\DFF_1240.Q ),
    .y(_02653_)
  );
  al_inv _07783_ (
    .a(\DFF_681.Q ),
    .y(_02654_)
  );
  al_aoi21ttf _07784_ (
    .a(_00577_),
    .b(_00425_),
    .c(_01394_),
    .y(_02655_)
  );
  al_ao21ftf _07785_ (
    .a(_01396_),
    .b(_02654_),
    .c(_02655_),
    .y(_02656_)
  );
  al_inv _07786_ (
    .a(\DFF_387.Q ),
    .y(_02657_)
  );
  al_oa21ftf _07787_ (
    .a(_02657_),
    .b(_01394_),
    .c(_00066_),
    .y(_02658_)
  );
  al_ao21 _07788_ (
    .a(_02658_),
    .b(_02656_),
    .c(_02653_),
    .y(\DFF_387.D )
  );
  al_and3 _07789_ (
    .a(\DFF_551.Q ),
    .b(_01832_),
    .c(_01815_),
    .y(_02659_)
  );
  al_nand3 _07790_ (
    .a(\DFF_351.Q ),
    .b(\DFF_508.Q ),
    .c(_02659_),
    .y(_02660_)
  );
  al_aoi21 _07791_ (
    .a(\DFF_201.Q ),
    .b(_02660_),
    .c(_01831_),
    .y(_02661_)
  );
  al_oai21 _07792_ (
    .a(\DFF_201.Q ),
    .b(_02660_),
    .c(_02661_),
    .y(_02662_)
  );
  al_aoi21ftf _07793_ (
    .a(\DFF_508.Q ),
    .b(_00066_),
    .c(_02662_),
    .y(\DFF_201.D )
  );
  al_aoi21 _07794_ (
    .a(\DFF_1027.Q ),
    .b(g35),
    .c(\DFF_1043.Q ),
    .y(_02663_)
  );
  al_and2 _07795_ (
    .a(g35),
    .b(\DFF_1043.Q ),
    .y(_02664_)
  );
  al_aoi21 _07796_ (
    .a(\DFF_1027.Q ),
    .b(_02664_),
    .c(_02663_),
    .y(\DFF_858.D )
  );
  al_and2ft _07797_ (
    .a(\DFF_519.Q ),
    .b(\DFF_385.Q ),
    .y(_02665_)
  );
  al_nand3 _07798_ (
    .a(_00499_),
    .b(_01467_),
    .c(_02665_),
    .y(_02666_)
  );
  al_ao21 _07799_ (
    .a(_02665_),
    .b(_01467_),
    .c(\DFF_1255.Q ),
    .y(_02667_)
  );
  al_nand3 _07800_ (
    .a(g35),
    .b(_02667_),
    .c(_02666_),
    .y(_02668_)
  );
  al_ao21ftf _07801_ (
    .a(g35),
    .b(\DFF_815.Q ),
    .c(_02668_),
    .y(\DFF_1255.D )
  );
  al_and2 _07802_ (
    .a(g35),
    .b(_01014_),
    .y(_02669_)
  );
  al_and3ftt _07803_ (
    .a(\DFF_120.Q ),
    .b(_01028_),
    .c(_02669_),
    .y(\DFF_120.D )
  );
  al_nand3fft _07804_ (
    .a(\DFF_350.Q ),
    .b(g73),
    .c(g72),
    .y(_02670_)
  );
  al_mux2l _07805_ (
    .a(_02670_),
    .b(\DFF_816.Q ),
    .s(_01208_),
    .y(\DFF_1330.D )
  );
  al_oa21ttf _07806_ (
    .a(g35),
    .b(\DFF_1384.Q ),
    .c(_02664_),
    .y(\DFF_1027.D )
  );
  al_nor2 _07807_ (
    .a(\DFF_1299.Q ),
    .b(g35),
    .y(_02671_)
  );
  al_nand3fft _07808_ (
    .a(\DFF_853.Q ),
    .b(_00410_),
    .c(_00998_),
    .y(_02672_)
  );
  al_oai21ftf _07809_ (
    .a(g90),
    .b(\DFF_1125.Q ),
    .c(\DFF_115.Q ),
    .y(_02673_)
  );
  al_nand2ft _07810_ (
    .a(\DFF_1379.Q ),
    .b(\DFF_115.Q ),
    .y(_02674_)
  );
  al_nand3ftt _07811_ (
    .a(\DFF_1084.Q ),
    .b(_02674_),
    .c(_02673_),
    .y(_02675_)
  );
  al_nand2ft _07812_ (
    .a(\DFF_1415.Q ),
    .b(\DFF_1084.Q ),
    .y(_02676_)
  );
  al_ao21 _07813_ (
    .a(_02676_),
    .b(_00605_),
    .c(\DFF_115.Q ),
    .y(_02677_)
  );
  al_nand3ftt _07814_ (
    .a(\DFF_853.Q ),
    .b(_02675_),
    .c(_02677_),
    .y(_02678_)
  );
  al_nand2 _07815_ (
    .a(g35),
    .b(_00608_),
    .y(_02679_)
  );
  al_aoi21 _07816_ (
    .a(_00410_),
    .b(_02678_),
    .c(_02679_),
    .y(_02680_)
  );
  al_aoi21 _07817_ (
    .a(_02680_),
    .b(_02672_),
    .c(_02671_),
    .y(\DFF_26.D )
  );
  al_mux2h _07818_ (
    .a(\DFF_1113.Q ),
    .b(_01039_),
    .s(g35),
    .y(\DFF_975.D )
  );
  al_mux2l _07819_ (
    .a(\DFF_339.Q ),
    .b(\DFF_828.Q ),
    .s(g35),
    .y(\DFF_343.D )
  );
  al_mux2h _07820_ (
    .a(\DFF_1238.Q ),
    .b(_01337_),
    .s(g35),
    .y(\DFF_787.D )
  );
  al_and2ft _07821_ (
    .a(\DFF_271.Q ),
    .b(\DFF_522.Q ),
    .y(_02681_)
  );
  al_and2 _07822_ (
    .a(\DFF_803.Q ),
    .b(\DFF_35.Q ),
    .y(_02682_)
  );
  al_nand3 _07823_ (
    .a(_00499_),
    .b(_02681_),
    .c(_02682_),
    .y(_02683_)
  );
  al_ao21 _07824_ (
    .a(_02681_),
    .b(_02682_),
    .c(\DFF_1410.Q ),
    .y(_02684_)
  );
  al_nand3 _07825_ (
    .a(g35),
    .b(_02684_),
    .c(_02683_),
    .y(_02685_)
  );
  al_ao21ftf _07826_ (
    .a(g35),
    .b(\DFF_225.Q ),
    .c(_02685_),
    .y(\DFF_1410.D )
  );
  al_nand2ft _07827_ (
    .a(\DFF_111.Q ),
    .b(\DFF_759.Q ),
    .y(_02686_)
  );
  al_and3fft _07828_ (
    .a(_02686_),
    .b(_01131_),
    .c(_01125_),
    .y(_02687_)
  );
  al_ao21ftt _07829_ (
    .a(_02686_),
    .b(_01125_),
    .c(\DFF_968.Q ),
    .y(_02688_)
  );
  al_or3fft _07830_ (
    .a(g35),
    .b(_02688_),
    .c(_02687_),
    .y(_02689_)
  );
  al_ao21ftf _07831_ (
    .a(g35),
    .b(\DFF_504.Q ),
    .c(_02689_),
    .y(\DFF_968.D )
  );
  al_ao21 _07832_ (
    .a(\DFF_351.Q ),
    .b(_02659_),
    .c(\DFF_508.Q ),
    .y(_02690_)
  );
  al_ao21 _07833_ (
    .a(_02660_),
    .b(_02690_),
    .c(_01831_),
    .y(_02691_)
  );
  al_aoi21ftf _07834_ (
    .a(\DFF_351.Q ),
    .b(_00066_),
    .c(_02691_),
    .y(\DFF_508.D )
  );
  al_or2ft _07835_ (
    .a(\DFF_1260.Q ),
    .b(_00361_),
    .y(_02692_)
  );
  al_inv _07836_ (
    .a(\DFF_1383.Q ),
    .y(_02693_)
  );
  al_or2ft _07837_ (
    .a(g35),
    .b(_00361_),
    .y(_02694_)
  );
  al_ao21ftf _07838_ (
    .a(_02693_),
    .b(_00987_),
    .c(_02694_),
    .y(_02695_)
  );
  al_and3ftt _07839_ (
    .a(_00987_),
    .b(_02693_),
    .c(_02694_),
    .y(_02696_)
  );
  al_aoi21 _07840_ (
    .a(_02692_),
    .b(_02695_),
    .c(_02696_),
    .y(\DFF_1260.D )
  );
  al_and3ftt _07841_ (
    .a(\DFF_1037.Q ),
    .b(\DFF_173.Q ),
    .c(\DFF_552.Q ),
    .y(_02697_)
  );
  al_and3ftt _07842_ (
    .a(\DFF_1375.Q ),
    .b(\DFF_1137.Q ),
    .c(\DFF_1037.Q ),
    .y(_02698_)
  );
  al_and2ft _07843_ (
    .a(\DFF_1037.Q ),
    .b(\DFF_1375.Q ),
    .y(_02699_)
  );
  al_ao21 _07844_ (
    .a(\DFF_16.Q ),
    .b(_02699_),
    .c(_02698_),
    .y(_02700_)
  );
  al_nand3 _07845_ (
    .a(\DFF_1375.Q ),
    .b(\DFF_1258.Q ),
    .c(\DFF_552.Q ),
    .y(_02701_)
  );
  al_and3fft _07846_ (
    .a(\DFF_1375.Q ),
    .b(\DFF_552.Q ),
    .c(\DFF_306.Q ),
    .y(_02702_)
  );
  al_and3ftt _07847_ (
    .a(\DFF_552.Q ),
    .b(\DFF_1037.Q ),
    .c(\DFF_41.Q ),
    .y(_02703_)
  );
  al_and3fft _07848_ (
    .a(_02703_),
    .b(_02702_),
    .c(_02701_),
    .y(_02704_)
  );
  al_nand3fft _07849_ (
    .a(_02697_),
    .b(_02700_),
    .c(_02704_),
    .y(_02705_)
  );
  al_mux2l _07850_ (
    .a(_02705_),
    .b(\DFF_1167.Q ),
    .s(_00546_),
    .y(_02706_)
  );
  al_mux2h _07851_ (
    .a(\DFF_1375.Q ),
    .b(_02706_),
    .s(g35),
    .y(\DFF_1167.D )
  );
  al_and2ft _07852_ (
    .a(\DFF_776.Q ),
    .b(\DFF_784.Q ),
    .y(_02707_)
  );
  al_nand3 _07853_ (
    .a(_00499_),
    .b(_00597_),
    .c(_02707_),
    .y(_02708_)
  );
  al_ao21 _07854_ (
    .a(_00597_),
    .b(_02707_),
    .c(\DFF_1128.Q ),
    .y(_02709_)
  );
  al_nand3 _07855_ (
    .a(g35),
    .b(_02709_),
    .c(_02708_),
    .y(_02710_)
  );
  al_ao21ftf _07856_ (
    .a(g35),
    .b(\DFF_1350.Q ),
    .c(_02710_),
    .y(\DFF_1128.D )
  );
  al_ao21ftf _07857_ (
    .a(g113),
    .b(_00342_),
    .c(\DFF_1036.Q ),
    .y(_02711_)
  );
  al_nand3ftt _07858_ (
    .a(_01559_),
    .b(_02711_),
    .c(_01272_),
    .y(_02712_)
  );
  al_ao21ftf _07859_ (
    .a(_01272_),
    .b(\DFF_1.Q ),
    .c(_02712_),
    .y(_02713_)
  );
  al_mux2h _07860_ (
    .a(\DFF_1288.Q ),
    .b(_02713_),
    .s(g35),
    .y(\DFF_1.D )
  );
  al_and2ft _07861_ (
    .a(\DFF_339.Q ),
    .b(g35),
    .y(_02714_)
  );
  al_oai21ftf _07862_ (
    .a(\DFF_339.Q ),
    .b(\DFF_261.Q ),
    .c(\DFF_1133.Q ),
    .y(_02715_)
  );
  al_ao21 _07863_ (
    .a(\DFF_1207.Q ),
    .b(_02715_),
    .c(_00066_),
    .y(_02716_)
  );
  al_ao21ftf _07864_ (
    .a(_02714_),
    .b(\DFF_1133.Q ),
    .c(_02716_),
    .y(\DFF_24.D )
  );
  al_mux2l _07865_ (
    .a(g116),
    .b(g114),
    .s(\DFF_767.Q ),
    .y(_02717_)
  );
  al_mux2h _07866_ (
    .a(\DFF_116.Q ),
    .b(_02717_),
    .s(g35),
    .y(\DFF_282.D )
  );
  al_ao21ttf _07867_ (
    .a(\DFF_953.Q ),
    .b(g35),
    .c(\DFF_896.Q ),
    .y(_02718_)
  );
  al_or3fft _07868_ (
    .a(\DFF_953.Q ),
    .b(_01175_),
    .c(_00953_),
    .y(_02719_)
  );
  al_ao21ftf _07869_ (
    .a(_02718_),
    .b(_02375_),
    .c(_02719_),
    .y(\DFF_953.D )
  );
  al_mux2l _07870_ (
    .a(\DFF_1275.Q ),
    .b(\DFF_481.Q ),
    .s(g35),
    .y(\DFF_395.D )
  );
  al_ao21ftt _07871_ (
    .a(_01460_),
    .b(\DFF_303.Q ),
    .c(_01462_),
    .y(_02720_)
  );
  al_or3fft _07872_ (
    .a(g35),
    .b(_02720_),
    .c(_01593_),
    .y(_02721_)
  );
  al_ao21ftf _07873_ (
    .a(g35),
    .b(\DFF_1241.Q ),
    .c(_02721_),
    .y(\DFF_303.D )
  );
  al_and2ft _07874_ (
    .a(\DFF_463.Q ),
    .b(\DFF_14.Q ),
    .y(_02722_)
  );
  al_nand2ft _07875_ (
    .a(\DFF_14.Q ),
    .b(\DFF_463.Q ),
    .y(_02723_)
  );
  al_nand2ft _07876_ (
    .a(_02722_),
    .b(_02723_),
    .y(_02724_)
  );
  al_mux2l _07877_ (
    .a(\DFF_679.Q ),
    .b(_02724_),
    .s(_01958_),
    .y(_02725_)
  );
  al_mux2h _07878_ (
    .a(\DFF_463.Q ),
    .b(_02725_),
    .s(g35),
    .y(\DFF_679.D )
  );
  al_and2 _07879_ (
    .a(g35),
    .b(_00734_),
    .y(_02726_)
  );
  al_and3ftt _07880_ (
    .a(\DFF_784.Q ),
    .b(_01270_),
    .c(_02726_),
    .y(\DFF_784.D )
  );
  al_ao21 _07881_ (
    .a(_00793_),
    .b(_00766_),
    .c(_00066_),
    .y(_02727_)
  );
  al_mux2l _07882_ (
    .a(\DFF_589.Q ),
    .b(\DFF_341.Q ),
    .s(_02727_),
    .y(\DFF_341.D )
  );
  al_mux2l _07883_ (
    .a(\DFF_39.Q ),
    .b(\DFF_1214.Q ),
    .s(\DFF_1312.Q ),
    .y(_02728_)
  );
  al_aoi21 _07884_ (
    .a(\DFF_536.Q ),
    .b(_02728_),
    .c(\DFF_574.Q ),
    .y(_02729_)
  );
  al_oai21 _07885_ (
    .a(\DFF_536.Q ),
    .b(_02728_),
    .c(_02729_),
    .y(_02730_)
  );
  al_and3ftt _07886_ (
    .a(\DFF_892.Q ),
    .b(\DFF_1199.Q ),
    .c(_00464_),
    .y(_02731_)
  );
  al_ao21ttf _07887_ (
    .a(_02731_),
    .b(_02730_),
    .c(_00766_),
    .y(_02732_)
  );
  al_or2 _07888_ (
    .a(\DFF_574.Q ),
    .b(_00766_),
    .y(_02733_)
  );
  al_and3 _07889_ (
    .a(g35),
    .b(_02732_),
    .c(_02733_),
    .y(\DFF_574.D )
  );
  al_mux2l _07890_ (
    .a(\DFF_840.Q ),
    .b(\DFF_224.Q ),
    .s(\DFF_1347.Q ),
    .y(_02734_)
  );
  al_aoi21 _07891_ (
    .a(\DFF_443.Q ),
    .b(_02734_),
    .c(\DFF_1206.Q ),
    .y(_02735_)
  );
  al_oai21 _07892_ (
    .a(\DFF_443.Q ),
    .b(_02734_),
    .c(_02735_),
    .y(_02736_)
  );
  al_ao21ftf _07893_ (
    .a(_01863_),
    .b(_02736_),
    .c(_02064_),
    .y(_02737_)
  );
  al_or2 _07894_ (
    .a(\DFF_1206.Q ),
    .b(_02064_),
    .y(_02738_)
  );
  al_and3 _07895_ (
    .a(g35),
    .b(_02737_),
    .c(_02738_),
    .y(\DFF_1206.D )
  );
  al_aoi21 _07896_ (
    .a(\DFF_1148.Q ),
    .b(\DFF_60.Q ),
    .c(\DFF_717.Q ),
    .y(_02739_)
  );
  al_ao21ftf _07897_ (
    .a(_00521_),
    .b(\DFF_1159.Q ),
    .c(_00965_),
    .y(_02740_)
  );
  al_and2 _07898_ (
    .a(g35),
    .b(_02740_),
    .y(_02741_)
  );
  al_ao21ftf _07899_ (
    .a(_02739_),
    .b(_02547_),
    .c(_02741_),
    .y(_02742_)
  );
  al_aoi21ftf _07900_ (
    .a(\DFF_1148.Q ),
    .b(_00066_),
    .c(_02742_),
    .y(\DFF_717.D )
  );
  al_nand3 _07901_ (
    .a(_00499_),
    .b(_02114_),
    .c(_02681_),
    .y(_02743_)
  );
  al_ao21 _07902_ (
    .a(_02114_),
    .b(_02681_),
    .c(\DFF_1166.Q ),
    .y(_02744_)
  );
  al_nand3 _07903_ (
    .a(g35),
    .b(_02744_),
    .c(_02743_),
    .y(_02745_)
  );
  al_ao21ftf _07904_ (
    .a(g35),
    .b(\DFF_1386.Q ),
    .c(_02745_),
    .y(\DFF_1166.D )
  );
  al_oai21ftf _07905_ (
    .a(\DFF_119.Q ),
    .b(_01237_),
    .c(_01229_),
    .y(_02746_)
  );
  al_nand3 _07906_ (
    .a(g35),
    .b(_01238_),
    .c(_02746_),
    .y(_02747_)
  );
  al_ao21ftf _07907_ (
    .a(g35),
    .b(\DFF_119.Q ),
    .c(_02747_),
    .y(\DFF_844.D )
  );
  al_nor2 _07908_ (
    .a(\DFF_889.Q ),
    .b(g35),
    .y(_02748_)
  );
  al_and3 _07909_ (
    .a(_00604_),
    .b(_00576_),
    .c(_00449_),
    .y(_02749_)
  );
  al_nand3ftt _07910_ (
    .a(\DFF_889.Q ),
    .b(\DFF_1091.Q ),
    .c(\DFF_379.Q ),
    .y(_02750_)
  );
  al_oai21ftf _07911_ (
    .a(\DFF_1091.Q ),
    .b(\DFF_889.Q ),
    .c(\DFF_379.Q ),
    .y(_02751_)
  );
  al_nand3 _07912_ (
    .a(_02750_),
    .b(_02751_),
    .c(_02749_),
    .y(_02752_)
  );
  al_oa21ftf _07913_ (
    .a(\DFF_462.Q ),
    .b(_02749_),
    .c(_00066_),
    .y(_02753_)
  );
  al_aoi21 _07914_ (
    .a(_02752_),
    .b(_02753_),
    .c(_02748_),
    .y(\DFF_462.D )
  );
  al_nor2 _07915_ (
    .a(\DFF_271.Q ),
    .b(\DFF_522.Q ),
    .y(_02754_)
  );
  al_nand3 _07916_ (
    .a(_00499_),
    .b(_02114_),
    .c(_02754_),
    .y(_02755_)
  );
  al_ao21 _07917_ (
    .a(_02114_),
    .b(_02754_),
    .c(\DFF_1218.Q ),
    .y(_02756_)
  );
  al_nand3 _07918_ (
    .a(g35),
    .b(_02756_),
    .c(_02755_),
    .y(_02757_)
  );
  al_ao21ftf _07919_ (
    .a(g35),
    .b(\DFF_1378.Q ),
    .c(_02757_),
    .y(\DFF_1218.D )
  );
  al_mux2l _07920_ (
    .a(g6749),
    .b(\DFF_383.Q ),
    .s(g35),
    .y(\DFF_911.D )
  );
  al_and2ft _07921_ (
    .a(\DFF_399.Q ),
    .b(\DFF_1131.Q ),
    .y(_02758_)
  );
  al_nand3 _07922_ (
    .a(\DFF_416.Q ),
    .b(g35),
    .c(_02758_),
    .y(_02759_)
  );
  al_aoi21ftf _07923_ (
    .a(\DFF_733.Q ),
    .b(_00066_),
    .c(_02759_),
    .y(\DFF_399.D )
  );
  al_oai21ftf _07924_ (
    .a(\DFF_371.Q ),
    .b(\DFF_168.Q ),
    .c(\DFF_1279.Q ),
    .y(_02760_)
  );
  al_nand3ftt _07925_ (
    .a(\DFF_861.Q ),
    .b(g35),
    .c(_02760_),
    .y(_02761_)
  );
  al_ao21ftf _07926_ (
    .a(g35),
    .b(\DFF_168.Q ),
    .c(_02761_),
    .y(\DFF_1279.D )
  );
  al_aoi21 _07927_ (
    .a(\DFF_869.Q ),
    .b(g35),
    .c(\DFF_636.Q ),
    .y(_02762_)
  );
  al_oa21ftt _07928_ (
    .a(g35),
    .b(\DFF_636.Q ),
    .c(\DFF_869.Q ),
    .y(_02763_)
  );
  al_aoi21 _07929_ (
    .a(g35),
    .b(_02763_),
    .c(_02762_),
    .y(\DFF_869.D )
  );
  al_oai21ftf _07930_ (
    .a(\DFF_861.Q ),
    .b(\DFF_603.Q ),
    .c(\DFF_732.Q ),
    .y(_02764_)
  );
  al_nand3ftt _07931_ (
    .a(\DFF_371.Q ),
    .b(g35),
    .c(_02764_),
    .y(_02765_)
  );
  al_ao21ftf _07932_ (
    .a(g35),
    .b(\DFF_603.Q ),
    .c(_02765_),
    .y(\DFF_732.D )
  );
  al_and3ftt _07933_ (
    .a(\DFF_849.Q ),
    .b(\DFF_894.Q ),
    .c(_00461_),
    .y(_02766_)
  );
  al_ao21 _07934_ (
    .a(_02766_),
    .b(_01222_),
    .c(_00066_),
    .y(_02767_)
  );
  al_aoi21 _07935_ (
    .a(_00461_),
    .b(_00455_),
    .c(\DFF_207.Q ),
    .y(_02768_)
  );
  al_ao21ftf _07936_ (
    .a(_02768_),
    .b(_01221_),
    .c(_01226_),
    .y(_02769_)
  );
  al_aoi21ftf _07937_ (
    .a(\DFF_647.Q ),
    .b(_02767_),
    .c(_02769_),
    .y(\DFF_207.D )
  );
  al_oai21ftf _07938_ (
    .a(\DFF_1316.Q ),
    .b(\DFF_377.Q ),
    .c(\DFF_838.Q ),
    .y(_02770_)
  );
  al_nand3ftt _07939_ (
    .a(\DFF_86.Q ),
    .b(g35),
    .c(_02770_),
    .y(_02771_)
  );
  al_ao21ftf _07940_ (
    .a(g35),
    .b(\DFF_377.Q ),
    .c(_02771_),
    .y(\DFF_838.D )
  );
  al_nand3 _07941_ (
    .a(_00499_),
    .b(_02682_),
    .c(_02754_),
    .y(_02772_)
  );
  al_ao21 _07942_ (
    .a(_02754_),
    .b(_02682_),
    .c(\DFF_670.Q ),
    .y(_02773_)
  );
  al_nand3 _07943_ (
    .a(g35),
    .b(_02773_),
    .c(_02772_),
    .y(_02774_)
  );
  al_ao21ftf _07944_ (
    .a(g35),
    .b(\DFF_370.Q ),
    .c(_02774_),
    .y(\DFF_670.D )
  );
  al_aoi21ftf _07945_ (
    .a(_00543_),
    .b(\DFF_319.Q ),
    .c(_00562_),
    .y(_02775_)
  );
  al_nand3 _07946_ (
    .a(\DFF_103.Q ),
    .b(\DFF_705.Q ),
    .c(_02775_),
    .y(_02776_)
  );
  al_nand2 _07947_ (
    .a(g35),
    .b(_02776_),
    .y(_02777_)
  );
  al_mux2l _07948_ (
    .a(\DFF_1184.Q ),
    .b(\DFF_1369.Q ),
    .s(_02777_),
    .y(\DFF_1369.D )
  );
  al_or2 _07949_ (
    .a(\DFF_468.Q ),
    .b(\DFF_942.Q ),
    .y(_02778_)
  );
  al_ao21ttf _07950_ (
    .a(\DFF_1420.Q ),
    .b(\DFF_468.Q ),
    .c(_02778_),
    .y(_02779_)
  );
  al_or3 _07951_ (
    .a(\DFF_220.Q ),
    .b(\DFF_81.Q ),
    .c(\DFF_34.Q ),
    .y(_02780_)
  );
  al_and3ftt _07952_ (
    .a(_02780_),
    .b(g35),
    .c(_02779_),
    .y(\DFF_1420.D )
  );
  al_or2 _07953_ (
    .a(_01614_),
    .b(_00641_),
    .y(_02781_)
  );
  al_and3ftt _07954_ (
    .a(_01844_),
    .b(_01615_),
    .c(_00641_),
    .y(_02782_)
  );
  al_nand2 _07955_ (
    .a(_02782_),
    .b(_02348_),
    .y(_02783_)
  );
  al_aoi21 _07956_ (
    .a(_02781_),
    .b(_02783_),
    .c(_00066_),
    .y(\DFF_713.D )
  );
  al_mux2h _07957_ (
    .a(\DFF_1423.Q ),
    .b(_01934_),
    .s(_00369_),
    .y(_02784_)
  );
  al_mux2h _07958_ (
    .a(\DFF_55.Q ),
    .b(_02784_),
    .s(g35),
    .y(\DFF_1423.D )
  );
  al_nand2ft _07959_ (
    .a(g35),
    .b(\DFF_154.Q ),
    .y(_02785_)
  );
  al_nand3 _07960_ (
    .a(\DFF_860.Q ),
    .b(\DFF_154.Q ),
    .c(_01761_),
    .y(_02786_)
  );
  al_aoi21ttf _07961_ (
    .a(_00355_),
    .b(_02786_),
    .c(_01760_),
    .y(_02787_)
  );
  al_ao21ftf _07962_ (
    .a(_01833_),
    .b(_02787_),
    .c(_02785_),
    .y(\DFF_411.D )
  );
  al_nand2 _07963_ (
    .a(\DFF_845.Q ),
    .b(_01964_),
    .y(_02788_)
  );
  al_or2 _07964_ (
    .a(\DFF_845.Q ),
    .b(_01964_),
    .y(_02789_)
  );
  al_ao21 _07965_ (
    .a(_02788_),
    .b(_02789_),
    .c(_01963_),
    .y(_02790_)
  );
  al_aoi21ftf _07966_ (
    .a(\DFF_746.Q ),
    .b(_00066_),
    .c(_02790_),
    .y(\DFF_845.D )
  );
  al_nand2ft _07967_ (
    .a(g35),
    .b(\DFF_599.Q ),
    .y(_02791_)
  );
  al_ao21ftf _07968_ (
    .a(\DFF_1404.Q ),
    .b(_00730_),
    .c(_02791_),
    .y(\DFF_1162.D )
  );
  al_oa21ftt _07969_ (
    .a(g35),
    .b(\DFF_57.Q ),
    .c(\DFF_1377.Q ),
    .y(\DFF_1249.D )
  );
  al_and2ft _07970_ (
    .a(\DFF_159.Q ),
    .b(\DFF_250.Q ),
    .y(_02792_)
  );
  al_ao21ftf _07971_ (
    .a(_02792_),
    .b(_00506_),
    .c(_00505_),
    .y(_02793_)
  );
  al_nand3 _07972_ (
    .a(g35),
    .b(_02793_),
    .c(_00981_),
    .y(_02794_)
  );
  al_aoi21ftf _07973_ (
    .a(\DFF_482.Q ),
    .b(_00066_),
    .c(_02794_),
    .y(\DFF_250.D )
  );
  al_inv _07974_ (
    .a(\DFF_403.Q ),
    .y(_02795_)
  );
  al_and3 _07975_ (
    .a(\DFF_1148.Q ),
    .b(\DFF_717.Q ),
    .c(\DFF_327.Q ),
    .y(_02796_)
  );
  al_nand3fft _07976_ (
    .a(\DFF_1092.Q ),
    .b(\DFF_595.Q ),
    .c(_00516_),
    .y(_02797_)
  );
  al_ao21ftf _07977_ (
    .a(\DFF_1092.Q ),
    .b(_00516_),
    .c(\DFF_595.Q ),
    .y(_02798_)
  );
  al_nand3 _07978_ (
    .a(_02796_),
    .b(_02797_),
    .c(_02798_),
    .y(_02799_)
  );
  al_nor2 _07979_ (
    .a(\DFF_182.Q ),
    .b(\DFF_822.Q ),
    .y(_02800_)
  );
  al_ao21 _07980_ (
    .a(_02800_),
    .b(_02796_),
    .c(\DFF_424.Q ),
    .y(_02801_)
  );
  al_nand3 _07981_ (
    .a(g35),
    .b(_02801_),
    .c(_02799_),
    .y(_02802_)
  );
  al_ao21ftf _07982_ (
    .a(_02795_),
    .b(_00066_),
    .c(_02802_),
    .y(\DFF_424.D )
  );
  al_inv _07983_ (
    .a(\DFF_104.Q ),
    .y(_02803_)
  );
  al_nand3 _07984_ (
    .a(\DFF_411.Q ),
    .b(_00556_),
    .c(_00357_),
    .y(_02804_)
  );
  al_nand3 _07985_ (
    .a(_02803_),
    .b(_02625_),
    .c(_02804_),
    .y(_02805_)
  );
  al_ao21ftf _07986_ (
    .a(g35),
    .b(\DFF_653.Q ),
    .c(_02805_),
    .y(\DFF_104.D )
  );
  al_nand2ft _07987_ (
    .a(\DFF_209.Q ),
    .b(\DFF_1010.Q ),
    .y(_02806_)
  );
  al_nand3ftt _07988_ (
    .a(_02806_),
    .b(_00526_),
    .c(_00530_),
    .y(_02807_)
  );
  al_ao21ftt _07989_ (
    .a(_02806_),
    .b(_00526_),
    .c(\DFF_625.Q ),
    .y(_02808_)
  );
  al_nand3 _07990_ (
    .a(g35),
    .b(_02808_),
    .c(_02807_),
    .y(_02809_)
  );
  al_ao21ftf _07991_ (
    .a(g35),
    .b(\DFF_469.Q ),
    .c(_02809_),
    .y(\DFF_625.D )
  );
  al_mux2l _07992_ (
    .a(\DFF_663.Q ),
    .b(\DFF_1221.Q ),
    .s(g35),
    .y(\DFF_159.D )
  );
  al_oa21ttf _07993_ (
    .a(\DFF_259.Q ),
    .b(\DFF_205.Q ),
    .c(\DFF_976.Q ),
    .y(_02810_)
  );
  al_nand3 _07994_ (
    .a(_02810_),
    .b(_01947_),
    .c(_01943_),
    .y(_02811_)
  );
  al_or3ftt _07995_ (
    .a(\DFF_976.Q ),
    .b(\DFF_259.Q ),
    .c(\DFF_205.Q ),
    .y(_02812_)
  );
  al_nand3 _07996_ (
    .a(g35),
    .b(_02812_),
    .c(_02811_),
    .y(_02813_)
  );
  al_aoi21ftf _07997_ (
    .a(\DFF_205.Q ),
    .b(_00066_),
    .c(_02813_),
    .y(\DFF_976.D )
  );
  al_mux2l _07998_ (
    .a(\DFF_994.Q ),
    .b(\DFF_1357.Q ),
    .s(g35),
    .y(\DFF_994.D )
  );
  al_mux2l _07999_ (
    .a(\DFF_445.Q ),
    .b(\DFF_941.Q ),
    .s(g35),
    .y(\DFF_445.D )
  );
  al_nand3ftt _08000_ (
    .a(_01311_),
    .b(_01408_),
    .c(_00499_),
    .y(_02814_)
  );
  al_ao21ftt _08001_ (
    .a(_01311_),
    .b(_01408_),
    .c(\DFF_602.Q ),
    .y(_02815_)
  );
  al_nand3 _08002_ (
    .a(g35),
    .b(_02814_),
    .c(_02815_),
    .y(_02816_)
  );
  al_ao21ftf _08003_ (
    .a(g35),
    .b(\DFF_750.Q ),
    .c(_02816_),
    .y(\DFF_602.D )
  );
  al_nand2 _08004_ (
    .a(\DFF_461.Q ),
    .b(_00459_),
    .y(_02817_)
  );
  al_or2 _08005_ (
    .a(\DFF_461.Q ),
    .b(_00459_),
    .y(_02818_)
  );
  al_and3 _08006_ (
    .a(_02817_),
    .b(_02818_),
    .c(_01731_),
    .y(_02819_)
  );
  al_mux2h _08007_ (
    .a(\DFF_1373.Q ),
    .b(_02819_),
    .s(g35),
    .y(\DFF_461.D )
  );
  al_and2 _08008_ (
    .a(\DFF_993.Q ),
    .b(\DFF_1091.Q ),
    .y(_02820_)
  );
  al_ao21 _08009_ (
    .a(_02820_),
    .b(_00576_),
    .c(_00066_),
    .y(_02821_)
  );
  al_mux2l _08010_ (
    .a(\DFF_835.Q ),
    .b(\DFF_558.Q ),
    .s(_02821_),
    .y(\DFF_558.D )
  );
  al_ao21 _08011_ (
    .a(\DFF_604.Q ),
    .b(_00459_),
    .c(\DFF_452.Q ),
    .y(_02822_)
  );
  al_nand3ftt _08012_ (
    .a(_01323_),
    .b(_02822_),
    .c(_01319_),
    .y(_02823_)
  );
  al_ao21ftf _08013_ (
    .a(g35),
    .b(\DFF_1191.Q ),
    .c(_02823_),
    .y(\DFF_452.D )
  );
  al_and2 _08014_ (
    .a(\DFF_278.Q ),
    .b(\DFF_870.Q ),
    .y(_02824_)
  );
  al_nand3 _08015_ (
    .a(\DFF_525.Q ),
    .b(_02824_),
    .c(_01050_),
    .y(_02825_)
  );
  al_aoi21ftf _08016_ (
    .a(\DFF_710.Q ),
    .b(_02825_),
    .c(_02027_),
    .y(_02826_)
  );
  al_ao21ftf _08017_ (
    .a(_02825_),
    .b(\DFF_710.Q ),
    .c(_02826_),
    .y(_02827_)
  );
  al_ao21ftf _08018_ (
    .a(g35),
    .b(\DFF_278.Q ),
    .c(_02827_),
    .y(\DFF_710.D )
  );
  al_nand3 _08019_ (
    .a(\DFF_913.Q ),
    .b(\DFF_454.Q ),
    .c(_01317_),
    .y(_02828_)
  );
  al_and2 _08020_ (
    .a(\DFF_1275.Q ),
    .b(\DFF_1109.Q ),
    .y(_02829_)
  );
  al_aoi21ftf _08021_ (
    .a(_02829_),
    .b(_02828_),
    .c(g35),
    .y(_02830_)
  );
  al_ao21ftf _08022_ (
    .a(_02828_),
    .b(\DFF_1109.Q ),
    .c(_02830_),
    .y(_02831_)
  );
  al_ao21ftf _08023_ (
    .a(g35),
    .b(\DFF_913.Q ),
    .c(_02831_),
    .y(\DFF_1109.D )
  );
  al_oa21 _08024_ (
    .a(_00705_),
    .b(_02114_),
    .c(_01359_),
    .y(_02832_)
  );
  al_mux2h _08025_ (
    .a(\DFF_35.Q ),
    .b(_02832_),
    .s(g35),
    .y(\DFF_803.D )
  );
  al_mux2l _08026_ (
    .a(\DFF_1275.Q ),
    .b(\DFF_171.Q ),
    .s(g35),
    .y(\DFF_67.D )
  );
  al_ao21 _08027_ (
    .a(\DFF_860.Q ),
    .b(_01761_),
    .c(\DFF_154.Q ),
    .y(_02833_)
  );
  al_ao21ttf _08028_ (
    .a(_02786_),
    .b(_02833_),
    .c(_01760_),
    .y(_02834_)
  );
  al_aoi21ftf _08029_ (
    .a(\DFF_860.Q ),
    .b(_00066_),
    .c(_02834_),
    .y(\DFF_154.D )
  );
  al_and2ft _08030_ (
    .a(g35),
    .b(\DFF_676.Q ),
    .y(_02835_)
  );
  al_mux2h _08031_ (
    .a(_01998_),
    .b(_01994_),
    .s(\DFF_676.Q ),
    .y(_02836_)
  );
  al_ao21ftf _08032_ (
    .a(_02836_),
    .b(_02164_),
    .c(\DFF_1246.Q ),
    .y(_02837_)
  );
  al_oa21ttf _08033_ (
    .a(\DFF_1246.Q ),
    .b(_02836_),
    .c(_00066_),
    .y(_02838_)
  );
  al_ao21 _08034_ (
    .a(_02838_),
    .b(_02837_),
    .c(_02835_),
    .y(\DFF_1246.D )
  );
  al_nor2 _08035_ (
    .a(g35),
    .b(\DFF_781.Q ),
    .y(_02839_)
  );
  al_and3fft _08036_ (
    .a(_00620_),
    .b(_00634_),
    .c(g35),
    .y(_02840_)
  );
  al_aoi21 _08037_ (
    .a(_00261_),
    .b(_02840_),
    .c(_02839_),
    .y(\DFF_223.D )
  );
  al_and2 _08038_ (
    .a(\DFF_88.Q ),
    .b(_01184_),
    .y(_02841_)
  );
  al_nand2ft _08039_ (
    .a(g35),
    .b(\DFF_7.Q ),
    .y(_02842_)
  );
  al_or2 _08040_ (
    .a(\DFF_88.Q ),
    .b(_01184_),
    .y(_02843_)
  );
  al_nand2 _08041_ (
    .a(\DFF_844.Q ),
    .b(\DFF_338.Q ),
    .y(_02844_)
  );
  al_and3 _08042_ (
    .a(_02276_),
    .b(_02844_),
    .c(_02843_),
    .y(_02845_)
  );
  al_ao21ftf _08043_ (
    .a(_02841_),
    .b(_02845_),
    .c(_02842_),
    .y(\DFF_88.D )
  );
  al_mux2l _08044_ (
    .a(\DFF_143.Q ),
    .b(\DFF_1194.Q ),
    .s(g35),
    .y(\DFF_1275.D )
  );
  al_nand3 _08045_ (
    .a(\DFF_286.Q ),
    .b(\DFF_517.Q ),
    .c(_00585_),
    .y(_02846_)
  );
  al_ao21 _08046_ (
    .a(\DFF_286.Q ),
    .b(_00585_),
    .c(\DFF_517.Q ),
    .y(_02847_)
  );
  al_and3 _08047_ (
    .a(_02846_),
    .b(_02847_),
    .c(_00588_),
    .y(_02848_)
  );
  al_mux2h _08048_ (
    .a(\DFF_286.Q ),
    .b(_02848_),
    .s(g35),
    .y(\DFF_517.D )
  );
  al_and2ft _08049_ (
    .a(g35),
    .b(\DFF_862.Q ),
    .y(_02849_)
  );
  al_ao21ftf _08050_ (
    .a(_01371_),
    .b(_01362_),
    .c(_02040_),
    .y(_02850_)
  );
  al_oa21ftf _08051_ (
    .a(_01361_),
    .b(_01363_),
    .c(_00066_),
    .y(_02851_)
  );
  al_ao21 _08052_ (
    .a(_02851_),
    .b(_02850_),
    .c(_02849_),
    .y(\DFF_1070.D )
  );
  al_and2ft _08053_ (
    .a(g35),
    .b(\DFF_713.Q ),
    .y(_02852_)
  );
  al_and3ftt _08054_ (
    .a(_00640_),
    .b(_00604_),
    .c(_02347_),
    .y(_02853_)
  );
  al_oai21ftt _08055_ (
    .a(\DFF_505.Q ),
    .b(\DFF_402.Q ),
    .c(\DFF_1181.Q ),
    .y(_02854_)
  );
  al_or3ftt _08056_ (
    .a(\DFF_505.Q ),
    .b(\DFF_402.Q ),
    .c(\DFF_1181.Q ),
    .y(_02855_)
  );
  al_nand3 _08057_ (
    .a(_02854_),
    .b(_02855_),
    .c(_02853_),
    .y(_02856_)
  );
  al_oa21ftf _08058_ (
    .a(_02345_),
    .b(_02853_),
    .c(_00066_),
    .y(_02857_)
  );
  al_ao21 _08059_ (
    .a(_02856_),
    .b(_02857_),
    .c(_02852_),
    .y(\DFF_594.D )
  );
  al_oa21ttf _08060_ (
    .a(\DFF_539.Q ),
    .b(\DFF_1392.Q ),
    .c(\DFF_191.Q ),
    .y(_02858_)
  );
  al_nand3 _08061_ (
    .a(_02858_),
    .b(_01335_),
    .c(_01337_),
    .y(_02859_)
  );
  al_and3fft _08062_ (
    .a(\DFF_539.Q ),
    .b(\DFF_1392.Q ),
    .c(\DFF_191.Q ),
    .y(_02860_)
  );
  al_nand3ftt _08063_ (
    .a(_02860_),
    .b(g35),
    .c(_02859_),
    .y(_02861_)
  );
  al_aoi21ftf _08064_ (
    .a(\DFF_1392.Q ),
    .b(_00066_),
    .c(_02861_),
    .y(\DFF_191.D )
  );
  al_nor2 _08065_ (
    .a(\DFF_519.Q ),
    .b(\DFF_385.Q ),
    .y(_02862_)
  );
  al_nand3 _08066_ (
    .a(_00499_),
    .b(_01467_),
    .c(_02862_),
    .y(_02863_)
  );
  al_ao21 _08067_ (
    .a(_02862_),
    .b(_01467_),
    .c(\DFF_877.Q ),
    .y(_02864_)
  );
  al_nand3 _08068_ (
    .a(g35),
    .b(_02864_),
    .c(_02863_),
    .y(_02865_)
  );
  al_ao21ftf _08069_ (
    .a(g35),
    .b(\DFF_192.Q ),
    .c(_02865_),
    .y(\DFF_877.D )
  );
  al_mux2l _08070_ (
    .a(\DFF_346.Q ),
    .b(\DFF_652.Q ),
    .s(_00478_),
    .y(_02866_)
  );
  al_mux2h _08071_ (
    .a(\DFF_533.Q ),
    .b(_02866_),
    .s(g35),
    .y(\DFF_652.D )
  );
  al_nor2 _08072_ (
    .a(\DFF_237.Q ),
    .b(g35),
    .y(_02867_)
  );
  al_oa21ftf _08073_ (
    .a(_01579_),
    .b(_00911_),
    .c(_02867_),
    .y(_02868_)
  );
  al_oa21 _08074_ (
    .a(\DFF_1315.Q ),
    .b(_01174_),
    .c(_02868_),
    .y(\DFF_1315.D )
  );
  al_aoi21 _08075_ (
    .a(\DFF_90.Q ),
    .b(g35),
    .c(\DFF_295.Q ),
    .y(_02869_)
  );
  al_and2 _08076_ (
    .a(\DFF_90.Q ),
    .b(\DFF_295.Q ),
    .y(_02870_)
  );
  al_aoi21 _08077_ (
    .a(g35),
    .b(_02870_),
    .c(_02869_),
    .y(\DFF_90.D )
  );
  al_and2ft _08078_ (
    .a(\DFF_723.Q ),
    .b(\DFF_734.Q ),
    .y(_02871_)
  );
  al_nand3 _08079_ (
    .a(_00499_),
    .b(_02665_),
    .c(_02871_),
    .y(_02872_)
  );
  al_ao21 _08080_ (
    .a(_02665_),
    .b(_02871_),
    .c(\DFF_1058.Q ),
    .y(_02873_)
  );
  al_nand3 _08081_ (
    .a(g35),
    .b(_02873_),
    .c(_02872_),
    .y(_02874_)
  );
  al_ao21ftf _08082_ (
    .a(g35),
    .b(\DFF_1291.Q ),
    .c(_02874_),
    .y(\DFF_1058.D )
  );
  al_nor2 _08083_ (
    .a(\DFF_174.Q ),
    .b(g35),
    .y(_02875_)
  );
  al_and3 _08084_ (
    .a(_00604_),
    .b(_02775_),
    .c(_00430_),
    .y(_02876_)
  );
  al_nand3ftt _08085_ (
    .a(\DFF_174.Q ),
    .b(\DFF_103.Q ),
    .c(\DFF_379.Q ),
    .y(_02877_)
  );
  al_oai21ftf _08086_ (
    .a(\DFF_103.Q ),
    .b(\DFF_174.Q ),
    .c(\DFF_379.Q ),
    .y(_02878_)
  );
  al_nand3 _08087_ (
    .a(_02877_),
    .b(_02878_),
    .c(_02876_),
    .y(_02879_)
  );
  al_oa21ftf _08088_ (
    .a(\DFF_1063.Q ),
    .b(_02876_),
    .c(_00066_),
    .y(_02880_)
  );
  al_aoi21 _08089_ (
    .a(_02879_),
    .b(_02880_),
    .c(_02875_),
    .y(\DFF_1063.D )
  );
  al_mux2h _08090_ (
    .a(\DFF_787.Q ),
    .b(_01335_),
    .s(g35),
    .y(\DFF_1367.D )
  );
  al_mux2h _08091_ (
    .a(\DFF_548.Q ),
    .b(_01637_),
    .s(g35),
    .y(\DFF_1385.D )
  );
  al_nor2 _08092_ (
    .a(g35),
    .b(\DFF_1254.Q ),
    .y(_02881_)
  );
  al_and2 _08093_ (
    .a(\DFF_622.Q ),
    .b(_00328_),
    .y(_02882_)
  );
  al_nand3 _08094_ (
    .a(\DFF_1181.Q ),
    .b(_00604_),
    .c(_02882_),
    .y(_02883_)
  );
  al_nand3 _08095_ (
    .a(\DFF_1143.Q ),
    .b(_00974_),
    .c(_02883_),
    .y(_02884_)
  );
  al_oa21ftf _08096_ (
    .a(\DFF_265.Q ),
    .b(_00974_),
    .c(_00066_),
    .y(_02885_)
  );
  al_aoi21 _08097_ (
    .a(_02885_),
    .b(_02884_),
    .c(_02881_),
    .y(\DFF_265.D )
  );
  al_nand3 _08098_ (
    .a(_00499_),
    .b(_01045_),
    .c(_02010_),
    .y(_02886_)
  );
  al_ao21 _08099_ (
    .a(_01045_),
    .b(_02010_),
    .c(\DFF_321.Q ),
    .y(_02887_)
  );
  al_nand3 _08100_ (
    .a(g35),
    .b(_02887_),
    .c(_02886_),
    .y(_02888_)
  );
  al_ao21ftf _08101_ (
    .a(g35),
    .b(\DFF_1259.Q ),
    .c(_02888_),
    .y(\DFF_321.D )
  );
  al_and3fft _08102_ (
    .a(\DFF_912.Q ),
    .b(\DFF_42.Q ),
    .c(g35),
    .y(_02889_)
  );
  al_oai21ftt _08103_ (
    .a(g35),
    .b(\DFF_42.Q ),
    .c(\DFF_912.Q ),
    .y(_02890_)
  );
  al_nand2ft _08104_ (
    .a(_02889_),
    .b(_02890_),
    .y(_02891_)
  );
  al_mux2l _08105_ (
    .a(_02891_),
    .b(\DFF_1179.Q ),
    .s(_01127_),
    .y(\DFF_1179.D )
  );
  al_and2ft _08106_ (
    .a(g35),
    .b(\DFF_467.Q ),
    .y(_02892_)
  );
  al_oa21ttf _08107_ (
    .a(\DFF_587.Q ),
    .b(_00733_),
    .c(_02694_),
    .y(_02893_)
  );
  al_ao21 _08108_ (
    .a(_02893_),
    .b(_00734_),
    .c(_02892_),
    .y(\DFF_587.D )
  );
  al_aoi21ftt _08109_ (
    .a(\DFF_66.Q ),
    .b(\DFF_1343.Q ),
    .c(_01696_),
    .y(_02894_)
  );
  al_and2ft _08110_ (
    .a(\DFF_211.Q ),
    .b(\DFF_1343.Q ),
    .y(_02895_)
  );
  al_mux2l _08111_ (
    .a(_02895_),
    .b(\DFF_211.Q ),
    .s(_02894_),
    .y(_02896_)
  );
  al_mux2h _08112_ (
    .a(\DFF_66.Q ),
    .b(_02896_),
    .s(g35),
    .y(\DFF_211.D )
  );
  al_or3fft _08113_ (
    .a(_00329_),
    .b(_00974_),
    .c(_00977_),
    .y(_02897_)
  );
  al_ao21 _08114_ (
    .a(_00329_),
    .b(_00974_),
    .c(\DFF_959.Q ),
    .y(_02898_)
  );
  al_nand3 _08115_ (
    .a(g35),
    .b(_02898_),
    .c(_02897_),
    .y(_02899_)
  );
  al_ao21ftf _08116_ (
    .a(g35),
    .b(\DFF_887.Q ),
    .c(_02899_),
    .y(\DFF_959.D )
  );
  al_oai21ftt _08117_ (
    .a(g35),
    .b(_00563_),
    .c(\DFF_989.Q ),
    .y(_02900_)
  );
  al_nand3 _08118_ (
    .a(\DFF_726.Q ),
    .b(g35),
    .c(_01009_),
    .y(_02901_)
  );
  al_and2ft _08119_ (
    .a(_02900_),
    .b(_02901_),
    .y(_02902_)
  );
  al_or2ft _08120_ (
    .a(_02900_),
    .b(_02901_),
    .y(_02903_)
  );
  al_nand2ft _08121_ (
    .a(_02902_),
    .b(_02903_),
    .y(\DFF_726.D )
  );
  al_oa21ftt _08122_ (
    .a(g35),
    .b(\DFF_250.Q ),
    .c(\DFF_159.Q ),
    .y(_02904_)
  );
  al_nor2 _08123_ (
    .a(_00503_),
    .b(_00505_),
    .y(_02905_)
  );
  al_ao21 _08124_ (
    .a(g35),
    .b(_02905_),
    .c(_02904_),
    .y(\DFF_234.D )
  );
  al_nand3ftt _08125_ (
    .a(\DFF_20.Q ),
    .b(\DFF_916.Q ),
    .c(\DFF_104.Q ),
    .y(_02906_)
  );
  al_aoi21ftf _08126_ (
    .a(\DFF_92.Q ),
    .b(_02906_),
    .c(g35),
    .y(_02907_)
  );
  al_ao21ftf _08127_ (
    .a(_02906_),
    .b(_00499_),
    .c(_02907_),
    .y(_02908_)
  );
  al_ao21ftf _08128_ (
    .a(g35),
    .b(\DFF_1123.Q ),
    .c(_02908_),
    .y(\DFF_92.D )
  );
  al_nand3 _08129_ (
    .a(_00499_),
    .b(_00567_),
    .c(_01312_),
    .y(_02909_)
  );
  al_ao21 _08130_ (
    .a(_01312_),
    .b(_00567_),
    .c(\DFF_1406.Q ),
    .y(_02910_)
  );
  al_nand3 _08131_ (
    .a(g35),
    .b(_02910_),
    .c(_02909_),
    .y(_02911_)
  );
  al_ao21ftf _08132_ (
    .a(g35),
    .b(\DFF_950.Q ),
    .c(_02911_),
    .y(\DFF_1406.D )
  );
  al_and2 _08133_ (
    .a(\DFF_655.Q ),
    .b(\DFF_165.Q ),
    .y(_02912_)
  );
  al_and3 _08134_ (
    .a(\DFF_927.Q ),
    .b(\DFF_906.Q ),
    .c(_02912_),
    .y(_02913_)
  );
  al_aoi21 _08135_ (
    .a(\DFF_141.Q ),
    .b(_02913_),
    .c(_00066_),
    .y(_02914_)
  );
  al_oai21 _08136_ (
    .a(\DFF_141.Q ),
    .b(_02913_),
    .c(_02914_),
    .y(_02915_)
  );
  al_ao21ftf _08137_ (
    .a(g35),
    .b(\DFF_281.Q ),
    .c(_02915_),
    .y(\DFF_141.D )
  );
  al_nand3fft _08138_ (
    .a(\DFF_1092.Q ),
    .b(\DFF_774.Q ),
    .c(_00516_),
    .y(_02916_)
  );
  al_ao21ftf _08139_ (
    .a(\DFF_1092.Q ),
    .b(_00516_),
    .c(\DFF_774.Q ),
    .y(_02917_)
  );
  al_nand3 _08140_ (
    .a(_01260_),
    .b(_02916_),
    .c(_02917_),
    .y(_02918_)
  );
  al_ao21 _08141_ (
    .a(_01260_),
    .b(_02800_),
    .c(\DFF_169.Q ),
    .y(_02919_)
  );
  al_nand3 _08142_ (
    .a(g35),
    .b(_02919_),
    .c(_02918_),
    .y(_02920_)
  );
  al_ao21ftf _08143_ (
    .a(g35),
    .b(\DFF_182.Q ),
    .c(_02920_),
    .y(\DFF_169.D )
  );
  al_and2ft _08144_ (
    .a(g35),
    .b(\DFF_777.Q ),
    .y(_02921_)
  );
  al_and2ft _08145_ (
    .a(\DFF_705.Q ),
    .b(\DFF_174.Q ),
    .y(_02922_)
  );
  al_nand2 _08146_ (
    .a(_02922_),
    .b(_02775_),
    .y(_02923_)
  );
  al_nand2ft _08147_ (
    .a(\DFF_832.Q ),
    .b(\DFF_777.Q ),
    .y(_02924_)
  );
  al_nand2ft _08148_ (
    .a(\DFF_777.Q ),
    .b(\DFF_832.Q ),
    .y(_02925_)
  );
  al_or3fft _08149_ (
    .a(_02924_),
    .b(_02925_),
    .c(_02923_),
    .y(_02926_)
  );
  al_aoi21ftf _08150_ (
    .a(\DFF_1216.Q ),
    .b(_02923_),
    .c(g35),
    .y(_02927_)
  );
  al_ao21 _08151_ (
    .a(_02926_),
    .b(_02927_),
    .c(_02921_),
    .y(\DFF_1216.D )
  );
  al_ao21 _08152_ (
    .a(\DFF_812.Q ),
    .b(_01236_),
    .c(\DFF_751.Q ),
    .y(_02928_)
  );
  al_nand3 _08153_ (
    .a(_02276_),
    .b(_01237_),
    .c(_02928_),
    .y(_02929_)
  );
  al_ao21ftf _08154_ (
    .a(g35),
    .b(\DFF_812.Q ),
    .c(_02929_),
    .y(\DFF_751.D )
  );
  al_nor2 _08155_ (
    .a(\DFF_20.Q ),
    .b(\DFF_916.Q ),
    .y(_02930_)
  );
  al_nand3 _08156_ (
    .a(_00499_),
    .b(_02930_),
    .c(_02625_),
    .y(_02931_)
  );
  al_ao21 _08157_ (
    .a(_02930_),
    .b(_02625_),
    .c(\DFF_1366.Q ),
    .y(_02932_)
  );
  al_nand3 _08158_ (
    .a(g35),
    .b(_02932_),
    .c(_02931_),
    .y(_02933_)
  );
  al_ao21ftf _08159_ (
    .a(g35),
    .b(\DFF_397.Q ),
    .c(_02933_),
    .y(\DFF_1366.D )
  );
  al_mux2h _08160_ (
    .a(\DFF_1356.Q ),
    .b(_01934_),
    .s(_00378_),
    .y(_02934_)
  );
  al_mux2h _08161_ (
    .a(\DFF_1177.Q ),
    .b(_02934_),
    .s(g35),
    .y(\DFF_1356.D )
  );
  al_nand3ftt _08162_ (
    .a(_02686_),
    .b(_00431_),
    .c(_02775_),
    .y(_02935_)
  );
  al_ao21 _08163_ (
    .a(_00431_),
    .b(_02775_),
    .c(\DFF_1202.Q ),
    .y(_02936_)
  );
  al_nand3 _08164_ (
    .a(g35),
    .b(_02935_),
    .c(_02936_),
    .y(_02937_)
  );
  al_ao21ftf _08165_ (
    .a(g35),
    .b(\DFF_2.Q ),
    .c(_02937_),
    .y(\DFF_1202.D )
  );
  al_ao21 _08166_ (
    .a(g35),
    .b(\DFF_1134.Q ),
    .c(\DFF_58.Q ),
    .y(_02938_)
  );
  al_aoi21 _08167_ (
    .a(g35),
    .b(_00809_),
    .c(_02938_),
    .y(_02939_)
  );
  al_ao21ttf _08168_ (
    .a(_00793_),
    .b(_00766_),
    .c(\DFF_688.Q ),
    .y(_02940_)
  );
  al_nand2 _08169_ (
    .a(\DFF_58.Q ),
    .b(\DFF_1134.Q ),
    .y(_02941_)
  );
  al_oa21ftf _08170_ (
    .a(_02941_),
    .b(_00809_),
    .c(_00066_),
    .y(_02942_)
  );
  al_aoi21 _08171_ (
    .a(_02940_),
    .b(_02942_),
    .c(_02939_),
    .y(\DFF_688.D )
  );
  al_nand2 _08172_ (
    .a(\DFF_1148.Q ),
    .b(\DFF_60.Q ),
    .y(_02943_)
  );
  al_nor2 _08173_ (
    .a(\DFF_1148.Q ),
    .b(\DFF_60.Q ),
    .y(_02944_)
  );
  al_nand2ft _08174_ (
    .a(_02944_),
    .b(_02943_),
    .y(_02945_)
  );
  al_aoi21 _08175_ (
    .a(_02945_),
    .b(_02740_),
    .c(_00066_),
    .y(\DFF_1148.D )
  );
  al_nor2 _08176_ (
    .a(\DFF_516.Q ),
    .b(g35),
    .y(_02946_)
  );
  al_mux2l _08177_ (
    .a(\DFF_478.Q ),
    .b(\DFF_405.Q ),
    .s(\DFF_516.Q ),
    .y(_02947_)
  );
  al_nand3ftt _08178_ (
    .a(_02947_),
    .b(\DFF_475.Q ),
    .c(_01642_),
    .y(_02948_)
  );
  al_aoi21ftf _08179_ (
    .a(\DFF_475.Q ),
    .b(_02947_),
    .c(g35),
    .y(_02949_)
  );
  al_aoi21 _08180_ (
    .a(_02949_),
    .b(_02948_),
    .c(_02946_),
    .y(\DFF_475.D )
  );
  al_nand3ftt _08181_ (
    .a(_01920_),
    .b(_00305_),
    .c(_00852_),
    .y(_02950_)
  );
  al_mux2l _08182_ (
    .a(\DFF_247.Q ),
    .b(\DFF_282.Q ),
    .s(_02950_),
    .y(_02951_)
  );
  al_mux2h _08183_ (
    .a(\DFF_114.Q ),
    .b(_02951_),
    .s(g35),
    .y(\DFF_247.D )
  );
  al_and2ft _08184_ (
    .a(g35),
    .b(\DFF_1413.Q ),
    .y(_02952_)
  );
  al_and3ftt _08185_ (
    .a(_01149_),
    .b(_00604_),
    .c(_00323_),
    .y(_02953_)
  );
  al_oai21ftt _08186_ (
    .a(\DFF_996.Q ),
    .b(\DFF_671.Q ),
    .c(\DFF_1181.Q ),
    .y(_02954_)
  );
  al_or3ftt _08187_ (
    .a(\DFF_996.Q ),
    .b(\DFF_671.Q ),
    .c(\DFF_1181.Q ),
    .y(_02955_)
  );
  al_nand3 _08188_ (
    .a(_02954_),
    .b(_02955_),
    .c(_02953_),
    .y(_02956_)
  );
  al_oa21ftf _08189_ (
    .a(_02591_),
    .b(_02953_),
    .c(_00066_),
    .y(_02957_)
  );
  al_ao21 _08190_ (
    .a(_02956_),
    .b(_02957_),
    .c(_02952_),
    .y(\DFF_472.D )
  );
  al_oa21ftt _08191_ (
    .a(g35),
    .b(\DFF_636.Q ),
    .c(\DFF_415.Q ),
    .y(_02958_)
  );
  al_oa21ftf _08192_ (
    .a(\DFF_572.Q ),
    .b(\DFF_466.Q ),
    .c(\DFF_636.Q ),
    .y(_02959_)
  );
  al_ao21ftf _08193_ (
    .a(\DFF_415.Q ),
    .b(_02959_),
    .c(_00886_),
    .y(_02960_)
  );
  al_ao21 _08194_ (
    .a(g35),
    .b(_02960_),
    .c(_02958_),
    .y(\DFF_636.D )
  );
  al_and2 _08195_ (
    .a(\DFF_700.Q ),
    .b(_00937_),
    .y(_02961_)
  );
  al_aoi21 _08196_ (
    .a(\DFF_359.Q ),
    .b(_02961_),
    .c(_00066_),
    .y(_02962_)
  );
  al_aoi21ftt _08197_ (
    .a(\DFF_708.Q ),
    .b(_00066_),
    .c(_02962_),
    .y(\DFF_258.D )
  );
  al_nor2 _08198_ (
    .a(g35),
    .b(\DFF_484.Q ),
    .y(_02963_)
  );
  al_nand2ft _08199_ (
    .a(\DFF_118.Q ),
    .b(\DFF_139.Q ),
    .y(_02964_)
  );
  al_nand2 _08200_ (
    .a(\DFF_123.Q ),
    .b(\DFF_314.Q ),
    .y(_02965_)
  );
  al_nand2 _08201_ (
    .a(\DFF_1123.Q ),
    .b(\DFF_898.Q ),
    .y(_02966_)
  );
  al_aoi21 _08202_ (
    .a(_02965_),
    .b(_02966_),
    .c(_02964_),
    .y(_02967_)
  );
  al_and2ft _08203_ (
    .a(\DFF_139.Q ),
    .b(\DFF_118.Q ),
    .y(_02968_)
  );
  al_nand2 _08204_ (
    .a(\DFF_92.Q ),
    .b(\DFF_53.Q ),
    .y(_02969_)
  );
  al_nand2 _08205_ (
    .a(\DFF_945.Q ),
    .b(\DFF_1119.Q ),
    .y(_02970_)
  );
  al_ao21ttf _08206_ (
    .a(_02969_),
    .b(_02970_),
    .c(_02968_),
    .y(_02971_)
  );
  al_and3fft _08207_ (
    .a(\DFF_118.Q ),
    .b(\DFF_139.Q ),
    .c(\DFF_905.Q ),
    .y(_02972_)
  );
  al_ao21 _08208_ (
    .a(\DFF_59.Q ),
    .b(_02972_),
    .c(\DFF_1005.Q ),
    .y(_02973_)
  );
  al_nand2 _08209_ (
    .a(\DFF_634.Q ),
    .b(\DFF_970.Q ),
    .y(_02974_)
  );
  al_nand2 _08210_ (
    .a(\DFF_554.Q ),
    .b(\DFF_158.Q ),
    .y(_02975_)
  );
  al_ao21ttf _08211_ (
    .a(_02974_),
    .b(_02975_),
    .c(_00394_),
    .y(_02976_)
  );
  al_and3ftt _08212_ (
    .a(_02973_),
    .b(_02971_),
    .c(_02976_),
    .y(_02977_)
  );
  al_nand3 _08213_ (
    .a(\DFF_1366.Q ),
    .b(\DFF_898.Q ),
    .c(_00394_),
    .y(_02978_)
  );
  al_nand3 _08214_ (
    .a(\DFF_397.Q ),
    .b(\DFF_905.Q ),
    .c(_02968_),
    .y(_02979_)
  );
  al_and3 _08215_ (
    .a(\DFF_1005.Q ),
    .b(_02979_),
    .c(_02978_),
    .y(_02980_)
  );
  al_or2 _08216_ (
    .a(\DFF_118.Q ),
    .b(\DFF_139.Q ),
    .y(_02981_)
  );
  al_nand2 _08217_ (
    .a(\DFF_579.Q ),
    .b(\DFF_1119.Q ),
    .y(_02982_)
  );
  al_nand2 _08218_ (
    .a(\DFF_337.Q ),
    .b(\DFF_53.Q ),
    .y(_02983_)
  );
  al_ao21 _08219_ (
    .a(_02982_),
    .b(_02983_),
    .c(_02981_),
    .y(_02984_)
  );
  al_nand2 _08220_ (
    .a(\DFF_1011.Q ),
    .b(\DFF_970.Q ),
    .y(_02985_)
  );
  al_nand2 _08221_ (
    .a(\DFF_554.Q ),
    .b(\DFF_494.Q ),
    .y(_02986_)
  );
  al_ao21 _08222_ (
    .a(_02985_),
    .b(_02986_),
    .c(_02964_),
    .y(_02987_)
  );
  al_nand3 _08223_ (
    .a(_02984_),
    .b(_02987_),
    .c(_02980_),
    .y(_02988_)
  );
  al_ao21ftf _08224_ (
    .a(_02967_),
    .b(_02977_),
    .c(_02988_),
    .y(_02989_)
  );
  al_nand2 _08225_ (
    .a(\DFF_484.Q ),
    .b(_01664_),
    .y(_02990_)
  );
  al_nor3fft _08226_ (
    .a(\DFF_188.Q ),
    .b(\DFF_483.Q ),
    .c(_02981_),
    .y(_02991_)
  );
  al_and3 _08227_ (
    .a(\DFF_315.Q ),
    .b(\DFF_298.Q ),
    .c(_02968_),
    .y(_02992_)
  );
  al_nor2 _08228_ (
    .a(\DFF_1005.Q ),
    .b(\DFF_554.Q ),
    .y(_02993_)
  );
  al_nand2 _08229_ (
    .a(\DFF_1005.Q ),
    .b(\DFF_554.Q ),
    .y(_02994_)
  );
  al_or3fft _08230_ (
    .a(\DFF_474.Q ),
    .b(\DFF_82.Q ),
    .c(_02964_),
    .y(_02995_)
  );
  al_and3ftt _08231_ (
    .a(_02993_),
    .b(_02994_),
    .c(_02995_),
    .y(_02996_)
  );
  al_nand3fft _08232_ (
    .a(_02991_),
    .b(_02992_),
    .c(_02996_),
    .y(_02997_)
  );
  al_nor3fft _08233_ (
    .a(\DFF_315.Q ),
    .b(\DFF_1307.Q ),
    .c(_02981_),
    .y(_02998_)
  );
  al_nand2ft _08234_ (
    .a(_02993_),
    .b(_02994_),
    .y(_02999_)
  );
  al_and3 _08235_ (
    .a(\DFF_188.Q ),
    .b(\DFF_179.Q ),
    .c(_02968_),
    .y(_03000_)
  );
  al_nand3 _08236_ (
    .a(\DFF_474.Q ),
    .b(\DFF_904.Q ),
    .c(_00394_),
    .y(_03001_)
  );
  al_and3ftt _08237_ (
    .a(_03000_),
    .b(_03001_),
    .c(_02999_),
    .y(_03002_)
  );
  al_ao21ftf _08238_ (
    .a(_02998_),
    .b(_03002_),
    .c(_02997_),
    .y(_03003_)
  );
  al_nand3 _08239_ (
    .a(_02990_),
    .b(_03003_),
    .c(_02989_),
    .y(_03004_)
  );
  al_nand2 _08240_ (
    .a(_01663_),
    .b(_03004_),
    .y(_03005_)
  );
  al_oa21ftf _08241_ (
    .a(\DFF_493.Q ),
    .b(_01663_),
    .c(_00066_),
    .y(_03006_)
  );
  al_aoi21 _08242_ (
    .a(_03006_),
    .b(_03005_),
    .c(_02963_),
    .y(\DFF_493.D )
  );
  al_aoi21 _08243_ (
    .a(\DFF_933.Q ),
    .b(_00642_),
    .c(_00066_),
    .y(_03007_)
  );
  al_oai21 _08244_ (
    .a(\DFF_933.Q ),
    .b(_00642_),
    .c(_03007_),
    .y(_03008_)
  );
  al_aoi21ftf _08245_ (
    .a(\DFF_1071.Q ),
    .b(_00066_),
    .c(_03008_),
    .y(\DFF_933.D )
  );
  al_ao21 _08246_ (
    .a(\DFF_62.Q ),
    .b(_01323_),
    .c(\DFF_894.Q ),
    .y(_03009_)
  );
  al_and3 _08247_ (
    .a(\DFF_894.Q ),
    .b(\DFF_62.Q ),
    .c(_01323_),
    .y(_03010_)
  );
  al_nand3ftt _08248_ (
    .a(_03010_),
    .b(_03009_),
    .c(_01319_),
    .y(_03011_)
  );
  al_ao21ftf _08249_ (
    .a(g35),
    .b(\DFF_62.Q ),
    .c(_03011_),
    .y(\DFF_894.D )
  );
  al_ao21ftt _08250_ (
    .a(\DFF_164.Q ),
    .b(_00550_),
    .c(\DFF_1036.Q ),
    .y(_03012_)
  );
  al_and2ft _08251_ (
    .a(g35),
    .b(\DFF_451.Q ),
    .y(_03013_)
  );
  al_ao21 _08252_ (
    .a(_00552_),
    .b(_03012_),
    .c(_03013_),
    .y(\DFF_1036.D )
  );
  al_nand3 _08253_ (
    .a(_00499_),
    .b(_02862_),
    .c(_02871_),
    .y(_03014_)
  );
  al_ao21 _08254_ (
    .a(_02871_),
    .b(_02862_),
    .c(\DFF_398.Q ),
    .y(_03015_)
  );
  al_nand3 _08255_ (
    .a(g35),
    .b(_03015_),
    .c(_03014_),
    .y(_03016_)
  );
  al_ao21ftf _08256_ (
    .a(g35),
    .b(\DFF_267.Q ),
    .c(_03016_),
    .y(\DFF_398.D )
  );
  al_nor2 _08257_ (
    .a(g35),
    .b(\DFF_1356.Q ),
    .y(_03017_)
  );
  al_oa21ftf _08258_ (
    .a(\DFF_535.Q ),
    .b(_00766_),
    .c(_00066_),
    .y(_03018_)
  );
  al_aoi21 _08259_ (
    .a(_03018_),
    .b(_00808_),
    .c(_03017_),
    .y(\DFF_535.D )
  );
  al_oa21ftt _08260_ (
    .a(g35),
    .b(\DFF_1190.Q ),
    .c(\DFF_73.Q ),
    .y(_03019_)
  );
  al_or3fft _08261_ (
    .a(\DFF_215.Q ),
    .b(g35),
    .c(_03019_),
    .y(_03020_)
  );
  al_aoi21ttf _08262_ (
    .a(\DFF_215.Q ),
    .b(g35),
    .c(_03019_),
    .y(_03021_)
  );
  al_nand2ft _08263_ (
    .a(_03021_),
    .b(_03020_),
    .y(\DFF_215.D )
  );
  al_oa21ftt _08264_ (
    .a(g35),
    .b(_00745_),
    .c(\DFF_699.Q ),
    .y(\DFF_635.D )
  );
  al_nand3fft _08265_ (
    .a(_01128_),
    .b(_01646_),
    .c(_01125_),
    .y(_03022_)
  );
  al_aoi21ftf _08266_ (
    .a(\DFF_2.Q ),
    .b(_03022_),
    .c(g35),
    .y(_03023_)
  );
  al_oai21 _08267_ (
    .a(_01131_),
    .b(_03022_),
    .c(_03023_),
    .y(_03024_)
  );
  al_ao21ftf _08268_ (
    .a(g35),
    .b(\DFF_968.Q ),
    .c(_03024_),
    .y(\DFF_2.D )
  );
  al_mux2l _08269_ (
    .a(\DFF_274.Q ),
    .b(\DFF_1383.Q ),
    .s(_02694_),
    .y(\DFF_1383.D )
  );
  al_nor3ftt _08270_ (
    .a(\DFF_1195.Q ),
    .b(_00499_),
    .c(_00361_),
    .y(_03025_)
  );
  al_oa21ftt _08271_ (
    .a(\DFF_1195.Q ),
    .b(_00361_),
    .c(_00499_),
    .y(_03026_)
  );
  al_nor3ftt _08272_ (
    .a(g35),
    .b(_03025_),
    .c(_03026_),
    .y(\DFF_1195.D )
  );
  al_and2 _08273_ (
    .a(\DFF_806.Q ),
    .b(\DFF_1158.Q ),
    .y(_03027_)
  );
  al_and3 _08274_ (
    .a(\DFF_1196.Q ),
    .b(\DFF_1248.Q ),
    .c(_03027_),
    .y(_03028_)
  );
  al_aoi21 _08275_ (
    .a(\DFF_198.Q ),
    .b(_03028_),
    .c(_00066_),
    .y(_03029_)
  );
  al_oai21 _08276_ (
    .a(\DFF_198.Q ),
    .b(_03028_),
    .c(_03029_),
    .y(_03030_)
  );
  al_ao21ftf _08277_ (
    .a(g35),
    .b(\DFF_1023.Q ),
    .c(_03030_),
    .y(\DFF_198.D )
  );
  al_mux2l _08278_ (
    .a(\DFF_496.Q ),
    .b(\DFF_1106.Q ),
    .s(_01557_),
    .y(_03031_)
  );
  al_mux2h _08279_ (
    .a(\DFF_771.Q ),
    .b(_03031_),
    .s(g35),
    .y(\DFF_496.D )
  );
  al_oai21ttf _08280_ (
    .a(\DFF_927.Q ),
    .b(\DFF_655.Q ),
    .c(_02912_),
    .y(_03032_)
  );
  al_nand2ft _08281_ (
    .a(\DFF_566.Q ),
    .b(\DFF_616.Q ),
    .y(_03033_)
  );
  al_nand2ft _08282_ (
    .a(\DFF_906.Q ),
    .b(\DFF_566.Q ),
    .y(_03034_)
  );
  al_aoi21ftf _08283_ (
    .a(\DFF_927.Q ),
    .b(\DFF_906.Q ),
    .c(_03034_),
    .y(_03035_)
  );
  al_and3 _08284_ (
    .a(g35),
    .b(_03033_),
    .c(_03035_),
    .y(_03036_)
  );
  al_and3ftt _08285_ (
    .a(_02913_),
    .b(_03032_),
    .c(_03036_),
    .y(\DFF_165.D )
  );
  al_oa21ftt _08286_ (
    .a(g35),
    .b(\DFF_1113.Q ),
    .c(\DFF_975.Q ),
    .y(\DFF_907.D )
  );
  al_nand3 _08287_ (
    .a(\DFF_463.Q ),
    .b(_01958_),
    .c(_02325_),
    .y(_03037_)
  );
  al_ao21 _08288_ (
    .a(\DFF_463.Q ),
    .b(_01958_),
    .c(_02325_),
    .y(_03038_)
  );
  al_nand3 _08289_ (
    .a(g35),
    .b(_03037_),
    .c(_03038_),
    .y(_03039_)
  );
  al_aoi21ftf _08290_ (
    .a(\DFF_14.Q ),
    .b(_00066_),
    .c(_03039_),
    .y(\DFF_463.D )
  );
  al_nand3 _08291_ (
    .a(_00499_),
    .b(_01701_),
    .c(_01744_),
    .y(_03040_)
  );
  al_ao21 _08292_ (
    .a(_01701_),
    .b(_01744_),
    .c(\DFF_1355.Q ),
    .y(_03041_)
  );
  al_nand3 _08293_ (
    .a(g35),
    .b(_03041_),
    .c(_03040_),
    .y(_03042_)
  );
  al_ao21ftf _08294_ (
    .a(g35),
    .b(\DFF_392.Q ),
    .c(_03042_),
    .y(\DFF_1355.D )
  );
  al_mux2l _08295_ (
    .a(\DFF_941.Q ),
    .b(\DFF_507.Q ),
    .s(g35),
    .y(\DFF_941.D )
  );
  al_oai21ftf _08296_ (
    .a(\DFF_525.Q ),
    .b(_02024_),
    .c(\DFF_278.Q ),
    .y(_03043_)
  );
  al_nand3 _08297_ (
    .a(_02027_),
    .b(_02825_),
    .c(_03043_),
    .y(_03044_)
  );
  al_ao21ftf _08298_ (
    .a(g35),
    .b(\DFF_525.Q ),
    .c(_03044_),
    .y(\DFF_278.D )
  );
  al_oa21ftf _08299_ (
    .a(\DFF_1348.Q ),
    .b(_00373_),
    .c(_00066_),
    .y(_03045_)
  );
  al_ao21ftf _08300_ (
    .a(_00499_),
    .b(_00373_),
    .c(_03045_),
    .y(_03046_)
  );
  al_aoi21ftf _08301_ (
    .a(\DFF_779.Q ),
    .b(_00066_),
    .c(_03046_),
    .y(\DFF_1348.D )
  );
  al_nand3 _08302_ (
    .a(\DFF_23.Q ),
    .b(\DFF_113.Q ),
    .c(_01050_),
    .y(_03047_)
  );
  al_nand3 _08303_ (
    .a(\DFF_524.Q ),
    .b(\DFF_872.Q ),
    .c(_03047_),
    .y(_03048_)
  );
  al_and3 _08304_ (
    .a(\DFF_23.Q ),
    .b(\DFF_1161.Q ),
    .c(_00477_),
    .y(_03049_)
  );
  al_nand3ftt _08305_ (
    .a(_02026_),
    .b(\DFF_113.Q ),
    .c(_03049_),
    .y(_03050_)
  );
  al_nand3 _08306_ (
    .a(g35),
    .b(_03050_),
    .c(_03048_),
    .y(_03051_)
  );
  al_aoi21ftf _08307_ (
    .a(\DFF_113.Q ),
    .b(_00066_),
    .c(_03051_),
    .y(\DFF_524.D )
  );
  al_mux2l _08308_ (
    .a(\DFF_731.Q ),
    .b(\DFF_543.Q ),
    .s(\DFF_833.Q ),
    .y(_03052_)
  );
  al_aoi21 _08309_ (
    .a(\DFF_429.Q ),
    .b(_03052_),
    .c(\DFF_647.Q ),
    .y(_03053_)
  );
  al_oai21 _08310_ (
    .a(\DFF_429.Q ),
    .b(_03052_),
    .c(_03053_),
    .y(_03054_)
  );
  al_ao21ttf _08311_ (
    .a(_02766_),
    .b(_03054_),
    .c(_01956_),
    .y(_03055_)
  );
  al_or2 _08312_ (
    .a(\DFF_647.Q ),
    .b(_01956_),
    .y(_03056_)
  );
  al_and3 _08313_ (
    .a(g35),
    .b(_03055_),
    .c(_03056_),
    .y(\DFF_647.D )
  );
  al_nand3ftt _08314_ (
    .a(_01921_),
    .b(_00305_),
    .c(_00852_),
    .y(_03057_)
  );
  al_mux2l _08315_ (
    .a(\DFF_114.Q ),
    .b(\DFF_282.Q ),
    .s(_03057_),
    .y(_03058_)
  );
  al_mux2h _08316_ (
    .a(\DFF_1152.Q ),
    .b(_03058_),
    .s(g35),
    .y(\DFF_114.D )
  );
  al_mux2l _08317_ (
    .a(\DFF_573.Q ),
    .b(\DFF_1365.Q ),
    .s(_01054_),
    .y(\DFF_1365.D )
  );
  al_inv _08318_ (
    .a(\DFF_567.Q ),
    .y(_03059_)
  );
  al_and2 _08319_ (
    .a(\DFF_272.Q ),
    .b(_01889_),
    .y(_03060_)
  );
  al_nand3 _08320_ (
    .a(\DFF_1181.Q ),
    .b(_00604_),
    .c(_00334_),
    .y(_03061_)
  );
  al_oa21ftf _08321_ (
    .a(\DFF_500.Q ),
    .b(_01889_),
    .c(_00066_),
    .y(_03062_)
  );
  al_ao21ttf _08322_ (
    .a(_03060_),
    .b(_03061_),
    .c(_03062_),
    .y(_03063_)
  );
  al_aoi21ftf _08323_ (
    .a(g35),
    .b(_03059_),
    .c(_03063_),
    .y(\DFF_500.D )
  );
  al_or3 _08324_ (
    .a(\DFF_803.Q ),
    .b(\DFF_35.Q ),
    .c(\DFF_54.Q ),
    .y(_03064_)
  );
  al_nand3ftt _08325_ (
    .a(_03064_),
    .b(_00499_),
    .c(_02681_),
    .y(_03065_)
  );
  al_ao21ftt _08326_ (
    .a(_03064_),
    .b(_02681_),
    .c(\DFF_1386.Q ),
    .y(_03066_)
  );
  al_nand3 _08327_ (
    .a(g35),
    .b(_03065_),
    .c(_03066_),
    .y(_03067_)
  );
  al_ao21ftf _08328_ (
    .a(g35),
    .b(\DFF_1263.Q ),
    .c(_03067_),
    .y(\DFF_1386.D )
  );
  al_oa21 _08329_ (
    .a(\DFF_1221.Q ),
    .b(\DFF_1397.Q ),
    .c(g35),
    .y(_03068_)
  );
  al_or3 _08330_ (
    .a(\DFF_688.Q ),
    .b(\DFF_742.Q ),
    .c(\DFF_1409.Q ),
    .y(_03069_)
  );
  al_ao21 _08331_ (
    .a(g35),
    .b(_03069_),
    .c(_03068_),
    .y(_03070_)
  );
  al_or2 _08332_ (
    .a(\DFF_1021.Q ),
    .b(\DFF_1121.Q ),
    .y(_03071_)
  );
  al_oai21ttf _08333_ (
    .a(\DFF_679.Q ),
    .b(_03071_),
    .c(_00066_),
    .y(_03072_)
  );
  al_oai21 _08334_ (
    .a(\DFF_987.Q ),
    .b(\DFF_1203.Q ),
    .c(g35),
    .y(_03073_)
  );
  al_and2 _08335_ (
    .a(_03073_),
    .b(_03072_),
    .y(_03074_)
  );
  al_nand3fft _08336_ (
    .a(\DFF_781.Q ),
    .b(_03070_),
    .c(_03074_),
    .y(_03075_)
  );
  al_mux2h _08337_ (
    .a(\DFF_1182.Q ),
    .b(_03075_),
    .s(g35),
    .y(\DFF_781.D )
  );
  al_mux2l _08338_ (
    .a(\DFF_538.Q ),
    .b(\DFF_259.Q ),
    .s(g35),
    .y(\DFF_1256.D )
  );
  al_nand3fft _08339_ (
    .a(\DFF_894.Q ),
    .b(\DFF_849.Q ),
    .c(_00461_),
    .y(_03076_)
  );
  al_ao21ftf _08340_ (
    .a(\DFF_609.Q ),
    .b(_03076_),
    .c(_01221_),
    .y(_03077_)
  );
  al_nand3 _08341_ (
    .a(g35),
    .b(_01222_),
    .c(_03077_),
    .y(_03078_)
  );
  al_ao21ftf _08342_ (
    .a(_03076_),
    .b(_01222_),
    .c(g35),
    .y(_03079_)
  );
  al_aoi21ftf _08343_ (
    .a(\DFF_254.Q ),
    .b(_03079_),
    .c(_03078_),
    .y(\DFF_609.D )
  );
  al_ao21ftf _08344_ (
    .a(g35),
    .b(\DFF_555.Q ),
    .c(_00494_),
    .y(\DFF_708.D )
  );
  al_or3 _08345_ (
    .a(\DFF_221.Q ),
    .b(g73),
    .c(g72),
    .y(_03080_)
  );
  al_mux2l _08346_ (
    .a(_03080_),
    .b(\DFF_384.Q ),
    .s(_01208_),
    .y(\DFF_1296.D )
  );
  al_and2 _08347_ (
    .a(\DFF_271.Q ),
    .b(g35),
    .y(\DFF_317.D )
  );
  al_nor2 _08348_ (
    .a(\DFF_432.Q ),
    .b(g35),
    .y(_03081_)
  );
  al_nor3ftt _08349_ (
    .a(\DFF_1192.Q ),
    .b(_01086_),
    .c(_01089_),
    .y(_03082_)
  );
  al_nand3 _08350_ (
    .a(_03082_),
    .b(_01100_),
    .c(_01096_),
    .y(_03083_)
  );
  al_oai21ttf _08351_ (
    .a(_01086_),
    .b(_01089_),
    .c(\DFF_1192.Q ),
    .y(_03084_)
  );
  al_and2 _08352_ (
    .a(g35),
    .b(_03084_),
    .y(_03085_)
  );
  al_aoi21 _08353_ (
    .a(_03085_),
    .b(_03083_),
    .c(_03081_),
    .y(\DFF_1192.D )
  );
  al_and2 _08354_ (
    .a(g35),
    .b(\DFF_1157.Q ),
    .y(\DFF_1157.D )
  );
  al_mux2l _08355_ (
    .a(\DFF_652.Q ),
    .b(\DFF_10.Q ),
    .s(_01109_),
    .y(\DFF_10.D )
  );
  al_oa21ftt _08356_ (
    .a(g35),
    .b(\DFF_969.Q ),
    .c(\DFF_1183.Q ),
    .y(_03086_)
  );
  al_aoi21ftf _08357_ (
    .a(\DFF_1062.Q ),
    .b(g35),
    .c(_03086_),
    .y(_03087_)
  );
  al_or3fft _08358_ (
    .a(\DFF_266.Q ),
    .b(g35),
    .c(_03087_),
    .y(_03088_)
  );
  al_aoi21ftf _08359_ (
    .a(_00066_),
    .b(\DFF_266.Q ),
    .c(_03087_),
    .y(_03089_)
  );
  al_nand2ft _08360_ (
    .a(_03089_),
    .b(_03088_),
    .y(\DFF_266.D )
  );
  al_and2ft _08361_ (
    .a(g35),
    .b(\DFF_1252.Q ),
    .y(_03090_)
  );
  al_nand3 _08362_ (
    .a(_00587_),
    .b(_01689_),
    .c(_00406_),
    .y(_03091_)
  );
  al_nand2ft _08363_ (
    .a(_00407_),
    .b(_01689_),
    .y(_03092_)
  );
  al_ao21 _08364_ (
    .a(\DFF_1252.Q ),
    .b(_01689_),
    .c(\DFF_1283.Q ),
    .y(_03093_)
  );
  al_and3 _08365_ (
    .a(g35),
    .b(_03092_),
    .c(_03093_),
    .y(_03094_)
  );
  al_ao21 _08366_ (
    .a(_03094_),
    .b(_03091_),
    .c(_03090_),
    .y(\DFF_1283.D )
  );
  al_oa21 _08367_ (
    .a(\DFF_956.Q ),
    .b(\DFF_593.Q ),
    .c(g35),
    .y(\DFF_593.D )
  );
  al_ao21 _08368_ (
    .a(\DFF_893.Q ),
    .b(\DFF_962.Q ),
    .c(\DFF_746.Q ),
    .y(_03095_)
  );
  al_nand3fft _08369_ (
    .a(_01963_),
    .b(_01964_),
    .c(_03095_),
    .y(_03096_)
  );
  al_ao21ftf _08370_ (
    .a(g35),
    .b(\DFF_893.Q ),
    .c(_03096_),
    .y(\DFF_746.D )
  );
  al_mux2h _08371_ (
    .a(\DFF_183.Q ),
    .b(_01934_),
    .s(_00358_),
    .y(_03097_)
  );
  al_mux2h _08372_ (
    .a(\DFF_336.Q ),
    .b(_03097_),
    .s(g35),
    .y(\DFF_183.D )
  );
  al_mux2l _08373_ (
    .a(\DFF_42.Q ),
    .b(\DFF_912.Q ),
    .s(_01127_),
    .y(\DFF_912.D )
  );
  al_nand2 _08374_ (
    .a(\DFF_1370.Q ),
    .b(\DFF_145.Q ),
    .y(_03098_)
  );
  al_nor2 _08375_ (
    .a(\DFF_1370.Q ),
    .b(\DFF_145.Q ),
    .y(_03099_)
  );
  al_nand2ft _08376_ (
    .a(_03099_),
    .b(_03098_),
    .y(_03100_)
  );
  al_mux2l _08377_ (
    .a(\DFF_456.Q ),
    .b(_03100_),
    .s(_01651_),
    .y(_03101_)
  );
  al_mux2h _08378_ (
    .a(\DFF_145.Q ),
    .b(_03101_),
    .s(g35),
    .y(\DFF_456.D )
  );
  al_nor3ftt _08379_ (
    .a(\DFF_136.Q ),
    .b(_00499_),
    .c(_00376_),
    .y(_03102_)
  );
  al_oa21ftt _08380_ (
    .a(\DFF_136.Q ),
    .b(_00376_),
    .c(_00499_),
    .y(_03103_)
  );
  al_nor3ftt _08381_ (
    .a(g35),
    .b(_03102_),
    .c(_03103_),
    .y(\DFF_136.D )
  );
  al_nand3 _08382_ (
    .a(_00499_),
    .b(_00691_),
    .c(_02707_),
    .y(_03104_)
  );
  al_ao21 _08383_ (
    .a(_02707_),
    .b(_00691_),
    .c(\DFF_479.Q ),
    .y(_03105_)
  );
  al_nand3 _08384_ (
    .a(g35),
    .b(_03105_),
    .c(_03104_),
    .y(_03106_)
  );
  al_ao21ftf _08385_ (
    .a(g35),
    .b(\DFF_340.Q ),
    .c(_03106_),
    .y(\DFF_479.D )
  );
  al_nor2 _08386_ (
    .a(g35),
    .b(\DFF_1164.Q ),
    .y(_03107_)
  );
  al_nor2ft _08387_ (
    .a(\DFF_669.Q ),
    .b(_01582_),
    .y(_03108_)
  );
  al_ao21ttf _08388_ (
    .a(_01826_),
    .b(_00920_),
    .c(_03108_),
    .y(_03109_)
  );
  al_mux2l _08389_ (
    .a(\DFF_736.Q ),
    .b(\DFF_669.Q ),
    .s(\DFF_799.Q ),
    .y(_03110_)
  );
  al_nor2ft _08390_ (
    .a(g35),
    .b(_03110_),
    .y(_03111_)
  );
  al_aoi21 _08391_ (
    .a(_03111_),
    .b(_03109_),
    .c(_03107_),
    .y(\DFF_736.D )
  );
  al_and2 _08392_ (
    .a(g35),
    .b(_02804_),
    .y(_03112_)
  );
  al_oai21 _08393_ (
    .a(_01169_),
    .b(_01344_),
    .c(_03112_),
    .y(_03113_)
  );
  al_ao21ftf _08394_ (
    .a(g35),
    .b(\DFF_925.Q ),
    .c(_03113_),
    .y(\DFF_653.D )
  );
  al_and3ftt _08395_ (
    .a(\DFF_893.Q ),
    .b(\DFF_1288.Q ),
    .c(\DFF_962.Q ),
    .y(_03114_)
  );
  al_aoi21 _08396_ (
    .a(\DFF_319.Q ),
    .b(_00561_),
    .c(_03114_),
    .y(_03115_)
  );
  al_and3 _08397_ (
    .a(\DFF_931.Q ),
    .b(\DFF_893.Q ),
    .c(\DFF_962.Q ),
    .y(_03116_)
  );
  al_aoi21 _08398_ (
    .a(\DFF_1.Q ),
    .b(_00575_),
    .c(_03116_),
    .y(_03117_)
  );
  al_ao21ttf _08399_ (
    .a(_03115_),
    .b(_03117_),
    .c(_01732_),
    .y(_03118_)
  );
  al_nand3ftt _08400_ (
    .a(\DFF_1310.Q ),
    .b(\DFF_893.Q ),
    .c(\DFF_962.Q ),
    .y(_03119_)
  );
  al_aoi21ftf _08401_ (
    .a(\DFF_772.Q ),
    .b(_00561_),
    .c(_03119_),
    .y(_03120_)
  );
  al_or3ftt _08402_ (
    .a(\DFF_962.Q ),
    .b(\DFF_893.Q ),
    .c(\DFF_1167.Q ),
    .y(_03121_)
  );
  al_aoi21ftf _08403_ (
    .a(\DFF_1069.Q ),
    .b(_00575_),
    .c(_03121_),
    .y(_03122_)
  );
  al_ao21 _08404_ (
    .a(_03120_),
    .b(_03122_),
    .c(_01732_),
    .y(_03123_)
  );
  al_nand3 _08405_ (
    .a(g35),
    .b(_03118_),
    .c(_03123_),
    .y(_03124_)
  );
  al_ao21ftf _08406_ (
    .a(g35),
    .b(\DFF_865.Q ),
    .c(_03124_),
    .y(\DFF_1033.D )
  );
  al_and2 _08407_ (
    .a(\DFF_1371.Q ),
    .b(\DFF_372.Q ),
    .y(_03125_)
  );
  al_aoi21 _08408_ (
    .a(\DFF_1371.Q ),
    .b(g35),
    .c(\DFF_372.Q ),
    .y(_03126_)
  );
  al_aoi21 _08409_ (
    .a(g35),
    .b(_03125_),
    .c(_03126_),
    .y(\DFF_1371.D )
  );
  al_nand3fft _08410_ (
    .a(_00066_),
    .b(\DFF_66.Q ),
    .c(_01696_),
    .y(_03127_)
  );
  al_aoi21ftf _08411_ (
    .a(\DFF_1419.Q ),
    .b(_00066_),
    .c(_03127_),
    .y(_03128_)
  );
  al_aoi21ftf _08412_ (
    .a(_00066_),
    .b(_02894_),
    .c(_03128_),
    .y(\DFF_66.D )
  );
  al_ao21 _08413_ (
    .a(\DFF_1080.Q ),
    .b(_01965_),
    .c(\DFF_1020.Q ),
    .y(_03129_)
  );
  al_and2ft _08414_ (
    .a(g35),
    .b(\DFF_1080.Q ),
    .y(_03130_)
  );
  al_ao21 _08415_ (
    .a(_03129_),
    .b(_01966_),
    .c(_03130_),
    .y(\DFF_1020.D )
  );
  al_aoi21 _08416_ (
    .a(\DFF_1080.Q ),
    .b(_01965_),
    .c(_01963_),
    .y(_03131_)
  );
  al_ao21ftf _08417_ (
    .a(_01965_),
    .b(_00427_),
    .c(_03131_),
    .y(_03132_)
  );
  al_ao21ftf _08418_ (
    .a(g35),
    .b(\DFF_1364.Q ),
    .c(_03132_),
    .y(\DFF_1080.D )
  );
  al_mux2l _08419_ (
    .a(\DFF_1357.Q ),
    .b(\DFF_608.Q ),
    .s(g35),
    .y(\DFF_1357.D )
  );
  al_or2 _08420_ (
    .a(\DFF_875.Q ),
    .b(_00369_),
    .y(_03133_)
  );
  al_nand2 _08421_ (
    .a(\DFF_875.Q ),
    .b(_00369_),
    .y(_03134_)
  );
  al_ao21 _08422_ (
    .a(_03134_),
    .b(_03133_),
    .c(_00066_),
    .y(_03135_)
  );
  al_aoi21ftf _08423_ (
    .a(\DFF_1021.Q ),
    .b(_00066_),
    .c(_03135_),
    .y(\DFF_875.D )
  );
  al_nand3 _08424_ (
    .a(_00499_),
    .b(_02624_),
    .c(_01169_),
    .y(_03136_)
  );
  al_ao21 _08425_ (
    .a(_01169_),
    .b(_02624_),
    .c(\DFF_82.Q ),
    .y(_03137_)
  );
  al_nand3 _08426_ (
    .a(g35),
    .b(_03137_),
    .c(_03136_),
    .y(_03138_)
  );
  al_ao21ftf _08427_ (
    .a(g35),
    .b(\DFF_483.Q ),
    .c(_03138_),
    .y(\DFF_82.D )
  );
  al_oa21ftt _08428_ (
    .a(g35),
    .b(\DFF_787.Q ),
    .c(\DFF_1367.Q ),
    .y(\DFF_668.D )
  );
  al_and2ft _08429_ (
    .a(g35),
    .b(\DFF_874.Q ),
    .y(_03139_)
  );
  al_ao21ftt _08430_ (
    .a(_00226_),
    .b(_01183_),
    .c(_02430_),
    .y(_03140_)
  );
  al_aoi21 _08431_ (
    .a(\DFF_966.Q ),
    .b(_02430_),
    .c(_00066_),
    .y(_03141_)
  );
  al_ao21 _08432_ (
    .a(_03140_),
    .b(_03141_),
    .c(_03139_),
    .y(\DFF_966.D )
  );
  al_nand3ftt _08433_ (
    .a(_01311_),
    .b(_00499_),
    .c(_01952_),
    .y(_03142_)
  );
  al_ao21ftt _08434_ (
    .a(_01311_),
    .b(_01952_),
    .c(\DFF_390.Q ),
    .y(_03143_)
  );
  al_nand3 _08435_ (
    .a(g35),
    .b(_03142_),
    .c(_03143_),
    .y(_03144_)
  );
  al_ao21ftf _08436_ (
    .a(g35),
    .b(\DFF_1040.Q ),
    .c(_03144_),
    .y(\DFF_390.D )
  );
  al_ao21 _08437_ (
    .a(\DFF_270.Q ),
    .b(g35),
    .c(\DFF_635.Q ),
    .y(_03145_)
  );
  al_nand3 _08438_ (
    .a(\DFF_635.Q ),
    .b(\DFF_270.Q ),
    .c(g35),
    .y(_03146_)
  );
  al_nand2 _08439_ (
    .a(_03145_),
    .b(_03146_),
    .y(_03147_)
  );
  al_oa21ftf _08440_ (
    .a(g35),
    .b(_00745_),
    .c(_03147_),
    .y(\DFF_270.D )
  );
  al_and2ft _08441_ (
    .a(g35),
    .b(\DFF_894.Q ),
    .y(_03148_)
  );
  al_or2 _08442_ (
    .a(\DFF_849.Q ),
    .b(_03010_),
    .y(_03149_)
  );
  al_aoi21ftf _08443_ (
    .a(_01224_),
    .b(_01324_),
    .c(_03149_),
    .y(_03150_)
  );
  al_ao21 _08444_ (
    .a(_03150_),
    .b(_01319_),
    .c(_03148_),
    .y(\DFF_849.D )
  );
  al_aoi21 _08445_ (
    .a(\DFF_1261.Q ),
    .b(_01195_),
    .c(_00066_),
    .y(_03151_)
  );
  al_oai21 _08446_ (
    .a(\DFF_1261.Q ),
    .b(_01195_),
    .c(_03151_),
    .y(_03152_)
  );
  al_aoi21ftf _08447_ (
    .a(\DFF_322.Q ),
    .b(_00066_),
    .c(_03152_),
    .y(\DFF_1261.D )
  );
  al_oai21 _08448_ (
    .a(_01409_),
    .b(_01976_),
    .c(_01496_),
    .y(_03153_)
  );
  al_ao21ftf _08449_ (
    .a(g35),
    .b(\DFF_407.Q ),
    .c(_03153_),
    .y(\DFF_1304.D )
  );
  al_oa21ttf _08450_ (
    .a(\DFF_329.Q ),
    .b(\DFF_396.Q ),
    .c(\DFF_426.Q ),
    .y(_03154_)
  );
  al_nand3 _08451_ (
    .a(_03154_),
    .b(_02004_),
    .c(_02006_),
    .y(_03155_)
  );
  al_or3ftt _08452_ (
    .a(\DFF_426.Q ),
    .b(\DFF_329.Q ),
    .c(\DFF_396.Q ),
    .y(_03156_)
  );
  al_nand3 _08453_ (
    .a(g35),
    .b(_03156_),
    .c(_03155_),
    .y(_03157_)
  );
  al_aoi21ftf _08454_ (
    .a(\DFF_329.Q ),
    .b(_00066_),
    .c(_03157_),
    .y(\DFF_426.D )
  );
  al_nor3fft _08455_ (
    .a(\DFF_591.Q ),
    .b(g35),
    .c(_01348_),
    .y(_03158_)
  );
  al_ao21 _08456_ (
    .a(\DFF_447.Q ),
    .b(_01351_),
    .c(_03158_),
    .y(\DFF_591.D )
  );
  al_mux2l _08457_ (
    .a(\DFF_141.Q ),
    .b(\DFF_1065.Q ),
    .s(g35),
    .y(\DFF_545.D )
  );
  al_nor2 _08458_ (
    .a(\DFF_639.Q ),
    .b(g35),
    .y(_03159_)
  );
  al_mux2l _08459_ (
    .a(_01874_),
    .b(_01871_),
    .s(_01869_),
    .y(_03160_)
  );
  al_or3fft _08460_ (
    .a(\DFF_1238.Q ),
    .b(_02565_),
    .c(_03160_),
    .y(_03161_)
  );
  al_aoi21ftf _08461_ (
    .a(\DFF_1238.Q ),
    .b(_03160_),
    .c(g35),
    .y(_03162_)
  );
  al_aoi21 _08462_ (
    .a(_03161_),
    .b(_03162_),
    .c(_03159_),
    .y(\DFF_1238.D )
  );
  al_mux2l _08463_ (
    .a(\DFF_1275.Q ),
    .b(\DFF_1072.Q ),
    .s(\DFF_1110.Q ),
    .y(_03163_)
  );
  al_mux2h _08464_ (
    .a(\DFF_395.Q ),
    .b(_03163_),
    .s(g35),
    .y(\DFF_1072.D )
  );
  al_or2 _08465_ (
    .a(_01534_),
    .b(_00974_),
    .y(_03164_)
  );
  al_and3ftt _08466_ (
    .a(_00975_),
    .b(_01535_),
    .c(_00974_),
    .y(_03165_)
  );
  al_nand2 _08467_ (
    .a(_03165_),
    .b(_02883_),
    .y(_03166_)
  );
  al_aoi21 _08468_ (
    .a(_03164_),
    .b(_03166_),
    .c(_00066_),
    .y(\DFF_1143.D )
  );
  al_nand3fft _08469_ (
    .a(\DFF_42.Q ),
    .b(_00066_),
    .c(_02776_),
    .y(_03167_)
  );
  al_or3fft _08470_ (
    .a(\DFF_42.Q ),
    .b(g35),
    .c(_02776_),
    .y(_03168_)
  );
  al_or2 _08471_ (
    .a(g35),
    .b(\DFF_1216.Q ),
    .y(_03169_)
  );
  al_and3 _08472_ (
    .a(_03169_),
    .b(_03167_),
    .c(_03168_),
    .y(\DFF_42.D )
  );
  al_and2 _08473_ (
    .a(\DFF_538.Q ),
    .b(g35),
    .y(_03170_)
  );
  al_aoi21ttf _08474_ (
    .a(_03170_),
    .b(_00714_),
    .c(\DFF_224.Q ),
    .y(\DFF_840.D )
  );
  al_nand3 _08475_ (
    .a(_00499_),
    .b(_02367_),
    .c(_01266_),
    .y(_03171_)
  );
  al_ao21 _08476_ (
    .a(_01266_),
    .b(_02367_),
    .c(\DFF_1013.Q ),
    .y(_03172_)
  );
  al_nand3 _08477_ (
    .a(g35),
    .b(_03172_),
    .c(_03171_),
    .y(_03173_)
  );
  al_ao21ftf _08478_ (
    .a(g35),
    .b(\DFF_917.Q ),
    .c(_03173_),
    .y(\DFF_1013.D )
  );
  al_aoi21ttf _08479_ (
    .a(\DFF_73.Q ),
    .b(g35),
    .c(\DFF_1190.Q ),
    .y(_03174_)
  );
  al_ao21 _08480_ (
    .a(\DFF_73.Q ),
    .b(\DFF_1190.D ),
    .c(_03174_),
    .y(\DFF_73.D )
  );
  al_and3 _08481_ (
    .a(_00695_),
    .b(\DFF_746.Q ),
    .c(_00549_),
    .y(_03175_)
  );
  al_aoi21ftf _08482_ (
    .a(g113),
    .b(_00342_),
    .c(\DFF_470.Q ),
    .y(_03176_)
  );
  al_nand3fft _08483_ (
    .a(_00698_),
    .b(_03176_),
    .c(_03175_),
    .y(_03177_)
  );
  al_ao21ftf _08484_ (
    .a(_03175_),
    .b(\DFF_284.Q ),
    .c(_03177_),
    .y(_03178_)
  );
  al_mux2h _08485_ (
    .a(\DFF_302.Q ),
    .b(_03178_),
    .s(g35),
    .y(\DFF_284.D )
  );
  al_aoi21ttf _08486_ (
    .a(_00577_),
    .b(_00430_),
    .c(_02775_),
    .y(_03179_)
  );
  al_oa21ttf _08487_ (
    .a(\DFF_103.Q ),
    .b(_02922_),
    .c(_00066_),
    .y(_03180_)
  );
  al_inv _08488_ (
    .a(\DFF_1202.Q ),
    .y(_03181_)
  );
  al_or3ftt _08489_ (
    .a(g35),
    .b(\DFF_705.Q ),
    .c(_02775_),
    .y(_03182_)
  );
  al_ao21ftf _08490_ (
    .a(g35),
    .b(_03181_),
    .c(_03182_),
    .y(_03183_)
  );
  al_aoi21 _08491_ (
    .a(_03180_),
    .b(_03179_),
    .c(_03183_),
    .y(\DFF_705.D )
  );
  al_and3ftt _08492_ (
    .a(\DFF_793.Q ),
    .b(\DFF_1025.Q ),
    .c(\DFF_1331.Q ),
    .y(_03184_)
  );
  al_and3ftt _08493_ (
    .a(\DFF_793.Q ),
    .b(\DFF_148.Q ),
    .c(\DFF_887.Q ),
    .y(_03185_)
  );
  al_ao21 _08494_ (
    .a(\DFF_959.Q ),
    .b(_00441_),
    .c(_03185_),
    .y(_03186_)
  );
  al_and3ftt _08495_ (
    .a(\DFF_1331.Q ),
    .b(\DFF_793.Q ),
    .c(\DFF_930.Q ),
    .y(_03187_)
  );
  al_and3fft _08496_ (
    .a(\DFF_1331.Q ),
    .b(\DFF_148.Q ),
    .c(\DFF_1171.Q ),
    .y(_03188_)
  );
  al_nand3 _08497_ (
    .a(\DFF_273.Q ),
    .b(\DFF_1331.Q ),
    .c(\DFF_148.Q ),
    .y(_03189_)
  );
  al_and3fft _08498_ (
    .a(_03187_),
    .b(_03188_),
    .c(_03189_),
    .y(_03190_)
  );
  al_nand3fft _08499_ (
    .a(_03184_),
    .b(_03186_),
    .c(_03190_),
    .y(_03191_)
  );
  al_mux2l _08500_ (
    .a(_03191_),
    .b(\DFF_989.Q ),
    .s(_00563_),
    .y(_03192_)
  );
  al_mux2h _08501_ (
    .a(\DFF_148.Q ),
    .b(_03192_),
    .s(g35),
    .y(\DFF_989.D )
  );
  al_and2ft _08502_ (
    .a(\DFF_1354.Q ),
    .b(\DFF_1155.Q ),
    .y(_03193_)
  );
  al_oai21ttf _08503_ (
    .a(\DFF_529.Q ),
    .b(\DFF_1038.Q ),
    .c(_00713_),
    .y(_03194_)
  );
  al_or2 _08504_ (
    .a(\DFF_1293.Q ),
    .b(\DFF_1354.Q ),
    .y(_03195_)
  );
  al_ao21ttf _08505_ (
    .a(\DFF_1293.Q ),
    .b(\DFF_1038.Q ),
    .c(_03195_),
    .y(_03196_)
  );
  al_and3ftt _08506_ (
    .a(_03193_),
    .b(_03196_),
    .c(_03194_),
    .y(_03197_)
  );
  al_and3ftt _08507_ (
    .a(_00714_),
    .b(g35),
    .c(_03197_),
    .y(\DFF_819.D )
  );
  al_nand3 _08508_ (
    .a(_00499_),
    .b(_02367_),
    .c(_00596_),
    .y(_03198_)
  );
  al_ao21 _08509_ (
    .a(_02367_),
    .b(_00596_),
    .c(\DFF_414.Q ),
    .y(_03199_)
  );
  al_nand3 _08510_ (
    .a(g35),
    .b(_03198_),
    .c(_03199_),
    .y(_03200_)
  );
  al_ao21ftf _08511_ (
    .a(g35),
    .b(\DFF_1013.Q ),
    .c(_03200_),
    .y(\DFF_414.D )
  );
  al_nand3 _08512_ (
    .a(_00499_),
    .b(_00567_),
    .c(_01840_),
    .y(_03201_)
  );
  al_ao21 _08513_ (
    .a(_01840_),
    .b(_00567_),
    .c(\DFF_659.Q ),
    .y(_03202_)
  );
  al_nand3 _08514_ (
    .a(g35),
    .b(_03202_),
    .c(_03201_),
    .y(_03203_)
  );
  al_ao21ftf _08515_ (
    .a(g35),
    .b(\DFF_773.Q ),
    .c(_03203_),
    .y(\DFF_659.D )
  );
  al_mux2l _08516_ (
    .a(\DFF_767.Q ),
    .b(\DFF_673.Q ),
    .s(g35),
    .y(\DFF_767.D )
  );
  al_or2 _08517_ (
    .a(\DFF_358.Q ),
    .b(_00603_),
    .y(_03204_)
  );
  al_nand3ftt _08518_ (
    .a(_02226_),
    .b(_01505_),
    .c(_03204_),
    .y(_03205_)
  );
  al_ao21ftf _08519_ (
    .a(g35),
    .b(\DFF_115.Q ),
    .c(_03205_),
    .y(\DFF_358.D )
  );
  al_mux2l _08520_ (
    .a(\DFF_673.Q ),
    .b(\DFF_1000.Q ),
    .s(g35),
    .y(\DFF_673.D )
  );
  al_inv _08521_ (
    .a(\DFF_21.Q ),
    .y(_03206_)
  );
  al_nand3fft _08522_ (
    .a(_03206_),
    .b(_00940_),
    .c(_00954_),
    .y(_03207_)
  );
  al_ao21 _08523_ (
    .a(_00278_),
    .b(_03207_),
    .c(_01837_),
    .y(_03208_)
  );
  al_ao21ftf _08524_ (
    .a(g35),
    .b(\DFF_21.Q ),
    .c(_03208_),
    .y(\DFF_142.D )
  );
  al_mux2h _08525_ (
    .a(\DFF_1272.Q ),
    .b(_00982_),
    .s(g35),
    .y(\DFF_980.D )
  );
  al_aoi21 _08526_ (
    .a(\DFF_1243.Q ),
    .b(_00547_),
    .c(_00066_),
    .y(_03209_)
  );
  al_oai21 _08527_ (
    .a(\DFF_1243.Q ),
    .b(_00547_),
    .c(_03209_),
    .y(_03210_)
  );
  al_aoi21ftf _08528_ (
    .a(g35),
    .b(_01486_),
    .c(_03210_),
    .y(\DFF_1243.D )
  );
  al_nor2 _08529_ (
    .a(\DFF_1105.Q ),
    .b(g35),
    .y(_03211_)
  );
  al_or2 _08530_ (
    .a(\DFF_1105.Q ),
    .b(_01682_),
    .y(_03212_)
  );
  al_aoi21ftf _08531_ (
    .a(_01681_),
    .b(_01679_),
    .c(_03212_),
    .y(_03213_)
  );
  al_nand3 _08532_ (
    .a(\DFF_940.Q ),
    .b(_01039_),
    .c(_03213_),
    .y(_03214_)
  );
  al_oa21ttf _08533_ (
    .a(\DFF_940.Q ),
    .b(_03213_),
    .c(_00066_),
    .y(_03215_)
  );
  al_aoi21 _08534_ (
    .a(_03214_),
    .b(_03215_),
    .c(_03211_),
    .y(\DFF_940.D )
  );
  al_and2ft _08535_ (
    .a(\DFF_1344.Q ),
    .b(g35),
    .y(_03216_)
  );
  al_or3fft _08536_ (
    .a(_02018_),
    .b(g35),
    .c(_01056_),
    .y(_03217_)
  );
  al_ao21ftf _08537_ (
    .a(\DFF_342.Q ),
    .b(_00066_),
    .c(_03217_),
    .y(_03218_)
  );
  al_aoi21 _08538_ (
    .a(_03216_),
    .b(_01058_),
    .c(_03218_),
    .y(\DFF_794.D )
  );
  al_ao21ttf _08539_ (
    .a(_02820_),
    .b(_00576_),
    .c(\DFF_232.Q ),
    .y(_03219_)
  );
  al_nand3ftt _08540_ (
    .a(\DFF_232.Q ),
    .b(_02820_),
    .c(_00576_),
    .y(_03220_)
  );
  al_nand3 _08541_ (
    .a(g35),
    .b(_03220_),
    .c(_03219_),
    .y(_03221_)
  );
  al_aoi21ftf _08542_ (
    .a(\DFF_301.Q ),
    .b(_00066_),
    .c(_03221_),
    .y(\DFF_232.D )
  );
  al_nand3 _08543_ (
    .a(\DFF_90.Q ),
    .b(\DFF_295.Q ),
    .c(\DFF_1057.Q ),
    .y(_03222_)
  );
  al_mux2l _08544_ (
    .a(\DFF_363.Q ),
    .b(_00344_),
    .s(_03222_),
    .y(_03223_)
  );
  al_mux2h _08545_ (
    .a(\DFF_1057.Q ),
    .b(_03223_),
    .s(g35),
    .y(\DFF_363.D )
  );
  al_oa21ftf _08546_ (
    .a(_01682_),
    .b(_01679_),
    .c(_01681_),
    .y(_03224_)
  );
  al_nand3 _08547_ (
    .a(\DFF_1105.Q ),
    .b(_01039_),
    .c(_01041_),
    .y(_03225_)
  );
  al_nand3ftt _08548_ (
    .a(_01679_),
    .b(_01682_),
    .c(_03225_),
    .y(_03226_)
  );
  al_nand3fft _08549_ (
    .a(_00066_),
    .b(_03224_),
    .c(_03226_),
    .y(_03227_)
  );
  al_ao21ftf _08550_ (
    .a(g35),
    .b(\DFF_850.Q ),
    .c(_03227_),
    .y(\DFF_1105.D )
  );
  al_oai21ftf _08551_ (
    .a(g35),
    .b(_01058_),
    .c(\DFF_1064.Q ),
    .y(_03228_)
  );
  al_aoi21ftf _08552_ (
    .a(\DFF_1344.Q ),
    .b(_01063_),
    .c(_03228_),
    .y(\DFF_1344.D )
  );
  al_mux2l _08553_ (
    .a(\DFF_1404.Q ),
    .b(\DFF_1162.Q ),
    .s(\DFF_1252.Q ),
    .y(_03229_)
  );
  al_aoi21 _08554_ (
    .a(\DFF_1283.Q ),
    .b(_03229_),
    .c(\DFF_254.Q ),
    .y(_03230_)
  );
  al_oai21 _08555_ (
    .a(\DFF_1283.Q ),
    .b(_03229_),
    .c(_03230_),
    .y(_03231_)
  );
  al_ao21ftf _08556_ (
    .a(_03076_),
    .b(_03231_),
    .c(_01689_),
    .y(_03232_)
  );
  al_or2 _08557_ (
    .a(\DFF_254.Q ),
    .b(_01689_),
    .y(_03233_)
  );
  al_and3 _08558_ (
    .a(g35),
    .b(_03232_),
    .c(_03233_),
    .y(\DFF_254.D )
  );
  al_and2ft _08559_ (
    .a(g35),
    .b(\DFF_176.Q ),
    .y(_03234_)
  );
  al_aoi21ftt _08560_ (
    .a(_01945_),
    .b(_01941_),
    .c(_02136_),
    .y(_03235_)
  );
  al_ao21ftf _08561_ (
    .a(_01944_),
    .b(_01940_),
    .c(_03235_),
    .y(_03236_)
  );
  al_ao21ftf _08562_ (
    .a(_01939_),
    .b(_01947_),
    .c(_03236_),
    .y(_03237_)
  );
  al_oa21ftf _08563_ (
    .a(\DFF_618.Q ),
    .b(_03236_),
    .c(_00066_),
    .y(_03238_)
  );
  al_ao21 _08564_ (
    .a(_03237_),
    .b(_03238_),
    .c(_03234_),
    .y(\DFF_618.D )
  );
  al_and2ft _08565_ (
    .a(g35),
    .b(\DFF_769.Q ),
    .y(_03239_)
  );
  al_and3ftt _08566_ (
    .a(_01281_),
    .b(_00604_),
    .c(_02638_),
    .y(_03240_)
  );
  al_oai21ftt _08567_ (
    .a(\DFF_1047.Q ),
    .b(\DFF_1141.Q ),
    .c(\DFF_1181.Q ),
    .y(_03241_)
  );
  al_or3ftt _08568_ (
    .a(\DFF_1047.Q ),
    .b(\DFF_1141.Q ),
    .c(\DFF_1181.Q ),
    .y(_03242_)
  );
  al_nand3 _08569_ (
    .a(_03241_),
    .b(_03242_),
    .c(_03240_),
    .y(_03243_)
  );
  al_oa21ttf _08570_ (
    .a(\DFF_658.Q ),
    .b(_03240_),
    .c(_00066_),
    .y(_03244_)
  );
  al_ao21 _08571_ (
    .a(_03243_),
    .b(_03244_),
    .c(_03239_),
    .y(\DFF_658.D )
  );
  al_nand2 _08572_ (
    .a(g35),
    .b(_03222_),
    .y(_03245_)
  );
  al_aoi21ttf _08573_ (
    .a(\DFF_1103.Q ),
    .b(g35),
    .c(\DFF_363.Q ),
    .y(_03246_)
  );
  al_mux2l _08574_ (
    .a(_03246_),
    .b(\DFF_1103.Q ),
    .s(_03245_),
    .y(\DFF_1103.D )
  );
  al_and2ft _08575_ (
    .a(g35),
    .b(\DFF_502.Q ),
    .y(_03247_)
  );
  al_ao21ftf _08576_ (
    .a(_01098_),
    .b(_01094_),
    .c(_01092_),
    .y(_03248_)
  );
  al_ao21ftf _08577_ (
    .a(_01093_),
    .b(_01100_),
    .c(_03248_),
    .y(_03249_)
  );
  al_oa21ftf _08578_ (
    .a(\DFF_0.Q ),
    .b(_03248_),
    .c(_00066_),
    .y(_03250_)
  );
  al_ao21 _08579_ (
    .a(_03249_),
    .b(_03250_),
    .c(_03247_),
    .y(\DFF_0.D )
  );
  al_nand3ftt _08580_ (
    .a(_03064_),
    .b(_00499_),
    .c(_02754_),
    .y(_03251_)
  );
  al_ao21ftt _08581_ (
    .a(_03064_),
    .b(_02754_),
    .c(\DFF_1378.Q ),
    .y(_03252_)
  );
  al_nand3 _08582_ (
    .a(g35),
    .b(_03251_),
    .c(_03252_),
    .y(_03253_)
  );
  al_ao21ftf _08583_ (
    .a(g35),
    .b(\DFF_271.Q ),
    .c(_03253_),
    .y(\DFF_1378.D )
  );
  al_nand2 _08584_ (
    .a(\DFF_1261.Q ),
    .b(\DFF_264.Q ),
    .y(_03254_)
  );
  al_nor2 _08585_ (
    .a(\DFF_1261.Q ),
    .b(\DFF_264.Q ),
    .y(_03255_)
  );
  al_nand2ft _08586_ (
    .a(_03255_),
    .b(_03254_),
    .y(_03256_)
  );
  al_mux2l _08587_ (
    .a(\DFF_1213.Q ),
    .b(_03256_),
    .s(_01364_),
    .y(_03257_)
  );
  al_mux2h _08588_ (
    .a(\DFF_264.Q ),
    .b(_03257_),
    .s(g35),
    .y(\DFF_1213.D )
  );
  al_mux2l _08589_ (
    .a(\DFF_1053.Q ),
    .b(\DFF_601.Q ),
    .s(_01174_),
    .y(\DFF_601.D )
  );
  al_aoi21 _08590_ (
    .a(\DFF_5.Q ),
    .b(_00882_),
    .c(_00066_),
    .y(_03258_)
  );
  al_nand2ft _08591_ (
    .a(g35),
    .b(\DFF_5.Q ),
    .y(_03259_)
  );
  al_ao21ftf _08592_ (
    .a(\DFF_347.Q ),
    .b(_03258_),
    .c(_03259_),
    .y(\DFF_423.D )
  );
  al_nand2ft _08593_ (
    .a(g35),
    .b(\DFF_956.Q ),
    .y(_03260_)
  );
  al_ao21ftf _08594_ (
    .a(\DFF_1061.Q ),
    .b(g35),
    .c(_03260_),
    .y(\DFF_612.D )
  );
  al_ao21 _08595_ (
    .a(\DFF_1183.Q ),
    .b(g35),
    .c(_01384_),
    .y(_03261_)
  );
  al_and3 _08596_ (
    .a(\DFF_1183.Q ),
    .b(g35),
    .c(_01384_),
    .y(_03262_)
  );
  al_and2ft _08597_ (
    .a(_03262_),
    .b(_03261_),
    .y(\DFF_1183.D )
  );
  al_nand3 _08598_ (
    .a(_00499_),
    .b(_01070_),
    .c(_02010_),
    .y(_03263_)
  );
  al_ao21 _08599_ (
    .a(_01070_),
    .b(_02010_),
    .c(\DFF_108.Q ),
    .y(_03264_)
  );
  al_nand3 _08600_ (
    .a(g35),
    .b(_03264_),
    .c(_03263_),
    .y(_03265_)
  );
  al_ao21ftf _08601_ (
    .a(g35),
    .b(\DFF_12.Q ),
    .c(_03265_),
    .y(\DFF_108.D )
  );
  al_nand3 _08602_ (
    .a(_00499_),
    .b(_01266_),
    .c(_02426_),
    .y(_03266_)
  );
  al_ao21 _08603_ (
    .a(_01266_),
    .b(_02426_),
    .c(\DFF_1160.Q ),
    .y(_03267_)
  );
  al_nand3 _08604_ (
    .a(g35),
    .b(_03267_),
    .c(_03266_),
    .y(_03268_)
  );
  al_ao21ftf _08605_ (
    .a(g35),
    .b(\DFF_986.Q ),
    .c(_03268_),
    .y(\DFF_1160.D )
  );
  al_and3 _08606_ (
    .a(\DFF_845.Q ),
    .b(_00696_),
    .c(_00549_),
    .y(_03269_)
  );
  al_aoi21ftf _08607_ (
    .a(g113),
    .b(_00342_),
    .c(\DFF_534.Q ),
    .y(_03270_)
  );
  al_nand3fft _08608_ (
    .a(_00698_),
    .b(_03270_),
    .c(_03269_),
    .y(_03271_)
  );
  al_ao21ftf _08609_ (
    .a(_03269_),
    .b(\DFF_302.Q ),
    .c(_03271_),
    .y(_03272_)
  );
  al_mux2h _08610_ (
    .a(\DFF_233.Q ),
    .b(_03272_),
    .s(g35),
    .y(\DFF_302.D )
  );
  al_oai21ttf _08611_ (
    .a(\DFF_806.Q ),
    .b(\DFF_1196.Q ),
    .c(_03027_),
    .y(_03273_)
  );
  al_nand2ft _08612_ (
    .a(\DFF_1185.Q ),
    .b(\DFF_163.Q ),
    .y(_03274_)
  );
  al_nand2ft _08613_ (
    .a(\DFF_1248.Q ),
    .b(\DFF_1185.Q ),
    .y(_03275_)
  );
  al_aoi21ftf _08614_ (
    .a(\DFF_1196.Q ),
    .b(\DFF_1248.Q ),
    .c(_03275_),
    .y(_03276_)
  );
  al_and3 _08615_ (
    .a(g35),
    .b(_03274_),
    .c(_03276_),
    .y(_03277_)
  );
  al_and3ftt _08616_ (
    .a(_03028_),
    .b(_03273_),
    .c(_03277_),
    .y(\DFF_1158.D )
  );
  al_mux2l _08617_ (
    .a(\DFF_771.Q ),
    .b(\DFF_561.Q ),
    .s(_01557_),
    .y(_03278_)
  );
  al_mux2h _08618_ (
    .a(\DFF_382.Q ),
    .b(_03278_),
    .s(g35),
    .y(\DFF_771.D )
  );
  al_oai21ftt _08619_ (
    .a(g35),
    .b(_01425_),
    .c(\DFF_692.Q ),
    .y(_03279_)
  );
  al_ao21ftf _08620_ (
    .a(_00066_),
    .b(\DFF_687.Q ),
    .c(_03279_),
    .y(\DFF_490.D )
  );
  al_and3ftt _08621_ (
    .a(\DFF_331.Q ),
    .b(_01406_),
    .c(_01505_),
    .y(\DFF_331.D )
  );
  al_nand3ftt _08622_ (
    .a(\DFF_916.Q ),
    .b(\DFF_20.Q ),
    .c(\DFF_104.Q ),
    .y(_03280_)
  );
  al_aoi21ftf _08623_ (
    .a(\DFF_314.Q ),
    .b(_03280_),
    .c(g35),
    .y(_03281_)
  );
  al_ao21ftf _08624_ (
    .a(_03280_),
    .b(_00499_),
    .c(_03281_),
    .y(_03282_)
  );
  al_ao21ftf _08625_ (
    .a(g35),
    .b(\DFF_1307.Q ),
    .c(_03282_),
    .y(\DFF_314.D )
  );
  al_nand3ftt _08626_ (
    .a(\DFF_843.Q ),
    .b(\DFF_126.Q ),
    .c(g35),
    .y(_03283_)
  );
  al_ao21ftf _08627_ (
    .a(g35),
    .b(\DFF_448.Q ),
    .c(_03283_),
    .y(\DFF_843.D )
  );
  al_nor2 _08628_ (
    .a(\DFF_217.Q ),
    .b(g35),
    .y(_03284_)
  );
  al_mux2h _08629_ (
    .a(_01447_),
    .b(_01450_),
    .s(\DFF_217.Q ),
    .y(_03285_)
  );
  al_nand3ftt _08630_ (
    .a(_03285_),
    .b(\DFF_1170.Q ),
    .c(_01455_),
    .y(_03286_)
  );
  al_aoi21ftf _08631_ (
    .a(\DFF_1170.Q ),
    .b(_03285_),
    .c(g35),
    .y(_03287_)
  );
  al_aoi21 _08632_ (
    .a(_03287_),
    .b(_03286_),
    .c(_03284_),
    .y(\DFF_1170.D )
  );
  al_nand2 _08633_ (
    .a(\DFF_1034.Q ),
    .b(\DFF_1276.Q ),
    .y(_03288_)
  );
  al_nor2 _08634_ (
    .a(\DFF_1034.Q ),
    .b(\DFF_1276.Q ),
    .y(_03289_)
  );
  al_nand2ft _08635_ (
    .a(_03289_),
    .b(_03288_),
    .y(_03290_)
  );
  al_mux2l _08636_ (
    .a(\DFF_499.Q ),
    .b(_03290_),
    .s(_01437_),
    .y(_03291_)
  );
  al_mux2h _08637_ (
    .a(\DFF_1276.Q ),
    .b(_03291_),
    .s(g35),
    .y(\DFF_499.D )
  );
  al_nand3 _08638_ (
    .a(_01028_),
    .b(_01046_),
    .c(_01014_),
    .y(_03292_)
  );
  al_ao21ftf _08639_ (
    .a(g35),
    .b(\DFF_27.Q ),
    .c(_03292_),
    .y(\DFF_245.D )
  );
  al_and2ft _08640_ (
    .a(g35),
    .b(\DFF_1077.Q ),
    .y(_03293_)
  );
  al_oai21 _08641_ (
    .a(\DFF_1077.Q ),
    .b(_01632_),
    .c(_01630_),
    .y(_03294_)
  );
  al_ao21ttf _08642_ (
    .a(\DFF_335.Q ),
    .b(_01642_),
    .c(_03294_),
    .y(_03295_)
  );
  al_oa21ftf _08643_ (
    .a(\DFF_335.Q ),
    .b(_03294_),
    .c(_00066_),
    .y(_03296_)
  );
  al_ao21 _08644_ (
    .a(_03296_),
    .b(_03295_),
    .c(_03293_),
    .y(\DFF_335.D )
  );
  al_nand3ftt _08645_ (
    .a(\DFF_1150.Q ),
    .b(\DFF_1273.Q ),
    .c(\DFF_1068.Q ),
    .y(_03297_)
  );
  al_aoi21ftf _08646_ (
    .a(\DFF_1024.Q ),
    .b(_03297_),
    .c(g35),
    .y(_03298_)
  );
  al_ao21ftf _08647_ (
    .a(_03297_),
    .b(_00499_),
    .c(_03298_),
    .y(_03299_)
  );
  al_ao21ftf _08648_ (
    .a(g35),
    .b(\DFF_378.Q ),
    .c(_03299_),
    .y(\DFF_1024.D )
  );
  al_and2 _08649_ (
    .a(\DFF_75.Q ),
    .b(g35),
    .y(\DFF_75.D )
  );
  al_or2 _08650_ (
    .a(_01885_),
    .b(_01889_),
    .y(_03300_)
  );
  al_and3ftt _08651_ (
    .a(_01575_),
    .b(_01884_),
    .c(_01889_),
    .y(_03301_)
  );
  al_nand2 _08652_ (
    .a(_03301_),
    .b(_03061_),
    .y(_03302_)
  );
  al_aoi21 _08653_ (
    .a(_03300_),
    .b(_03302_),
    .c(_00066_),
    .y(\DFF_272.D )
  );
  al_and2ft _08654_ (
    .a(g35),
    .b(\DFF_570.Q ),
    .y(_03303_)
  );
  al_inv _08655_ (
    .a(\DFF_1091.Q ),
    .y(_03304_)
  );
  al_ao21ftf _08656_ (
    .a(_00855_),
    .b(_03304_),
    .c(_00578_),
    .y(_03305_)
  );
  al_oa21ftf _08657_ (
    .a(_00574_),
    .b(_00576_),
    .c(_00066_),
    .y(_03306_)
  );
  al_ao21 _08658_ (
    .a(_03306_),
    .b(_03305_),
    .c(_03303_),
    .y(\DFF_993.D )
  );
  al_aoi21 _08659_ (
    .a(\DFF_88.Q ),
    .b(_01184_),
    .c(\DFF_728.Q ),
    .y(_03307_)
  );
  al_or3ftt _08660_ (
    .a(_02276_),
    .b(_01185_),
    .c(_03307_),
    .y(_03308_)
  );
  al_ao21ftf _08661_ (
    .a(g35),
    .b(\DFF_88.Q ),
    .c(_03308_),
    .y(\DFF_728.D )
  );
  al_nand3 _08662_ (
    .a(_00499_),
    .b(_01046_),
    .c(_02011_),
    .y(_03309_)
  );
  al_ao21 _08663_ (
    .a(_02011_),
    .b(_01046_),
    .c(\DFF_72.Q ),
    .y(_03310_)
  );
  al_nand3 _08664_ (
    .a(g35),
    .b(_03310_),
    .c(_03309_),
    .y(_03311_)
  );
  al_ao21ftf _08665_ (
    .a(g35),
    .b(\DFF_633.Q ),
    .c(_03311_),
    .y(\DFF_72.D )
  );
  al_nand2 _08666_ (
    .a(g35),
    .b(_01364_),
    .y(_03312_)
  );
  al_mux2l _08667_ (
    .a(\DFF_1261.Q ),
    .b(\DFF_264.Q ),
    .s(_03312_),
    .y(\DFF_264.D )
  );
  al_ao21ftf _08668_ (
    .a(_00882_),
    .b(_02393_),
    .c(_03258_),
    .y(_03313_)
  );
  al_ao21ftf _08669_ (
    .a(g35),
    .b(\DFF_995.Q ),
    .c(_03313_),
    .y(\DFF_5.D )
  );
  al_mux2l _08670_ (
    .a(\DFF_1041.Q ),
    .b(\DFF_974.Q ),
    .s(g35),
    .y(\DFF_1041.D )
  );
  al_aoi21 _08671_ (
    .a(\DFF_344.Q ),
    .b(g35),
    .c(\DFF_1287.Q ),
    .y(_03314_)
  );
  al_oa21ftt _08672_ (
    .a(g35),
    .b(\DFF_1287.Q ),
    .c(\DFF_344.Q ),
    .y(_03315_)
  );
  al_aoi21 _08673_ (
    .a(g35),
    .b(_03315_),
    .c(_03314_),
    .y(\DFF_344.D )
  );
  al_nand3 _08674_ (
    .a(\DFF_1194.Q ),
    .b(\DFF_375.Q ),
    .c(_03125_),
    .y(_03316_)
  );
  al_oai21ttf _08675_ (
    .a(_00960_),
    .b(_01696_),
    .c(_03316_),
    .y(_03317_)
  );
  al_and3fft _08676_ (
    .a(\DFF_1110.Q ),
    .b(\DFF_422.Q ),
    .c(_00520_),
    .y(_03318_)
  );
  al_and3 _08677_ (
    .a(g35),
    .b(_03318_),
    .c(_03317_),
    .y(\DFF_422.D )
  );
  al_and2ft _08678_ (
    .a(\DFF_1287.Q ),
    .b(g35),
    .y(_03319_)
  );
  al_nand3ftt _08679_ (
    .a(\DFF_1142.Q ),
    .b(_01256_),
    .c(_03319_),
    .y(_03320_)
  );
  al_oai21ftt _08680_ (
    .a(g35),
    .b(\DFF_1287.Q ),
    .c(\DFF_1142.Q ),
    .y(_03321_)
  );
  al_nand3ftt _08681_ (
    .a(\DFF_821.Q ),
    .b(\DFF_596.Q ),
    .c(g35),
    .y(_03322_)
  );
  al_nand3 _08682_ (
    .a(_03321_),
    .b(_03322_),
    .c(_03320_),
    .y(\DFF_1287.D )
  );
  al_nand2 _08683_ (
    .a(\DFF_775.Q ),
    .b(g35),
    .y(_03323_)
  );
  al_aoi21ftt _08684_ (
    .a(\DFF_827.Q ),
    .b(_03323_),
    .c(_00959_),
    .y(\DFF_775.D )
  );
  al_nand3ftt _08685_ (
    .a(_01547_),
    .b(_01763_),
    .c(_00499_),
    .y(_03324_)
  );
  al_ao21ftt _08686_ (
    .a(_01547_),
    .b(_01763_),
    .c(\DFF_1169.Q ),
    .y(_03325_)
  );
  al_nand3 _08687_ (
    .a(g35),
    .b(_03324_),
    .c(_03325_),
    .y(_03326_)
  );
  al_ao21ftf _08688_ (
    .a(g35),
    .b(\DFF_1024.Q ),
    .c(_03326_),
    .y(\DFF_1169.D )
  );
  al_nand3 _08689_ (
    .a(_00499_),
    .b(_00705_),
    .c(_02681_),
    .y(_03327_)
  );
  al_ao21 _08690_ (
    .a(_00705_),
    .b(_02681_),
    .c(\DFF_225.Q ),
    .y(_03328_)
  );
  al_nand3 _08691_ (
    .a(g35),
    .b(_03328_),
    .c(_03327_),
    .y(_03329_)
  );
  al_ao21ftf _08692_ (
    .a(g35),
    .b(\DFF_1166.Q ),
    .c(_03329_),
    .y(\DFF_225.D )
  );
  al_nand2 _08693_ (
    .a(\DFF_395.Q ),
    .b(_01279_),
    .y(_03330_)
  );
  al_aoi21ttf _08694_ (
    .a(_03330_),
    .b(_01283_),
    .c(_01282_),
    .y(_03331_)
  );
  al_or3fft _08695_ (
    .a(\DFF_374.Q ),
    .b(_03331_),
    .c(_01858_),
    .y(_03332_)
  );
  al_oai21ftf _08696_ (
    .a(\DFF_374.Q ),
    .b(_01858_),
    .c(_03331_),
    .y(_03333_)
  );
  al_ao21 _08697_ (
    .a(_03332_),
    .b(_03333_),
    .c(_00066_),
    .y(_03334_)
  );
  al_aoi21ftf _08698_ (
    .a(\DFF_1047.Q ),
    .b(_00066_),
    .c(_03334_),
    .y(\DFF_374.D )
  );
  al_oa21ftt _08699_ (
    .a(g35),
    .b(\DFF_883.Q ),
    .c(\DFF_1217.Q ),
    .y(_03335_)
  );
  al_aoi21ftf _08700_ (
    .a(\DFF_248.Q ),
    .b(g35),
    .c(_03335_),
    .y(_03336_)
  );
  al_or3fft _08701_ (
    .a(\DFF_1078.Q ),
    .b(g35),
    .c(_03336_),
    .y(_03337_)
  );
  al_aoi21ftf _08702_ (
    .a(_00066_),
    .b(\DFF_1078.Q ),
    .c(_03336_),
    .y(_03338_)
  );
  al_nand2ft _08703_ (
    .a(_03338_),
    .b(_03337_),
    .y(\DFF_1078.D )
  );
  al_nand2 _08704_ (
    .a(g35),
    .b(_01651_),
    .y(_03339_)
  );
  al_mux2l _08705_ (
    .a(\DFF_1370.Q ),
    .b(\DFF_145.Q ),
    .s(_03339_),
    .y(\DFF_145.D )
  );
  al_nor2 _08706_ (
    .a(\DFF_1037.Q ),
    .b(g35),
    .y(_03340_)
  );
  al_nand3 _08707_ (
    .a(_00604_),
    .b(_00546_),
    .c(_00434_),
    .y(_03341_)
  );
  al_oai21ftf _08708_ (
    .a(\DFF_1375.Q ),
    .b(\DFF_1037.Q ),
    .c(\DFF_379.Q ),
    .y(_03342_)
  );
  al_nand3ftt _08709_ (
    .a(\DFF_1037.Q ),
    .b(\DFF_1375.Q ),
    .c(\DFF_379.Q ),
    .y(_03343_)
  );
  al_or3fft _08710_ (
    .a(_03342_),
    .b(_03343_),
    .c(_03341_),
    .y(_03344_)
  );
  al_aoi21 _08711_ (
    .a(\DFF_153.Q ),
    .b(_03341_),
    .c(_00066_),
    .y(_03345_)
  );
  al_aoi21 _08712_ (
    .a(_03344_),
    .b(_03345_),
    .c(_03340_),
    .y(\DFF_153.D )
  );
  al_or3fft _08713_ (
    .a(_00337_),
    .b(_01282_),
    .c(_01284_),
    .y(_03346_)
  );
  al_ao21 _08714_ (
    .a(_00337_),
    .b(_01282_),
    .c(\DFF_1135.Q ),
    .y(_03347_)
  );
  al_nand3 _08715_ (
    .a(g35),
    .b(_03347_),
    .c(_03346_),
    .y(_03348_)
  );
  al_ao21ftf _08716_ (
    .a(g35),
    .b(\DFF_1030.Q ),
    .c(_03348_),
    .y(\DFF_1135.D )
  );
  al_ao21ftt _08717_ (
    .a(g35),
    .b(\DFF_52.Q ),
    .c(_02171_),
    .y(_03349_)
  );
  al_mux2l _08718_ (
    .a(_03349_),
    .b(\DFF_1004.Q ),
    .s(_02219_),
    .y(\DFF_1004.D )
  );
  al_ao21 _08719_ (
    .a(\DFF_1217.Q ),
    .b(g35),
    .c(_01289_),
    .y(_03350_)
  );
  al_and3 _08720_ (
    .a(\DFF_1217.Q ),
    .b(g35),
    .c(_01289_),
    .y(_03351_)
  );
  al_and2ft _08721_ (
    .a(_03351_),
    .b(_03350_),
    .y(\DFF_1217.D )
  );
  al_nand3ftt _08722_ (
    .a(_00497_),
    .b(_00499_),
    .c(_01745_),
    .y(_03352_)
  );
  al_ao21ftt _08723_ (
    .a(_00497_),
    .b(_01745_),
    .c(\DFF_333.Q ),
    .y(_03353_)
  );
  al_nand3 _08724_ (
    .a(g35),
    .b(_03352_),
    .c(_03353_),
    .y(_03354_)
  );
  al_ao21ftf _08725_ (
    .a(g35),
    .b(\DFF_575.Q ),
    .c(_03354_),
    .y(\DFF_333.D )
  );
  al_ao21 _08726_ (
    .a(\DFF_490.Q ),
    .b(_01675_),
    .c(\DFF_373.Q ),
    .y(\DFF_692.D )
  );
  al_nand3 _08727_ (
    .a(_00499_),
    .b(_01763_),
    .c(_01104_),
    .y(_03355_)
  );
  al_ao21 _08728_ (
    .a(_01104_),
    .b(_01763_),
    .c(\DFF_588.Q ),
    .y(_03356_)
  );
  al_nand3 _08729_ (
    .a(g35),
    .b(_03356_),
    .c(_03355_),
    .y(_03357_)
  );
  al_ao21ftf _08730_ (
    .a(g35),
    .b(\DFF_1169.Q ),
    .c(_03357_),
    .y(\DFF_588.D )
  );
  al_and2ft _08731_ (
    .a(\DFF_709.Q ),
    .b(\DFF_1149.Q ),
    .y(_03358_)
  );
  al_or3fft _08732_ (
    .a(g35),
    .b(_03358_),
    .c(_02255_),
    .y(_03359_)
  );
  al_ao21ftf _08733_ (
    .a(g35),
    .b(\DFF_654.Q ),
    .c(_03359_),
    .y(\DFF_1059.D )
  );
  al_nor3ftt _08734_ (
    .a(\DFF_915.Q ),
    .b(_01035_),
    .c(_01034_),
    .y(_03360_)
  );
  al_nand3 _08735_ (
    .a(_01039_),
    .b(_01041_),
    .c(_03360_),
    .y(_03361_)
  );
  al_oai21ttf _08736_ (
    .a(_01035_),
    .b(_01034_),
    .c(\DFF_915.Q ),
    .y(_03362_)
  );
  al_nand3 _08737_ (
    .a(g35),
    .b(_03362_),
    .c(_03361_),
    .y(_03363_)
  );
  al_aoi21ftf _08738_ (
    .a(\DFF_1056.Q ),
    .b(_00066_),
    .c(_03363_),
    .y(\DFF_915.D )
  );
  al_mux2l _08739_ (
    .a(\DFF_753.Q ),
    .b(\DFF_1059.Q ),
    .s(g35),
    .y(\DFF_709.D )
  );
  al_ao21 _08740_ (
    .a(g35),
    .b(_01696_),
    .c(_00820_),
    .y(_03364_)
  );
  al_nand2 _08741_ (
    .a(\DFF_577.Q ),
    .b(\DFF_316.Q ),
    .y(_03365_)
  );
  al_ao21ttf _08742_ (
    .a(_03365_),
    .b(_00826_),
    .c(_00829_),
    .y(_03366_)
  );
  al_and2 _08743_ (
    .a(\DFF_1343.Q ),
    .b(g35),
    .y(_03367_)
  );
  al_ao21ttf _08744_ (
    .a(_03367_),
    .b(_03366_),
    .c(_03364_),
    .y(\DFF_1343.D )
  );
  al_and3ftt _08745_ (
    .a(\DFF_350.Q ),
    .b(g73),
    .c(g72),
    .y(_03368_)
  );
  al_nand3ftt _08746_ (
    .a(\DFF_724.Q ),
    .b(\DFF_26.Q ),
    .c(g35),
    .y(_03369_)
  );
  al_aoi21ftf _08747_ (
    .a(g35),
    .b(\DFF_663.Q ),
    .c(_03369_),
    .y(_03370_)
  );
  al_ao21ftf _08748_ (
    .a(_03368_),
    .b(_01208_),
    .c(_03370_),
    .y(\DFF_1022.D )
  );
  al_nand3 _08749_ (
    .a(_00498_),
    .b(_00499_),
    .c(_01744_),
    .y(_03371_)
  );
  al_ao21 _08750_ (
    .a(_00498_),
    .b(_01744_),
    .c(\DFF_71.Q ),
    .y(_03372_)
  );
  al_nand3 _08751_ (
    .a(g35),
    .b(_03372_),
    .c(_03371_),
    .y(_03373_)
  );
  al_ao21ftf _08752_ (
    .a(g35),
    .b(\DFF_476.Q ),
    .c(_03373_),
    .y(\DFF_71.D )
  );
  al_ao21 _08753_ (
    .a(\DFF_700.Q ),
    .b(_00935_),
    .c(_00937_),
    .y(_03374_)
  );
  al_aoi21ttf _08754_ (
    .a(\DFF_700.Q ),
    .b(_00937_),
    .c(_03374_),
    .y(_03375_)
  );
  al_mux2h _08755_ (
    .a(\DFF_83.Q ),
    .b(_03375_),
    .s(g35),
    .y(\DFF_700.D )
  );
  al_ao21ttf _08756_ (
    .a(\DFF_1168.Q ),
    .b(\DFF_801.Q ),
    .c(g35),
    .y(_03376_)
  );
  al_and2 _08757_ (
    .a(\DFF_437.Q ),
    .b(_03376_),
    .y(_03377_)
  );
  al_or3fft _08758_ (
    .a(\DFF_180.Q ),
    .b(g35),
    .c(_03377_),
    .y(_03378_)
  );
  al_aoi21ftf _08759_ (
    .a(_00066_),
    .b(\DFF_180.Q ),
    .c(_03377_),
    .y(_03379_)
  );
  al_nand2ft _08760_ (
    .a(_03379_),
    .b(_03378_),
    .y(\DFF_180.D )
  );
  al_ao21 _08761_ (
    .a(_01436_),
    .b(_01394_),
    .c(_00066_),
    .y(_03380_)
  );
  al_mux2l _08762_ (
    .a(\DFF_1034.Q ),
    .b(\DFF_1276.Q ),
    .s(_03380_),
    .y(\DFF_1276.D )
  );
  al_inv _08763_ (
    .a(\DFF_45.Q ),
    .y(_03381_)
  );
  al_aoi21 _08764_ (
    .a(\DFF_1368.Q ),
    .b(_00760_),
    .c(_00066_),
    .y(_03382_)
  );
  al_oai21 _08765_ (
    .a(\DFF_1368.Q ),
    .b(_00760_),
    .c(_03382_),
    .y(_03383_)
  );
  al_aoi21ftf _08766_ (
    .a(g35),
    .b(_03381_),
    .c(_03383_),
    .y(\DFF_1368.D )
  );
  al_ao21 _08767_ (
    .a(_00878_),
    .b(_00550_),
    .c(\DFF_763.Q ),
    .y(_03384_)
  );
  al_and2ft _08768_ (
    .a(g35),
    .b(\DFF_1033.Q ),
    .y(_03385_)
  );
  al_ao21 _08769_ (
    .a(_00552_),
    .b(_03384_),
    .c(_03385_),
    .y(\DFF_763.D )
  );
  al_oai21 _08770_ (
    .a(_01497_),
    .b(_02010_),
    .c(_02669_),
    .y(_03386_)
  );
  al_ao21ftf _08771_ (
    .a(g35),
    .b(\DFF_120.Q ),
    .c(_03386_),
    .y(\DFF_27.D )
  );
  al_and2ft _08772_ (
    .a(g35),
    .b(\DFF_977.Q ),
    .y(_03387_)
  );
  al_nand2ft _08773_ (
    .a(\DFF_1114.Q ),
    .b(\DFF_977.Q ),
    .y(_03388_)
  );
  al_nand2ft _08774_ (
    .a(\DFF_977.Q ),
    .b(\DFF_1114.Q ),
    .y(_03389_)
  );
  al_or3fft _08775_ (
    .a(_03388_),
    .b(_03389_),
    .c(_02361_),
    .y(_03390_)
  );
  al_aoi21 _08776_ (
    .a(_01486_),
    .b(_02361_),
    .c(_00066_),
    .y(_03391_)
  );
  al_ao21 _08777_ (
    .a(_03390_),
    .b(_03391_),
    .c(_03387_),
    .y(\DFF_1051.D )
  );
  al_nor2 _08778_ (
    .a(g35),
    .b(\DFF_197.Q ),
    .y(_03392_)
  );
  al_nand3 _08779_ (
    .a(_00300_),
    .b(_00301_),
    .c(_00186_),
    .y(_03393_)
  );
  al_ao21ttf _08780_ (
    .a(_00300_),
    .b(_00301_),
    .c(_00303_),
    .y(_03394_)
  );
  al_and2ft _08781_ (
    .a(g54),
    .b(_00073_),
    .y(_03395_)
  );
  al_nand3 _08782_ (
    .a(_03395_),
    .b(_03393_),
    .c(_03394_),
    .y(_03396_)
  );
  al_and2ft _08783_ (
    .a(\DFF_413.Q ),
    .b(g35),
    .y(_03397_)
  );
  al_aoi21 _08784_ (
    .a(_03397_),
    .b(_03396_),
    .c(_03392_),
    .y(\DFF_413.D )
  );
  al_mux2l _08785_ (
    .a(\DFF_599.Q ),
    .b(\DFF_539.Q ),
    .s(g35),
    .y(\DFF_503.D )
  );
  al_or3 _08786_ (
    .a(_00066_),
    .b(_00516_),
    .c(_00718_),
    .y(g28041)
  );
  al_aoi21 _08787_ (
    .a(\DFF_745.Q ),
    .b(\DFF_802.Q ),
    .c(\DFF_106.Q ),
    .y(_03398_)
  );
  al_aoi21 _08788_ (
    .a(_00936_),
    .b(_00935_),
    .c(_03398_),
    .y(_03399_)
  );
  al_nand3 _08789_ (
    .a(g35),
    .b(_00935_),
    .c(_03399_),
    .y(_03400_)
  );
  al_ao21ftf _08790_ (
    .a(g35),
    .b(\DFF_745.Q ),
    .c(_03400_),
    .y(\DFF_106.D )
  );
  al_inv _08791_ (
    .a(\DFF_37.Q ),
    .y(_03401_)
  );
  al_oai21ftf _08792_ (
    .a(g35),
    .b(_00576_),
    .c(_03401_),
    .y(_03402_)
  );
  al_nand3 _08793_ (
    .a(\DFF_1328.Q ),
    .b(g35),
    .c(_00856_),
    .y(_03403_)
  );
  al_and2ft _08794_ (
    .a(_03402_),
    .b(_03403_),
    .y(_03404_)
  );
  al_or2ft _08795_ (
    .a(_03402_),
    .b(_03403_),
    .y(_03405_)
  );
  al_nand2ft _08796_ (
    .a(_03404_),
    .b(_03405_),
    .y(\DFF_1328.D )
  );
  al_and2ft _08797_ (
    .a(g35),
    .b(\DFF_1091.Q ),
    .y(_03406_)
  );
  al_and3fft _08798_ (
    .a(\DFF_993.Q ),
    .b(\DFF_1091.Q ),
    .c(\DFF_1026.Q ),
    .y(_03407_)
  );
  al_aoi21 _08799_ (
    .a(\DFF_1231.Q ),
    .b(_00855_),
    .c(_03407_),
    .y(_03408_)
  );
  al_nand3ftt _08800_ (
    .a(\DFF_889.Q ),
    .b(\DFF_993.Q ),
    .c(\DFF_204.Q ),
    .y(_03409_)
  );
  al_nand3ftt _08801_ (
    .a(\DFF_889.Q ),
    .b(\DFF_1091.Q ),
    .c(\DFF_1030.Q ),
    .y(_03410_)
  );
  al_and3ftt _08802_ (
    .a(\DFF_1091.Q ),
    .b(\DFF_1135.Q ),
    .c(\DFF_889.Q ),
    .y(_03411_)
  );
  al_aoi21 _08803_ (
    .a(\DFF_1096.Q ),
    .b(_02820_),
    .c(_03411_),
    .y(_03412_)
  );
  al_and3 _08804_ (
    .a(_03409_),
    .b(_03410_),
    .c(_03412_),
    .y(_03413_)
  );
  al_nand3 _08805_ (
    .a(_03408_),
    .b(_00576_),
    .c(_03413_),
    .y(_03414_)
  );
  al_oa21ftf _08806_ (
    .a(_03401_),
    .b(_00576_),
    .c(_00066_),
    .y(_03415_)
  );
  al_ao21 _08807_ (
    .a(_03414_),
    .b(_03415_),
    .c(_03406_),
    .y(\DFF_37.D )
  );
  al_nand3 _08808_ (
    .a(_00499_),
    .b(_02029_),
    .c(_01497_),
    .y(_03416_)
  );
  al_ao21 _08809_ (
    .a(_01497_),
    .b(_02029_),
    .c(\DFF_1244.Q ),
    .y(_03417_)
  );
  al_nand3 _08810_ (
    .a(g35),
    .b(_03417_),
    .c(_03416_),
    .y(_03418_)
  );
  al_ao21ftf _08811_ (
    .a(g35),
    .b(\DFF_628.Q ),
    .c(_03418_),
    .y(\DFF_1244.D )
  );
  al_mux2l _08812_ (
    .a(\DFF_339.Q ),
    .b(\DFF_185.Q ),
    .s(\DFF_1122.Q ),
    .y(_03419_)
  );
  al_mux2h _08813_ (
    .a(\DFF_343.Q ),
    .b(_03419_),
    .s(g35),
    .y(\DFF_185.D )
  );
  al_aoi21 _08814_ (
    .a(\DFF_1252.Q ),
    .b(_01689_),
    .c(_00066_),
    .y(_03420_)
  );
  al_and2ft _08815_ (
    .a(g35),
    .b(\DFF_1404.Q ),
    .y(_03421_)
  );
  al_ao21 _08816_ (
    .a(_01689_),
    .b(_03091_),
    .c(\DFF_1252.Q ),
    .y(_03422_)
  );
  al_ao21 _08817_ (
    .a(_03420_),
    .b(_03422_),
    .c(_03421_),
    .y(\DFF_1252.D )
  );
  al_nand3 _08818_ (
    .a(\DFF_1057.Q ),
    .b(\DFF_1103.Q ),
    .c(_02870_),
    .y(_03423_)
  );
  al_oai21ttf _08819_ (
    .a(_01474_),
    .b(_02056_),
    .c(_03423_),
    .y(_03424_)
  );
  al_and3fft _08820_ (
    .a(\DFF_711.Q ),
    .b(\DFF_643.Q ),
    .c(_01120_),
    .y(_03425_)
  );
  al_and3 _08821_ (
    .a(g35),
    .b(_03425_),
    .c(_03424_),
    .y(\DFF_711.D )
  );
  al_nand3ftt _08822_ (
    .a(\DFF_385.Q ),
    .b(\DFF_519.Q ),
    .c(\DFF_393.Q ),
    .y(_03426_)
  );
  al_aoi21ftf _08823_ (
    .a(\DFF_1201.Q ),
    .b(_03426_),
    .c(g35),
    .y(_03427_)
  );
  al_ao21ftf _08824_ (
    .a(_03426_),
    .b(_00499_),
    .c(_03427_),
    .y(_03428_)
  );
  al_ao21ftf _08825_ (
    .a(g35),
    .b(\DFF_471.Q ),
    .c(_03428_),
    .y(\DFF_1201.D )
  );
  al_nand3ftt _08826_ (
    .a(_01547_),
    .b(_00499_),
    .c(_01787_),
    .y(_03429_)
  );
  al_ao21ftt _08827_ (
    .a(_01547_),
    .b(_01787_),
    .c(\DFF_610.Q ),
    .y(_03430_)
  );
  al_nand3 _08828_ (
    .a(g35),
    .b(_03429_),
    .c(_03430_),
    .y(_03431_)
  );
  al_ao21ftf _08829_ (
    .a(g35),
    .b(\DFF_1175.Q ),
    .c(_03431_),
    .y(\DFF_610.D )
  );
  al_and2 _08830_ (
    .a(\DFF_343.Q ),
    .b(_00717_),
    .y(_03432_)
  );
  al_ao21ftf _08831_ (
    .a(_03432_),
    .b(_00724_),
    .c(_00721_),
    .y(_03433_)
  );
  al_or3fft _08832_ (
    .a(\DFF_293.Q ),
    .b(_00722_),
    .c(_03433_),
    .y(_03434_)
  );
  al_ao21ttf _08833_ (
    .a(\DFF_293.Q ),
    .b(_00722_),
    .c(_03433_),
    .y(_03435_)
  );
  al_ao21 _08834_ (
    .a(_03434_),
    .b(_03435_),
    .c(_00066_),
    .y(_03436_)
  );
  al_aoi21ftf _08835_ (
    .a(\DFF_646.Q ),
    .b(_00066_),
    .c(_03436_),
    .y(\DFF_293.D )
  );
  al_oa21ftt _08836_ (
    .a(\DFF_701.Q ),
    .b(\DFF_548.Q ),
    .c(g35),
    .y(_03437_)
  );
  al_nand3fft _08837_ (
    .a(\DFF_701.Q ),
    .b(\DFF_1385.Q ),
    .c(g35),
    .y(_03438_)
  );
  al_aoi21ttf _08838_ (
    .a(_03438_),
    .b(_03437_),
    .c(\DFF_631.Q ),
    .y(\DFF_495.D )
  );
  al_nand3ftt _08839_ (
    .a(\DFF_1425.Q ),
    .b(\DFF_724.Q ),
    .c(_00605_),
    .y(_03439_)
  );
  al_oa21 _08840_ (
    .a(\DFF_724.Q ),
    .b(\DFF_1296.Q ),
    .c(_03439_),
    .y(_03440_)
  );
  al_oa21ttf _08841_ (
    .a(_01670_),
    .b(_01719_),
    .c(_00066_),
    .y(_03441_)
  );
  al_oai21 _08842_ (
    .a(_00605_),
    .b(_03440_),
    .c(_03441_),
    .y(_03442_)
  );
  al_ao21ftf _08843_ (
    .a(g35),
    .b(\DFF_129.Q ),
    .c(_03442_),
    .y(\DFF_1265.D )
  );
  al_or3ftt _08844_ (
    .a(\DFF_289.Q ),
    .b(\DFF_575.Q ),
    .c(\DFF_910.Q ),
    .y(_03443_)
  );
  al_aoi21ftf _08845_ (
    .a(\DFF_307.Q ),
    .b(_03443_),
    .c(g35),
    .y(_03444_)
  );
  al_ao21ftf _08846_ (
    .a(_03443_),
    .b(_00499_),
    .c(_03444_),
    .y(_03445_)
  );
  al_ao21ftf _08847_ (
    .a(g35),
    .b(\DFF_884.Q ),
    .c(_03445_),
    .y(\DFF_307.D )
  );
  al_nand3fft _08848_ (
    .a(\DFF_24.Q ),
    .b(\DFF_1136.Q ),
    .c(_00718_),
    .y(_03446_)
  );
  al_ao21ftf _08849_ (
    .a(\DFF_24.Q ),
    .b(_00718_),
    .c(\DFF_1136.Q ),
    .y(_03447_)
  );
  al_nand3 _08850_ (
    .a(_01210_),
    .b(_03446_),
    .c(_03447_),
    .y(_03448_)
  );
  al_ao21 _08851_ (
    .a(_01210_),
    .b(_01005_),
    .c(\DFF_1274.Q ),
    .y(_03449_)
  );
  al_nand3 _08852_ (
    .a(g35),
    .b(_03449_),
    .c(_03448_),
    .y(_03450_)
  );
  al_ao21ftf _08853_ (
    .a(_00088_),
    .b(_00066_),
    .c(_03450_),
    .y(\DFF_1274.D )
  );
  al_and3fft _08854_ (
    .a(\DFF_1016.Q ),
    .b(\DFF_549.Q ),
    .c(g35),
    .y(_03451_)
  );
  al_ao21ftt _08855_ (
    .a(g35),
    .b(\DFF_965.Q ),
    .c(_03451_),
    .y(\DFF_724.D )
  );
  al_and2 _08856_ (
    .a(\DFF_196.Q ),
    .b(g35),
    .y(\DFF_196.D )
  );
  al_mux2l _08857_ (
    .a(g6749),
    .b(\DFF_121.Q ),
    .s(g35),
    .y(\DFF_808.D )
  );
  al_ao21ftf _08858_ (
    .a(\DFF_1425.Q ),
    .b(g73),
    .c(_01208_),
    .y(_03452_)
  );
  al_nand3ftt _08859_ (
    .a(g72),
    .b(\DFF_724.Q ),
    .c(g35),
    .y(_03453_)
  );
  al_aoi21ftf _08860_ (
    .a(g35),
    .b(\DFF_184.Q ),
    .c(_03453_),
    .y(_03454_)
  );
  al_nand3 _08861_ (
    .a(_03369_),
    .b(_03454_),
    .c(_03452_),
    .y(\DFF_624.D )
  );
  al_ao21 _08862_ (
    .a(\DFF_359.Q ),
    .b(_00935_),
    .c(_02961_),
    .y(_03455_)
  );
  al_and2ft _08863_ (
    .a(g35),
    .b(\DFF_700.Q ),
    .y(_03456_)
  );
  al_ao21 _08864_ (
    .a(_03455_),
    .b(_02962_),
    .c(_03456_),
    .y(\DFF_359.D )
  );
  al_and2ft _08865_ (
    .a(g35),
    .b(\DFF_425.Q ),
    .y(_03457_)
  );
  al_oai21ftf _08866_ (
    .a(\DFF_793.Q ),
    .b(\DFF_1331.Q ),
    .c(\DFF_148.Q ),
    .y(_03458_)
  );
  al_nand3 _08867_ (
    .a(_00563_),
    .b(_03458_),
    .c(_00815_),
    .y(_03459_)
  );
  al_oa21ftf _08868_ (
    .a(_00559_),
    .b(_00563_),
    .c(_00066_),
    .y(_03460_)
  );
  al_ao21 _08869_ (
    .a(_03460_),
    .b(_03459_),
    .c(_03457_),
    .y(\DFF_1331.D )
  );
  al_ao21ftf _08870_ (
    .a(_01480_),
    .b(\DFF_1237.Q ),
    .c(_01479_),
    .y(_03461_)
  );
  al_and2 _08871_ (
    .a(g35),
    .b(_03461_),
    .y(_03462_)
  );
  al_aoi21 _08872_ (
    .a(\DFF_214.Q ),
    .b(\DFF_675.Q ),
    .c(\DFF_563.Q ),
    .y(_03463_)
  );
  al_ao21ftf _08873_ (
    .a(_03463_),
    .b(_01067_),
    .c(_03462_),
    .y(_03464_)
  );
  al_aoi21ftf _08874_ (
    .a(\DFF_214.Q ),
    .b(_00066_),
    .c(_03464_),
    .y(\DFF_563.D )
  );
  al_and3 _08875_ (
    .a(\DFF_525.Q ),
    .b(\DFF_710.Q ),
    .c(_01050_),
    .y(_03465_)
  );
  al_aoi21ttf _08876_ (
    .a(\DFF_524.Q ),
    .b(_03049_),
    .c(\DFF_872.Q ),
    .y(_03466_)
  );
  al_nand2ft _08877_ (
    .a(\DFF_872.Q ),
    .b(\DFF_667.Q ),
    .y(_03467_)
  );
  al_aoi21ftf _08878_ (
    .a(_03467_),
    .b(_03049_),
    .c(g35),
    .y(_03468_)
  );
  al_ao21ftf _08879_ (
    .a(_03465_),
    .b(_03466_),
    .c(_03468_),
    .y(_03469_)
  );
  al_aoi21ftf _08880_ (
    .a(\DFF_667.Q ),
    .b(_00066_),
    .c(_03469_),
    .y(\DFF_872.D )
  );
  al_nand2 _08881_ (
    .a(\DFF_214.Q ),
    .b(\DFF_675.Q ),
    .y(_03470_)
  );
  al_nor2 _08882_ (
    .a(\DFF_214.Q ),
    .b(\DFF_675.Q ),
    .y(_03471_)
  );
  al_nand2ft _08883_ (
    .a(_03471_),
    .b(_03470_),
    .y(_03472_)
  );
  al_aoi21 _08884_ (
    .a(_03472_),
    .b(_03461_),
    .c(_00066_),
    .y(\DFF_214.D )
  );
  al_and2 _08885_ (
    .a(\DFF_80.Q ),
    .b(g35),
    .y(\DFF_80.D )
  );
  al_oa21ftf _08886_ (
    .a(\DFF_835.Q ),
    .b(_01858_),
    .c(_00066_),
    .y(_03473_)
  );
  al_ao21ftf _08887_ (
    .a(\DFF_835.Q ),
    .b(_01858_),
    .c(_03473_),
    .y(_03474_)
  );
  al_aoi21ftf _08888_ (
    .a(\DFF_841.Q ),
    .b(_00066_),
    .c(_03474_),
    .y(\DFF_835.D )
  );
  al_oa21ftt _08889_ (
    .a(_00310_),
    .b(_02570_),
    .c(_02573_),
    .y(_03475_)
  );
  al_ao21ttf _08890_ (
    .a(_02569_),
    .b(_02570_),
    .c(_03475_),
    .y(_03476_)
  );
  al_ao21ftf _08891_ (
    .a(g35),
    .b(\DFF_591.Q ),
    .c(_03476_),
    .y(\DFF_353.D )
  );
  al_nand3 _08892_ (
    .a(\DFF_952.Q ),
    .b(\DFF_878.Q ),
    .c(_02338_),
    .y(_03477_)
  );
  al_nand3 _08893_ (
    .a(_00587_),
    .b(_02338_),
    .c(_00411_),
    .y(_03478_)
  );
  al_ao21 _08894_ (
    .a(\DFF_952.Q ),
    .b(_02338_),
    .c(\DFF_878.Q ),
    .y(_03479_)
  );
  al_and3 _08895_ (
    .a(_03477_),
    .b(_03479_),
    .c(_03478_),
    .y(_03480_)
  );
  al_mux2h _08896_ (
    .a(\DFF_952.Q ),
    .b(_03480_),
    .s(g35),
    .y(\DFF_878.D )
  );
  al_nor2 _08897_ (
    .a(\DFF_122.Q ),
    .b(g35),
    .y(_03481_)
  );
  al_nor3ftt _08898_ (
    .a(\DFF_49.Q ),
    .b(_00901_),
    .c(_00900_),
    .y(_03482_)
  );
  al_nand3 _08899_ (
    .a(_03482_),
    .b(_00898_),
    .c(_00894_),
    .y(_03483_)
  );
  al_oai21ttf _08900_ (
    .a(_00901_),
    .b(_00900_),
    .c(\DFF_49.Q ),
    .y(_03484_)
  );
  al_and2 _08901_ (
    .a(g35),
    .b(_03484_),
    .y(_03485_)
  );
  al_aoi21 _08902_ (
    .a(_03485_),
    .b(_03483_),
    .c(_03481_),
    .y(\DFF_49.D )
  );
  al_ao21ftf _08903_ (
    .a(_00474_),
    .b(_00488_),
    .c(_00490_),
    .y(_03486_)
  );
  al_nand3 _08904_ (
    .a(g35),
    .b(_03486_),
    .c(_01244_),
    .y(_03487_)
  );
  al_ao21ftf _08905_ (
    .a(g35),
    .b(\DFF_1339.Q ),
    .c(_03487_),
    .y(\DFF_582.D )
  );
  al_ao21ttf _08906_ (
    .a(g35),
    .b(_00516_),
    .c(\DFF_1109.Q ),
    .y(_03488_)
  );
  al_aoi21 _08907_ (
    .a(g35),
    .b(_02828_),
    .c(_03488_),
    .y(\DFF_754.D )
  );
  al_oai21 _08908_ (
    .a(\DFF_1005.Q ),
    .b(_01555_),
    .c(_02121_),
    .y(_03489_)
  );
  al_ao21ftf _08909_ (
    .a(g35),
    .b(\DFF_53.Q ),
    .c(_03489_),
    .y(\DFF_1005.D )
  );
  al_and2 _08910_ (
    .a(\DFF_598.Q ),
    .b(g35),
    .y(\DFF_678.D )
  );
  al_oa21ftt _08911_ (
    .a(g35),
    .b(\DFF_801.Q ),
    .c(\DFF_1168.Q ),
    .y(_03490_)
  );
  al_aoi21ttf _08912_ (
    .a(\DFF_1168.Q ),
    .b(g35),
    .c(\DFF_801.Q ),
    .y(_03491_)
  );
  al_oai21ftf _08913_ (
    .a(\DFF_1168.Q ),
    .b(_03490_),
    .c(_03491_),
    .y(\DFF_1168.D )
  );
  al_ao21 _08914_ (
    .a(\DFF_339.Q ),
    .b(_02196_),
    .c(\DFF_261.Q ),
    .y(_03492_)
  );
  al_and3 _08915_ (
    .a(_02198_),
    .b(_02197_),
    .c(_03492_),
    .y(\DFF_261.D )
  );
  al_nand3 _08916_ (
    .a(_00499_),
    .b(_01344_),
    .c(_02930_),
    .y(_03493_)
  );
  al_ao21 _08917_ (
    .a(_01344_),
    .b(_02930_),
    .c(\DFF_1011.Q ),
    .y(_03494_)
  );
  al_nand3 _08918_ (
    .a(g35),
    .b(_03494_),
    .c(_03493_),
    .y(_03495_)
  );
  al_ao21ftf _08919_ (
    .a(g35),
    .b(\DFF_579.Q ),
    .c(_03495_),
    .y(\DFF_1011.D )
  );
  al_nand3ftt _08920_ (
    .a(\DFF_271.Q ),
    .b(\DFF_522.Q ),
    .c(\DFF_54.Q ),
    .y(_03496_)
  );
  al_aoi21ftf _08921_ (
    .a(\DFF_645.Q ),
    .b(_03496_),
    .c(g35),
    .y(_03497_)
  );
  al_ao21ftf _08922_ (
    .a(_03496_),
    .b(_00499_),
    .c(_03497_),
    .y(_03498_)
  );
  al_ao21ftf _08923_ (
    .a(g35),
    .b(\DFF_1410.Q ),
    .c(_03498_),
    .y(\DFF_645.D )
  );
  al_ao21 _08924_ (
    .a(\DFF_68.Q ),
    .b(\DFF_1098.Q ),
    .c(\DFF_598.Q ),
    .y(_03499_)
  );
  al_nand3ftt _08925_ (
    .a(_01458_),
    .b(_03499_),
    .c(_00557_),
    .y(_03500_)
  );
  al_ao21ftf _08926_ (
    .a(g35),
    .b(\DFF_68.Q ),
    .c(_03500_),
    .y(\DFF_598.D )
  );
  al_oai21ttf _08927_ (
    .a(\DFF_188.Q ),
    .b(\DFF_474.Q ),
    .c(_01554_),
    .y(_03501_)
  );
  al_nand2ft _08928_ (
    .a(\DFF_123.Q ),
    .b(\DFF_1119.Q ),
    .y(_03502_)
  );
  al_nand2ft _08929_ (
    .a(\DFF_315.Q ),
    .b(\DFF_123.Q ),
    .y(_03503_)
  );
  al_aoi21ftf _08930_ (
    .a(\DFF_474.Q ),
    .b(\DFF_315.Q ),
    .c(_03503_),
    .y(_03504_)
  );
  al_and3 _08931_ (
    .a(g35),
    .b(_03502_),
    .c(_03504_),
    .y(_03505_)
  );
  al_and3ftt _08932_ (
    .a(_01555_),
    .b(_03501_),
    .c(_03505_),
    .y(\DFF_554.D )
  );
  al_oa21ftt _08933_ (
    .a(g35),
    .b(\DFF_801.Q ),
    .c(\DFF_578.Q ),
    .y(_03506_)
  );
  al_oa21ftf _08934_ (
    .a(\DFF_1405.Q ),
    .b(\DFF_1239.Q ),
    .c(\DFF_801.Q ),
    .y(_03507_)
  );
  al_ao21ftf _08935_ (
    .a(\DFF_578.Q ),
    .b(_03507_),
    .c(_01511_),
    .y(_03508_)
  );
  al_ao21 _08936_ (
    .a(g35),
    .b(_03508_),
    .c(_03506_),
    .y(\DFF_801.D )
  );
  al_oai21ftf _08937_ (
    .a(g35),
    .b(\DFF_736.Q ),
    .c(\DFF_669.Q ),
    .y(_03509_)
  );
  al_and3ftt _08938_ (
    .a(\DFF_736.Q ),
    .b(\DFF_669.Q ),
    .c(g35),
    .y(_03510_)
  );
  al_and2ft _08939_ (
    .a(_03510_),
    .b(_03509_),
    .y(\DFF_799.D )
  );
  al_mux2l _08940_ (
    .a(\DFF_820.Q ),
    .b(\DFF_682.Q ),
    .s(_01110_),
    .y(\DFF_682.D )
  );
  al_oa21ftt _08941_ (
    .a(g35),
    .b(\DFF_827.Q ),
    .c(\DFF_1318.Q ),
    .y(_03511_)
  );
  al_nand2ft _08942_ (
    .a(\DFF_1377.Q ),
    .b(\DFF_1249.Q ),
    .y(_03512_)
  );
  al_oa21ftf _08943_ (
    .a(\DFF_1249.Q ),
    .b(\DFF_57.Q ),
    .c(\DFF_827.Q ),
    .y(_03513_)
  );
  al_ao21ftf _08944_ (
    .a(\DFF_1318.Q ),
    .b(_03513_),
    .c(_03512_),
    .y(_03514_)
  );
  al_ao21 _08945_ (
    .a(g35),
    .b(_03514_),
    .c(_03511_),
    .y(\DFF_827.D )
  );
  al_nand3ftt _08946_ (
    .a(_00701_),
    .b(_00499_),
    .c(_02665_),
    .y(_03515_)
  );
  al_ao21ftt _08947_ (
    .a(_00701_),
    .b(_02665_),
    .c(\DFF_1291.Q ),
    .y(_03516_)
  );
  al_nand3 _08948_ (
    .a(g35),
    .b(_03515_),
    .c(_03516_),
    .y(_03517_)
  );
  al_ao21ftf _08949_ (
    .a(g35),
    .b(\DFF_526.Q ),
    .c(_03517_),
    .y(\DFF_1291.D )
  );
  al_nor2 _08950_ (
    .a(g35),
    .b(\DFF_729.Q ),
    .y(_03518_)
  );
  al_oa21ftf _08951_ (
    .a(\DFF_697.Q ),
    .b(_02064_),
    .c(_00066_),
    .y(_03519_)
  );
  al_aoi21 _08952_ (
    .a(_03519_),
    .b(_02105_),
    .c(_03518_),
    .y(\DFF_697.D )
  );
  al_nand3 _08953_ (
    .a(_00499_),
    .b(_00596_),
    .c(_02426_),
    .y(_03520_)
  );
  al_ao21 _08954_ (
    .a(_02426_),
    .b(_00596_),
    .c(\DFF_550.Q ),
    .y(_03521_)
  );
  al_nand3 _08955_ (
    .a(g35),
    .b(_03521_),
    .c(_03520_),
    .y(_03522_)
  );
  al_ao21ftf _08956_ (
    .a(g35),
    .b(\DFF_1160.Q ),
    .c(_03522_),
    .y(\DFF_550.D )
  );
  al_and2ft _08957_ (
    .a(g35),
    .b(\DFF_1379.Q ),
    .y(_03523_)
  );
  al_oa21 _08958_ (
    .a(\DFF_1084.Q ),
    .b(_00609_),
    .c(_00607_),
    .y(_03524_)
  );
  al_ao21 _08959_ (
    .a(_01936_),
    .b(_03524_),
    .c(_03523_),
    .y(\DFF_1084.D )
  );
  al_nor3fft _08960_ (
    .a(_03073_),
    .b(_03072_),
    .c(_03070_),
    .y(_03525_)
  );
  al_and2ft _08961_ (
    .a(_03068_),
    .b(_03072_),
    .y(_03526_)
  );
  al_and3ftt _08962_ (
    .a(\DFF_1203.Q ),
    .b(\DFF_987.Q ),
    .c(g35),
    .y(_03527_)
  );
  al_nand3ftt _08963_ (
    .a(_03069_),
    .b(_03527_),
    .c(_03526_),
    .y(_03528_)
  );
  al_or2 _08964_ (
    .a(\DFF_688.Q ),
    .b(\DFF_1409.Q ),
    .y(_03529_)
  );
  al_ao21 _08965_ (
    .a(\DFF_688.Q ),
    .b(\DFF_1409.Q ),
    .c(\DFF_742.Q ),
    .y(_03530_)
  );
  al_nand3 _08966_ (
    .a(g35),
    .b(_03529_),
    .c(_03530_),
    .y(_03531_)
  );
  al_nand3 _08967_ (
    .a(_03070_),
    .b(_03531_),
    .c(_03074_),
    .y(_03532_)
  );
  al_and3 _08968_ (
    .a(g35),
    .b(_03069_),
    .c(_03068_),
    .y(_03533_)
  );
  al_ao21 _08969_ (
    .a(_03532_),
    .b(_03528_),
    .c(_03533_),
    .y(_03534_)
  );
  al_and2 _08970_ (
    .a(\DFF_1203.Q ),
    .b(g35),
    .y(_03535_)
  );
  al_ao21 _08971_ (
    .a(\DFF_1021.Q ),
    .b(\DFF_1121.Q ),
    .c(\DFF_679.Q ),
    .y(_03536_)
  );
  al_and3 _08972_ (
    .a(g35),
    .b(_03071_),
    .c(_03536_),
    .y(_03537_)
  );
  al_or3 _08973_ (
    .a(_03068_),
    .b(_03537_),
    .c(_03072_),
    .y(_03538_)
  );
  al_oa21ttf _08974_ (
    .a(\DFF_987.Q ),
    .b(_03069_),
    .c(_00066_),
    .y(_03539_)
  );
  al_oa21ftf _08975_ (
    .a(_03535_),
    .b(_03526_),
    .c(_03539_),
    .y(_03540_)
  );
  al_ao21ftf _08976_ (
    .a(_03535_),
    .b(_03538_),
    .c(_03540_),
    .y(_03541_)
  );
  al_nand3ftt _08977_ (
    .a(_03525_),
    .b(_03541_),
    .c(_03534_),
    .y(g31793)
  );
  al_ao21 _08978_ (
    .a(\DFF_853.Q ),
    .b(_00601_),
    .c(\DFF_1173.Q ),
    .y(_03542_)
  );
  al_nand3ftt _08979_ (
    .a(_01426_),
    .b(_03542_),
    .c(_01505_),
    .y(_03543_)
  );
  al_ao21ftf _08980_ (
    .a(g35),
    .b(\DFF_853.Q ),
    .c(_03543_),
    .y(\DFF_1173.D )
  );
  al_nand3 _08981_ (
    .a(_00499_),
    .b(_01772_),
    .c(_01702_),
    .y(_03544_)
  );
  al_ao21 _08982_ (
    .a(_01772_),
    .b(_01702_),
    .c(\DFF_55.Q ),
    .y(_03545_)
  );
  al_nand3 _08983_ (
    .a(g35),
    .b(_03544_),
    .c(_03545_),
    .y(_03546_)
  );
  al_ao21ftf _08984_ (
    .a(g35),
    .b(\DFF_1297.Q ),
    .c(_03546_),
    .y(\DFF_55.D )
  );
  al_and3fft _08985_ (
    .a(\DFF_212.Q ),
    .b(\DFF_446.Q ),
    .c(g35),
    .y(_03547_)
  );
  al_oai21ftt _08986_ (
    .a(g35),
    .b(\DFF_446.Q ),
    .c(\DFF_212.Q ),
    .y(_03548_)
  );
  al_nand2ft _08987_ (
    .a(_03547_),
    .b(_03548_),
    .y(_03549_)
  );
  al_mux2l _08988_ (
    .a(_03549_),
    .b(\DFF_1277.Q ),
    .s(_01569_),
    .y(\DFF_1277.D )
  );
  al_nand3ftt _08989_ (
    .a(_02157_),
    .b(g35),
    .c(_02152_),
    .y(g26877)
  );
  al_mux2l _08990_ (
    .a(\DFF_446.Q ),
    .b(\DFF_212.Q ),
    .s(_01569_),
    .y(\DFF_212.D )
  );
  al_and2ft _08991_ (
    .a(g35),
    .b(\DFF_568.Q ),
    .y(_03550_)
  );
  al_inv _08992_ (
    .a(\DFF_189.Q ),
    .y(_03551_)
  );
  al_nand3fft _08993_ (
    .a(\DFF_623.Q ),
    .b(_03551_),
    .c(_00758_),
    .y(_03552_)
  );
  al_nand2ft _08994_ (
    .a(\DFF_682.Q ),
    .b(\DFF_568.Q ),
    .y(_03553_)
  );
  al_nand2ft _08995_ (
    .a(\DFF_568.Q ),
    .b(\DFF_682.Q ),
    .y(_03554_)
  );
  al_or3fft _08996_ (
    .a(_03553_),
    .b(_03554_),
    .c(_03552_),
    .y(_03555_)
  );
  al_aoi21 _08997_ (
    .a(_03381_),
    .b(_03552_),
    .c(_00066_),
    .y(_03556_)
  );
  al_ao21 _08998_ (
    .a(_03555_),
    .b(_03556_),
    .c(_03550_),
    .y(\DFF_45.D )
  );
  al_nand3 _08999_ (
    .a(\DFF_1251.Q ),
    .b(_02824_),
    .c(_03465_),
    .y(_03557_)
  );
  al_ao21 _09000_ (
    .a(_02824_),
    .b(_03465_),
    .c(\DFF_1251.Q ),
    .y(_03558_)
  );
  al_nand3 _09001_ (
    .a(_02027_),
    .b(_03557_),
    .c(_03558_),
    .y(_03559_)
  );
  al_ao21ftf _09002_ (
    .a(g35),
    .b(\DFF_710.Q ),
    .c(_03559_),
    .y(\DFF_1251.D )
  );
  al_and2 _09003_ (
    .a(\DFF_575.Q ),
    .b(g35),
    .y(\DFF_630.D )
  );
  al_or2ft _09004_ (
    .a(\DFF_1284.Q ),
    .b(g26801),
    .y(_03560_)
  );
  al_inv _09005_ (
    .a(\DFF_1398.Q ),
    .y(_03561_)
  );
  al_and2ft _09006_ (
    .a(\DFF_1211.Q ),
    .b(g35),
    .y(_03562_)
  );
  al_ao21ftf _09007_ (
    .a(_03561_),
    .b(_03562_),
    .c(_01458_),
    .y(_03563_)
  );
  al_and3ftt _09008_ (
    .a(_03562_),
    .b(_03561_),
    .c(_01458_),
    .y(_03564_)
  );
  al_aoi21 _09009_ (
    .a(_03560_),
    .b(_03563_),
    .c(_03564_),
    .y(\DFF_1284.D )
  );
  al_ao21 _09010_ (
    .a(_00948_),
    .b(_00947_),
    .c(\DFF_876.Q ),
    .y(_03565_)
  );
  al_nand3fft _09011_ (
    .a(_01837_),
    .b(_01178_),
    .c(_03565_),
    .y(_03566_)
  );
  al_ao21ftf _09012_ (
    .a(g35),
    .b(\DFF_256.Q ),
    .c(_03566_),
    .y(\DFF_876.D )
  );
  al_mux2l _09013_ (
    .a(\DFF_1187.Q ),
    .b(\DFF_1230.Q ),
    .s(_02950_),
    .y(_03567_)
  );
  al_mux2h _09014_ (
    .a(\DFF_689.Q ),
    .b(_03567_),
    .s(g35),
    .y(\DFF_1187.D )
  );
  al_nor2 _09015_ (
    .a(\DFF_1236.Q ),
    .b(g35),
    .y(_03568_)
  );
  al_and3 _09016_ (
    .a(_00604_),
    .b(_01363_),
    .c(_00438_),
    .y(_03569_)
  );
  al_nand3ftt _09017_ (
    .a(\DFF_1236.Q ),
    .b(\DFF_1295.Q ),
    .c(\DFF_379.Q ),
    .y(_03570_)
  );
  al_oai21ftf _09018_ (
    .a(\DFF_1295.Q ),
    .b(\DFF_1236.Q ),
    .c(\DFF_379.Q ),
    .y(_03571_)
  );
  al_nand3 _09019_ (
    .a(_03570_),
    .b(_03571_),
    .c(_03569_),
    .y(_03572_)
  );
  al_oa21ftf _09020_ (
    .a(\DFF_1093.Q ),
    .b(_03569_),
    .c(_00066_),
    .y(_03573_)
  );
  al_aoi21 _09021_ (
    .a(_03572_),
    .b(_03573_),
    .c(_03568_),
    .y(\DFF_1093.D )
  );
  al_oai21 _09022_ (
    .a(_00592_),
    .b(_02871_),
    .c(_02365_),
    .y(_03574_)
  );
  al_ao21ftf _09023_ (
    .a(g35),
    .b(\DFF_734.Q ),
    .c(_03574_),
    .y(\DFF_723.D )
  );
  al_nor2 _09024_ (
    .a(g35),
    .b(\DFF_1403.Q ),
    .y(_03575_)
  );
  al_and3fft _09025_ (
    .a(\DFF_531.Q ),
    .b(\DFF_708.Q ),
    .c(g35),
    .y(_03576_)
  );
  al_aoi21 _09026_ (
    .a(_03576_),
    .b(_00515_),
    .c(_03575_),
    .y(\DFF_531.D )
  );
  al_oai21 _09027_ (
    .a(\DFF_919.Q ),
    .b(\DFF_1417.Q ),
    .c(g35),
    .y(_03577_)
  );
  al_ao21ftf _09028_ (
    .a(g35),
    .b(\DFF_325.Q ),
    .c(_03577_),
    .y(\DFF_1417.D )
  );
  al_nand3 _09029_ (
    .a(_01826_),
    .b(\DFF_719.Q ),
    .c(_01579_),
    .y(_03578_)
  );
  al_aoi21ftf _09030_ (
    .a(_01174_),
    .b(\DFF_1053.Q ),
    .c(_03578_),
    .y(_03579_)
  );
  al_ao21ftf _09031_ (
    .a(g35),
    .b(\DFF_542.Q ),
    .c(_03579_),
    .y(\DFF_1053.D )
  );
  al_nand3 _09032_ (
    .a(_00332_),
    .b(_00641_),
    .c(_01618_),
    .y(_03580_)
  );
  al_ao21 _09033_ (
    .a(_00332_),
    .b(_00641_),
    .c(\DFF_1380.Q ),
    .y(_03581_)
  );
  al_nand3 _09034_ (
    .a(g35),
    .b(_03581_),
    .c(_03580_),
    .y(_03582_)
  );
  al_ao21ftf _09035_ (
    .a(g35),
    .b(\DFF_1097.Q ),
    .c(_03582_),
    .y(\DFF_1380.D )
  );
  al_and3 _09036_ (
    .a(\DFF_1382.Q ),
    .b(_02242_),
    .c(_01211_),
    .y(_03583_)
  );
  al_or2 _09037_ (
    .a(_00255_),
    .b(_03583_),
    .y(_03584_)
  );
  al_nand2 _09038_ (
    .a(_00255_),
    .b(_03583_),
    .y(_03585_)
  );
  al_nand3 _09039_ (
    .a(g35),
    .b(_03585_),
    .c(_03584_),
    .y(_03586_)
  );
  al_aoi21ftf _09040_ (
    .a(\DFF_1382.Q ),
    .b(_00066_),
    .c(_03586_),
    .y(\DFF_137.D )
  );
  al_and2ft _09041_ (
    .a(g35),
    .b(\DFF_683.Q ),
    .y(_03587_)
  );
  al_ao21 _09042_ (
    .a(_02338_),
    .b(_03478_),
    .c(\DFF_952.Q ),
    .y(_03588_)
  );
  al_aoi21 _09043_ (
    .a(\DFF_952.Q ),
    .b(_02338_),
    .c(_00066_),
    .y(_03589_)
  );
  al_ao21 _09044_ (
    .a(_03589_),
    .b(_03588_),
    .c(_03587_),
    .y(\DFF_952.D )
  );
  al_nand3 _09045_ (
    .a(_00641_),
    .b(_01844_),
    .c(_01618_),
    .y(_03590_)
  );
  al_ao21 _09046_ (
    .a(_01844_),
    .b(_00641_),
    .c(\DFF_890.Q ),
    .y(_03591_)
  );
  al_nand3 _09047_ (
    .a(g35),
    .b(_03591_),
    .c(_03590_),
    .y(_03592_)
  );
  al_ao21ftf _09048_ (
    .a(g35),
    .b(\DFF_1380.Q ),
    .c(_03592_),
    .y(\DFF_890.D )
  );
  al_nand3ftt _09049_ (
    .a(_01768_),
    .b(_02624_),
    .c(_00499_),
    .y(_03593_)
  );
  al_ao21ftt _09050_ (
    .a(_01768_),
    .b(_02624_),
    .c(\DFF_158.Q ),
    .y(_03594_)
  );
  al_nand3 _09051_ (
    .a(g35),
    .b(_03593_),
    .c(_03594_),
    .y(_03595_)
  );
  al_ao21ftf _09052_ (
    .a(g35),
    .b(\DFF_92.Q ),
    .c(_03595_),
    .y(\DFF_158.D )
  );
  al_oa21ftt _09053_ (
    .a(g35),
    .b(\DFF_1287.Q ),
    .c(\DFF_978.Q ),
    .y(_03596_)
  );
  al_aoi21ftf _09054_ (
    .a(\DFF_344.Q ),
    .b(g35),
    .c(_03596_),
    .y(_03597_)
  );
  al_or3fft _09055_ (
    .a(\DFF_138.Q ),
    .b(g35),
    .c(_03597_),
    .y(_03598_)
  );
  al_aoi21ftf _09056_ (
    .a(_00066_),
    .b(\DFF_138.Q ),
    .c(_03597_),
    .y(_03599_)
  );
  al_nand2ft _09057_ (
    .a(_03599_),
    .b(_03598_),
    .y(\DFF_138.D )
  );
  al_nand3 _09058_ (
    .a(_00499_),
    .b(_00705_),
    .c(_02754_),
    .y(_03600_)
  );
  al_ao21 _09059_ (
    .a(_00705_),
    .b(_02754_),
    .c(\DFF_370.Q ),
    .y(_03601_)
  );
  al_nand3 _09060_ (
    .a(g35),
    .b(_03601_),
    .c(_03600_),
    .y(_03602_)
  );
  al_ao21ftf _09061_ (
    .a(g35),
    .b(\DFF_1218.Q ),
    .c(_03602_),
    .y(\DFF_370.D )
  );
  al_nand2ft _09062_ (
    .a(g126),
    .b(g120),
    .y(_03603_)
  );
  al_and3ftt _09063_ (
    .a(\DFF_673.Q ),
    .b(g35),
    .c(_03603_),
    .y(_03604_)
  );
  al_aoi21ftf _09064_ (
    .a(g120),
    .b(g126),
    .c(_03604_),
    .y(_03605_)
  );
  al_nand2ft _09065_ (
    .a(g35),
    .b(\DFF_1083.Q ),
    .y(_03606_)
  );
  al_and2ft _09066_ (
    .a(\DFF_767.Q ),
    .b(g35),
    .y(_03607_)
  );
  al_aoi21ftf _09067_ (
    .a(g115),
    .b(g114),
    .c(_03607_),
    .y(_03608_)
  );
  al_ao21ftf _09068_ (
    .a(g114),
    .b(g115),
    .c(_03608_),
    .y(_03609_)
  );
  al_or3fft _09069_ (
    .a(_03606_),
    .b(_03609_),
    .c(_03605_),
    .y(\DFF_116.D )
  );
  al_ao21 _09070_ (
    .a(\DFF_43.Q ),
    .b(\DFF_331.Q ),
    .c(\DFF_1412.Q ),
    .y(_03610_)
  );
  al_and3ftt _09071_ (
    .a(_01526_),
    .b(_03610_),
    .c(_01848_),
    .y(_03611_)
  );
  al_mux2h _09072_ (
    .a(\DFF_43.Q ),
    .b(_03611_),
    .s(g35),
    .y(\DFF_1412.D )
  );
  al_nand3 _09073_ (
    .a(\DFF_424.Q ),
    .b(_01261_),
    .c(_02796_),
    .y(_03612_)
  );
  al_inv _09074_ (
    .a(\DFF_595.Q ),
    .y(_03613_)
  );
  al_aoi21 _09075_ (
    .a(_03613_),
    .b(_03612_),
    .c(_00066_),
    .y(_03614_)
  );
  al_ao21ftf _09076_ (
    .a(_03612_),
    .b(\DFF_595.Q ),
    .c(_03614_),
    .y(_03615_)
  );
  al_ao21ftf _09077_ (
    .a(g35),
    .b(\DFF_424.Q ),
    .c(_03615_),
    .y(\DFF_595.D )
  );
  al_or2ft _09078_ (
    .a(\DFF_1198.Q ),
    .b(_00358_),
    .y(_03616_)
  );
  al_inv _09079_ (
    .a(\DFF_1332.Q ),
    .y(_03617_)
  );
  al_ao21ftf _09080_ (
    .a(_03617_),
    .b(_01961_),
    .c(_01393_),
    .y(_03618_)
  );
  al_and3ftt _09081_ (
    .a(_01961_),
    .b(_03617_),
    .c(_01393_),
    .y(_03619_)
  );
  al_aoi21 _09082_ (
    .a(_03616_),
    .b(_03618_),
    .c(_03619_),
    .y(\DFF_1198.D )
  );
  al_nand3 _09083_ (
    .a(\DFF_1141.Q ),
    .b(_01414_),
    .c(_01282_),
    .y(_03620_)
  );
  al_aoi21ftf _09084_ (
    .a(\DFF_1030.Q ),
    .b(_03620_),
    .c(g35),
    .y(_03621_)
  );
  al_oai21 _09085_ (
    .a(_01284_),
    .b(_03620_),
    .c(_03621_),
    .y(_03622_)
  );
  al_ao21ftf _09086_ (
    .a(g35),
    .b(\DFF_1231.Q ),
    .c(_03622_),
    .y(\DFF_1030.D )
  );
  al_nand3fft _09087_ (
    .a(\DFF_1010.Q ),
    .b(_00514_),
    .c(_00526_),
    .y(_03623_)
  );
  al_aoi21ftf _09088_ (
    .a(\DFF_65.Q ),
    .b(_03623_),
    .c(g35),
    .y(_03624_)
  );
  al_ao21ftf _09089_ (
    .a(_03623_),
    .b(_00530_),
    .c(_03624_),
    .y(_03625_)
  );
  al_ao21ftf _09090_ (
    .a(g35),
    .b(\DFF_4.Q ),
    .c(_03625_),
    .y(\DFF_65.D )
  );
  al_aoi21ttf _09091_ (
    .a(\DFF_1124.Q ),
    .b(g35),
    .c(\DFF_288.Q ),
    .y(_03626_)
  );
  al_mux2l _09092_ (
    .a(_01418_),
    .b(_03626_),
    .s(_01419_),
    .y(\DFF_722.D )
  );
  al_oa21ttf _09093_ (
    .a(\DFF_1298.Q ),
    .b(\DFF_805.Q ),
    .c(\DFF_36.Q ),
    .y(_03627_)
  );
  al_and3fft _09094_ (
    .a(\DFF_1298.Q ),
    .b(\DFF_805.Q ),
    .c(\DFF_36.Q ),
    .y(_03628_)
  );
  al_nor2ft _09095_ (
    .a(g35),
    .b(_03628_),
    .y(_03629_)
  );
  al_ao21ttf _09096_ (
    .a(_03627_),
    .b(_01455_),
    .c(_03629_),
    .y(_03630_)
  );
  al_aoi21ftf _09097_ (
    .a(\DFF_805.Q ),
    .b(_00066_),
    .c(_03630_),
    .y(\DFF_36.D )
  );
  al_oa21ftf _09098_ (
    .a(\DFF_1016.Q ),
    .b(\DFF_965.Q ),
    .c(\DFF_440.Q ),
    .y(_03631_)
  );
  al_nand2 _09099_ (
    .a(_03631_),
    .b(_01824_),
    .y(_03632_)
  );
  al_mux2h _09100_ (
    .a(\DFF_436.Q ),
    .b(_03632_),
    .s(g35),
    .y(\DFF_1016.D )
  );
  al_mux2l _09101_ (
    .a(\DFF_706.Q ),
    .b(\DFF_1125.Q ),
    .s(g35),
    .y(\DFF_706.D )
  );
  al_or3fft _09102_ (
    .a(g35),
    .b(_01078_),
    .c(_01082_),
    .y(g26876)
  );
  al_ao21 _09103_ (
    .a(\DFF_524.Q ),
    .b(_03049_),
    .c(_01606_),
    .y(_03633_)
  );
  al_nand3ftt _09104_ (
    .a(\DFF_23.Q ),
    .b(\DFF_1251.Q ),
    .c(_02824_),
    .y(_03634_)
  );
  al_ao21ttf _09105_ (
    .a(_03467_),
    .b(_03634_),
    .c(_01579_),
    .y(_03635_)
  );
  al_nand2ft _09106_ (
    .a(g35),
    .b(\DFF_23.Q ),
    .y(_03636_)
  );
  al_nand3 _09107_ (
    .a(_03636_),
    .b(_03635_),
    .c(_03633_),
    .y(\DFF_667.D )
  );
  al_mux2l _09108_ (
    .a(\DFF_510.Q ),
    .b(\DFF_544.Q ),
    .s(_01174_),
    .y(\DFF_544.D )
  );
  al_mux2l _09109_ (
    .a(\DFF_1211.Q ),
    .b(\DFF_1398.Q ),
    .s(_01458_),
    .y(\DFF_1398.D )
  );
  al_or2ft _09110_ (
    .a(\DFF_1161.Q ),
    .b(_01582_),
    .y(_03637_)
  );
  al_nand2ft _09111_ (
    .a(\DFF_1161.Q ),
    .b(_01582_),
    .y(_03638_)
  );
  al_nand3 _09112_ (
    .a(g35),
    .b(_03638_),
    .c(_03637_),
    .y(_03639_)
  );
  al_aoi21ftf _09113_ (
    .a(\DFF_798.Q ),
    .b(_00066_),
    .c(_03639_),
    .y(\DFF_1161.D )
  );
  al_nand3fft _09114_ (
    .a(_01755_),
    .b(_02597_),
    .c(_01150_),
    .y(_03640_)
  );
  al_aoi21ftf _09115_ (
    .a(\DFF_465.Q ),
    .b(_03640_),
    .c(g35),
    .y(_03641_)
  );
  al_oai21 _09116_ (
    .a(_01153_),
    .b(_03640_),
    .c(_03641_),
    .y(_03642_)
  );
  al_ao21ftf _09117_ (
    .a(g35),
    .b(\DFF_641.Q ),
    .c(_03642_),
    .y(\DFF_465.D )
  );
  al_nor2 _09118_ (
    .a(\DFF_308.Q ),
    .b(g35),
    .y(_03643_)
  );
  al_mux2l _09119_ (
    .a(_02000_),
    .b(_01996_),
    .s(_01993_),
    .y(_03644_)
  );
  al_or3fft _09120_ (
    .a(\DFF_1271.Q ),
    .b(_02164_),
    .c(_03644_),
    .y(_03645_)
  );
  al_aoi21ftf _09121_ (
    .a(\DFF_1271.Q ),
    .b(_03644_),
    .c(g35),
    .y(_03646_)
  );
  al_aoi21 _09122_ (
    .a(_03645_),
    .b(_03646_),
    .c(_03643_),
    .y(\DFF_1271.D )
  );
  al_and2ft _09123_ (
    .a(g35),
    .b(\DFF_39.Q ),
    .y(_03647_)
  );
  al_ao21 _09124_ (
    .a(_00766_),
    .b(_01219_),
    .c(\DFF_1312.Q ),
    .y(_03648_)
  );
  al_aoi21 _09125_ (
    .a(\DFF_1312.Q ),
    .b(_00766_),
    .c(_00066_),
    .y(_03649_)
  );
  al_ao21 _09126_ (
    .a(_03649_),
    .b(_03648_),
    .c(_03647_),
    .y(\DFF_1312.D )
  );
  al_nor2 _09127_ (
    .a(\DFF_1321.Q ),
    .b(g35),
    .y(_03650_)
  );
  al_nand3ftt _09128_ (
    .a(_01298_),
    .b(\DFF_97.Q ),
    .c(_00899_),
    .y(_03651_)
  );
  al_aoi21ftf _09129_ (
    .a(\DFF_97.Q ),
    .b(_01298_),
    .c(g35),
    .y(_03652_)
  );
  al_aoi21 _09130_ (
    .a(_03652_),
    .b(_03651_),
    .c(_03650_),
    .y(\DFF_97.D )
  );
  al_and2 _09131_ (
    .a(\DFF_1275.Q ),
    .b(\DFF_913.Q ),
    .y(_03653_)
  );
  al_ao21 _09132_ (
    .a(\DFF_454.Q ),
    .b(_01317_),
    .c(_03653_),
    .y(_03654_)
  );
  al_nand3 _09133_ (
    .a(g35),
    .b(_02828_),
    .c(_03654_),
    .y(_03655_)
  );
  al_ao21ftf _09134_ (
    .a(g35),
    .b(\DFF_454.Q ),
    .c(_03655_),
    .y(\DFF_913.D )
  );
  al_nand3 _09135_ (
    .a(\DFF_671.Q ),
    .b(_02597_),
    .c(_01150_),
    .y(_03656_)
  );
  al_aoi21ftf _09136_ (
    .a(\DFF_924.Q ),
    .b(_03656_),
    .c(g35),
    .y(_03657_)
  );
  al_oai21 _09137_ (
    .a(_01153_),
    .b(_03656_),
    .c(_03657_),
    .y(_03658_)
  );
  al_ao21ftf _09138_ (
    .a(g35),
    .b(\DFF_1394.Q ),
    .c(_03658_),
    .y(\DFF_924.D )
  );
  al_aoi21ftt _09139_ (
    .a(\DFF_486.Q ),
    .b(\DFF_979.Q ),
    .c(_02056_),
    .y(_03659_)
  );
  al_nand3fft _09140_ (
    .a(_00066_),
    .b(\DFF_486.Q ),
    .c(_02056_),
    .y(_03660_)
  );
  al_aoi21ftf _09141_ (
    .a(\DFF_131.Q ),
    .b(_00066_),
    .c(_03660_),
    .y(_03661_)
  );
  al_aoi21ftf _09142_ (
    .a(_00066_),
    .b(_03659_),
    .c(_03661_),
    .y(\DFF_486.D )
  );
  al_and3 _09143_ (
    .a(\DFF_563.Q ),
    .b(\DFF_214.Q ),
    .c(\DFF_600.Q ),
    .y(_03662_)
  );
  al_nand3 _09144_ (
    .a(\DFF_921.Q ),
    .b(_01211_),
    .c(_03662_),
    .y(_03663_)
  );
  al_nand2 _09145_ (
    .a(\DFF_1046.Q ),
    .b(_03663_),
    .y(_03664_)
  );
  al_or2 _09146_ (
    .a(\DFF_1046.Q ),
    .b(_03663_),
    .y(_03665_)
  );
  al_nand3 _09147_ (
    .a(g35),
    .b(_03664_),
    .c(_03665_),
    .y(_03666_)
  );
  al_aoi21ftf _09148_ (
    .a(\DFF_921.Q ),
    .b(_00066_),
    .c(_03666_),
    .y(\DFF_1046.D )
  );
  al_nand3 _09149_ (
    .a(_00499_),
    .b(_00592_),
    .c(_02665_),
    .y(_03667_)
  );
  al_ao21 _09150_ (
    .a(_00592_),
    .b(_02665_),
    .c(\DFF_815.Q ),
    .y(_03668_)
  );
  al_nand3 _09151_ (
    .a(g35),
    .b(_03668_),
    .c(_03667_),
    .y(_03669_)
  );
  al_ao21ftf _09152_ (
    .a(g35),
    .b(\DFF_1058.Q ),
    .c(_03669_),
    .y(\DFF_815.D )
  );
  al_inv _09153_ (
    .a(\DFF_511.Q ),
    .y(_03670_)
  );
  al_and2ft _09154_ (
    .a(\DFF_698.Q ),
    .b(\DFF_791.Q ),
    .y(_03671_)
  );
  al_nand2ft _09155_ (
    .a(\DFF_791.Q ),
    .b(\DFF_698.Q ),
    .y(_03672_)
  );
  al_nand2ft _09156_ (
    .a(_03671_),
    .b(_03672_),
    .y(_03673_)
  );
  al_and3fft _09157_ (
    .a(_01474_),
    .b(_02056_),
    .c(_03673_),
    .y(_03674_)
  );
  al_ao21 _09158_ (
    .a(g35),
    .b(_03674_),
    .c(_03670_),
    .y(_03675_)
  );
  al_and3 _09159_ (
    .a(_03670_),
    .b(g35),
    .c(_03674_),
    .y(_03676_)
  );
  al_nand2ft _09160_ (
    .a(_03676_),
    .b(_03675_),
    .y(\DFF_1207.D )
  );
  al_mux2h _09161_ (
    .a(\DFF_1124.Q ),
    .b(_01096_),
    .s(g35),
    .y(\DFF_1116.D )
  );
  al_oai21ftt _09162_ (
    .a(g35),
    .b(_02775_),
    .c(\DFF_772.Q ),
    .y(_03677_)
  );
  al_nand3 _09163_ (
    .a(\DFF_777.Q ),
    .b(g35),
    .c(_02923_),
    .y(_03678_)
  );
  al_and2ft _09164_ (
    .a(_03677_),
    .b(_03678_),
    .y(_03679_)
  );
  al_or2ft _09165_ (
    .a(_03677_),
    .b(_03678_),
    .y(_03680_)
  );
  al_nand2ft _09166_ (
    .a(_03679_),
    .b(_03680_),
    .y(\DFF_777.D )
  );
  al_and2ft _09167_ (
    .a(\DFF_170.Q ),
    .b(\DFF_300.Q ),
    .y(_03681_)
  );
  al_nand2ft _09168_ (
    .a(\DFF_300.Q ),
    .b(\DFF_170.Q ),
    .y(_03682_)
  );
  al_nand2ft _09169_ (
    .a(_03681_),
    .b(_03682_),
    .y(_03683_)
  );
  al_mux2l _09170_ (
    .a(\DFF_1203.Q ),
    .b(_03683_),
    .s(_01665_),
    .y(_03684_)
  );
  al_mux2h _09171_ (
    .a(\DFF_170.Q ),
    .b(_03684_),
    .s(g35),
    .y(\DFF_1203.D )
  );
  al_oai21 _09172_ (
    .a(_01266_),
    .b(_02707_),
    .c(_02726_),
    .y(_03685_)
  );
  al_ao21ftf _09173_ (
    .a(g35),
    .b(\DFF_784.Q ),
    .c(_03685_),
    .y(\DFF_776.D )
  );
  al_ao21 _09174_ (
    .a(_01832_),
    .b(_01815_),
    .c(\DFF_551.Q ),
    .y(_03686_)
  );
  al_nand3fft _09175_ (
    .a(_01831_),
    .b(_02659_),
    .c(_03686_),
    .y(_03687_)
  );
  al_ao21ftf _09176_ (
    .a(g35),
    .b(\DFF_411.Q ),
    .c(_03687_),
    .y(\DFF_551.D )
  );
  al_and2ft _09177_ (
    .a(g35),
    .b(\DFF_660.Q ),
    .y(_03688_)
  );
  al_oai21ftf _09178_ (
    .a(\DFF_660.Q ),
    .b(_02227_),
    .c(\DFF_807.Q ),
    .y(_03689_)
  );
  al_ao21 _09179_ (
    .a(_02228_),
    .b(_03689_),
    .c(_03688_),
    .y(\DFF_807.D )
  );
  al_nand3 _09180_ (
    .a(\DFF_170.Q ),
    .b(_01665_),
    .c(_03005_),
    .y(_03690_)
  );
  al_ao21 _09181_ (
    .a(\DFF_170.Q ),
    .b(_01665_),
    .c(_03005_),
    .y(_03691_)
  );
  al_nand3 _09182_ (
    .a(g35),
    .b(_03690_),
    .c(_03691_),
    .y(_03692_)
  );
  al_aoi21ftf _09183_ (
    .a(\DFF_300.Q ),
    .b(_00066_),
    .c(_03692_),
    .y(\DFF_170.D )
  );
  al_or2ft _09184_ (
    .a(g35),
    .b(_01210_),
    .y(_03693_)
  );
  al_mux2l _09185_ (
    .a(\DFF_1094.Q ),
    .b(\DFF_98.Q ),
    .s(_03693_),
    .y(\DFF_98.D )
  );
  al_oa21ttf _09186_ (
    .a(\DFF_405.Q ),
    .b(\DFF_478.Q ),
    .c(\DFF_516.Q ),
    .y(_03694_)
  );
  al_nand3 _09187_ (
    .a(_03694_),
    .b(_01641_),
    .c(_01637_),
    .y(_03695_)
  );
  al_and3fft _09188_ (
    .a(\DFF_405.Q ),
    .b(\DFF_478.Q ),
    .c(\DFF_516.Q ),
    .y(_03696_)
  );
  al_nand3ftt _09189_ (
    .a(_03696_),
    .b(g35),
    .c(_03695_),
    .y(_03697_)
  );
  al_aoi21ftf _09190_ (
    .a(\DFF_405.Q ),
    .b(_00066_),
    .c(_03697_),
    .y(\DFF_516.D )
  );
  al_aoi21 _09191_ (
    .a(_00556_),
    .b(_00368_),
    .c(_00066_),
    .y(_03698_)
  );
  al_and3ftt _09192_ (
    .a(\DFF_244.Q ),
    .b(_02192_),
    .c(_03698_),
    .y(\DFF_244.D )
  );
  al_nand3 _09193_ (
    .a(_00499_),
    .b(_01104_),
    .c(_01787_),
    .y(_03699_)
  );
  al_ao21 _09194_ (
    .a(_01104_),
    .b(_01787_),
    .c(\DFF_1294.Q ),
    .y(_03700_)
  );
  al_nand3 _09195_ (
    .a(g35),
    .b(_03700_),
    .c(_03699_),
    .y(_03701_)
  );
  al_ao21ftf _09196_ (
    .a(g35),
    .b(\DFF_610.Q ),
    .c(_03701_),
    .y(\DFF_1294.D )
  );
  al_or2ft _09197_ (
    .a(\DFF_332.Q ),
    .b(_00373_),
    .y(_03702_)
  );
  al_inv _09198_ (
    .a(\DFF_1154.Q ),
    .y(_03703_)
  );
  al_and2ft _09199_ (
    .a(\DFF_1278.Q ),
    .b(g35),
    .y(_03704_)
  );
  al_ao21ftf _09200_ (
    .a(_03703_),
    .b(_03704_),
    .c(_01429_),
    .y(_03705_)
  );
  al_and3ftt _09201_ (
    .a(_03704_),
    .b(_03703_),
    .c(_01429_),
    .y(_03706_)
  );
  al_aoi21 _09202_ (
    .a(_03702_),
    .b(_03705_),
    .c(_03706_),
    .y(\DFF_332.D )
  );
  al_nand3fft _09203_ (
    .a(\DFF_24.Q ),
    .b(\DFF_1046.Q ),
    .c(_00718_),
    .y(_03707_)
  );
  al_ao21ftf _09204_ (
    .a(\DFF_24.Q ),
    .b(_00718_),
    .c(\DFF_1046.Q ),
    .y(_03708_)
  );
  al_nand3 _09205_ (
    .a(_03662_),
    .b(_03707_),
    .c(_03708_),
    .y(_03709_)
  );
  al_ao21 _09206_ (
    .a(_01005_),
    .b(_03662_),
    .c(\DFF_921.Q ),
    .y(_03710_)
  );
  al_nand3 _09207_ (
    .a(g35),
    .b(_03710_),
    .c(_03709_),
    .y(_03711_)
  );
  al_ao21ftf _09208_ (
    .a(_00291_),
    .b(_00066_),
    .c(_03711_),
    .y(\DFF_921.D )
  );
  al_oai21 _09209_ (
    .a(\DFF_715.Q ),
    .b(\DFF_258.Q ),
    .c(g35),
    .y(_03712_)
  );
  al_ao21ftf _09210_ (
    .a(g35),
    .b(\DFF_489.Q ),
    .c(_03712_),
    .y(\DFF_715.D )
  );
  al_or2 _09211_ (
    .a(\DFF_70.Q ),
    .b(_00846_),
    .y(_03713_)
  );
  al_nand3 _09212_ (
    .a(g35),
    .b(_00847_),
    .c(_03713_),
    .y(_03714_)
  );
  al_ao21ftf _09213_ (
    .a(g35),
    .b(\DFF_421.Q ),
    .c(_03714_),
    .y(\DFF_70.D )
  );
  al_or3ftt _09214_ (
    .a(\DFF_245.Q ),
    .b(\DFF_1408.Q ),
    .c(\DFF_199.Q ),
    .y(_03715_)
  );
  al_aoi21ftf _09215_ (
    .a(\DFF_982.Q ),
    .b(_03715_),
    .c(g35),
    .y(_03716_)
  );
  al_ao21ftf _09216_ (
    .a(_03715_),
    .b(_00499_),
    .c(_03716_),
    .y(_03717_)
  );
  al_ao21ftf _09217_ (
    .a(g35),
    .b(\DFF_72.Q ),
    .c(_03717_),
    .y(\DFF_982.D )
  );
  al_and2ft _09218_ (
    .a(g35),
    .b(\DFF_409.Q ),
    .y(_03718_)
  );
  al_ao21 _09219_ (
    .a(\DFF_318.Q ),
    .b(_00488_),
    .c(_00491_),
    .y(_03719_)
  );
  al_aoi21 _09220_ (
    .a(\DFF_318.Q ),
    .b(_00491_),
    .c(_00066_),
    .y(_03720_)
  );
  al_ao21 _09221_ (
    .a(_03719_),
    .b(_03720_),
    .c(_03718_),
    .y(\DFF_318.D )
  );
  al_aoi21ttf _09222_ (
    .a(\DFF_437.Q ),
    .b(g35),
    .c(_03490_),
    .y(_03721_)
  );
  al_or3fft _09223_ (
    .a(\DFF_437.Q ),
    .b(g35),
    .c(_03490_),
    .y(_03722_)
  );
  al_nand2ft _09224_ (
    .a(_03721_),
    .b(_03722_),
    .y(\DFF_437.D )
  );
  al_or3fft _09225_ (
    .a(\DFF_696.Q ),
    .b(g35),
    .c(_02106_),
    .y(_03723_)
  );
  al_or2 _09226_ (
    .a(\DFF_1302.Q ),
    .b(g35),
    .y(_03724_)
  );
  al_and2ft _09227_ (
    .a(\DFF_696.Q ),
    .b(g35),
    .y(_03725_)
  );
  al_ao21ttf _09228_ (
    .a(_02090_),
    .b(_02064_),
    .c(_03725_),
    .y(_03726_)
  );
  al_and3 _09229_ (
    .a(_03724_),
    .b(_03726_),
    .c(_03723_),
    .y(\DFF_696.D )
  );
  al_nand3 _09230_ (
    .a(\DFF_280.Q ),
    .b(\DFF_859.Q ),
    .c(_01593_),
    .y(_03727_)
  );
  al_nand2 _09231_ (
    .a(\DFF_339.Q ),
    .b(\DFF_859.Q ),
    .y(_03728_)
  );
  al_aoi21ftf _09232_ (
    .a(_01463_),
    .b(_03728_),
    .c(_03727_),
    .y(_03729_)
  );
  al_mux2h _09233_ (
    .a(\DFF_280.Q ),
    .b(_03729_),
    .s(g35),
    .y(\DFF_859.D )
  );
  al_ao21ftt _09234_ (
    .a(\DFF_862.Q ),
    .b(_00550_),
    .c(\DFF_811.Q ),
    .y(_03730_)
  );
  al_and2ft _09235_ (
    .a(g35),
    .b(\DFF_946.Q ),
    .y(_03731_)
  );
  al_ao21 _09236_ (
    .a(_00552_),
    .b(_03730_),
    .c(_03731_),
    .y(\DFF_811.D )
  );
  al_aoi21 _09237_ (
    .a(_00464_),
    .b(_00470_),
    .c(\DFF_922.Q ),
    .y(_03732_)
  );
  al_ao21ftf _09238_ (
    .a(_03732_),
    .b(_01864_),
    .c(_02035_),
    .y(_03733_)
  );
  al_and3ftt _09239_ (
    .a(\DFF_1199.Q ),
    .b(\DFF_892.Q ),
    .c(_00464_),
    .y(_03734_)
  );
  al_ao21 _09240_ (
    .a(_03734_),
    .b(_01865_),
    .c(_00066_),
    .y(_03735_)
  );
  al_aoi21ftf _09241_ (
    .a(\DFF_229.Q ),
    .b(_03735_),
    .c(_03733_),
    .y(\DFF_922.D )
  );
  al_ao21 _09242_ (
    .a(\DFF_936.Q ),
    .b(_01481_),
    .c(\DFF_277.Q ),
    .y(_03736_)
  );
  al_nand3 _09243_ (
    .a(_01482_),
    .b(_03736_),
    .c(_03462_),
    .y(_03737_)
  );
  al_ao21ftf _09244_ (
    .a(g35),
    .b(\DFF_936.Q ),
    .c(_03737_),
    .y(\DFF_277.D )
  );
  al_aoi21 _09245_ (
    .a(g35),
    .b(\DFF_1265.Q ),
    .c(\DFF_228.Q ),
    .y(_03738_)
  );
  al_nand3 _09246_ (
    .a(g35),
    .b(\DFF_228.Q ),
    .c(\DFF_1265.Q ),
    .y(_03739_)
  );
  al_and2ft _09247_ (
    .a(_03738_),
    .b(_03739_),
    .y(\DFF_1397.D )
  );
  al_or2 _09248_ (
    .a(\DFF_684.Q ),
    .b(_02731_),
    .y(_03740_)
  );
  al_ao21ttf _09249_ (
    .a(_01864_),
    .b(_03740_),
    .c(_02035_),
    .y(_03741_)
  );
  al_ao21 _09250_ (
    .a(_02731_),
    .b(_01865_),
    .c(_00066_),
    .y(_03742_)
  );
  al_aoi21ftf _09251_ (
    .a(\DFF_574.Q ),
    .b(_03742_),
    .c(_03741_),
    .y(\DFF_684.D )
  );
  al_mux2l _09252_ (
    .a(\DFF_544.Q ),
    .b(\DFF_239.Q ),
    .s(_01174_),
    .y(\DFF_239.D )
  );
  al_or2 _09253_ (
    .a(\DFF_175.Q ),
    .b(_01178_),
    .y(_03743_)
  );
  al_or3fft _09254_ (
    .a(_01175_),
    .b(_03743_),
    .c(_00950_),
    .y(_03744_)
  );
  al_ao21ftf _09255_ (
    .a(g35),
    .b(\DFF_876.Q ),
    .c(_03744_),
    .y(\DFF_175.D )
  );
  al_or2 _09256_ (
    .a(\DFF_1000.Q ),
    .b(\DFF_685.Q ),
    .y(_03745_)
  );
  al_mux2h _09257_ (
    .a(\DFF_25.Q ),
    .b(_03745_),
    .s(g35),
    .y(\DFF_1000.D )
  );
  al_or2ft _09258_ (
    .a(\DFF_310.Q ),
    .b(_00369_),
    .y(_03746_)
  );
  al_inv _09259_ (
    .a(\DFF_388.Q ),
    .y(_03747_)
  );
  al_ao21ftf _09260_ (
    .a(_03747_),
    .b(_01694_),
    .c(_01353_),
    .y(_03748_)
  );
  al_and3ftt _09261_ (
    .a(_01694_),
    .b(_03747_),
    .c(_01353_),
    .y(_03749_)
  );
  al_aoi21 _09262_ (
    .a(_03746_),
    .b(_03748_),
    .c(_03749_),
    .y(\DFF_310.D )
  );
  al_nand2ft _09263_ (
    .a(\DFF_1232.Q ),
    .b(\DFF_798.Q ),
    .y(_03750_)
  );
  al_nand2ft _09264_ (
    .a(\DFF_798.Q ),
    .b(\DFF_1232.Q ),
    .y(_03751_)
  );
  al_nand3 _09265_ (
    .a(g35),
    .b(_03750_),
    .c(_03751_),
    .y(_03752_)
  );
  al_aoi21ftf _09266_ (
    .a(\DFF_1161.Q ),
    .b(_00066_),
    .c(_03752_),
    .y(\DFF_1232.D )
  );
  al_or3ftt _09267_ (
    .a(g73),
    .b(\DFF_350.Q ),
    .c(g72),
    .y(_03753_)
  );
  al_mux2l _09268_ (
    .a(_03753_),
    .b(\DFF_226.Q ),
    .s(_01208_),
    .y(\DFF_56.D )
  );
  al_aoi21 _09269_ (
    .a(\DFF_1150.Q ),
    .b(g35),
    .c(\DFF_1273.Q ),
    .y(_03754_)
  );
  al_inv _09270_ (
    .a(\DFF_1273.Q ),
    .y(_03755_)
  );
  al_ao21ftf _09271_ (
    .a(_03755_),
    .b(\DFF_1150.Q ),
    .c(_01900_),
    .y(_03756_)
  );
  al_aoi21 _09272_ (
    .a(g35),
    .b(_03756_),
    .c(_03754_),
    .y(\DFF_1150.D )
  );
  al_nor2 _09273_ (
    .a(\DFF_402.Q ),
    .b(g35),
    .y(_03757_)
  );
  al_nand3 _09274_ (
    .a(\DFF_402.Q ),
    .b(_00641_),
    .c(_02348_),
    .y(_03758_)
  );
  al_oa21ftf _09275_ (
    .a(\DFF_505.Q ),
    .b(_00641_),
    .c(_00066_),
    .y(_03759_)
  );
  al_aoi21 _09276_ (
    .a(_03759_),
    .b(_03758_),
    .c(_03757_),
    .y(\DFF_505.D )
  );
  al_nand3 _09277_ (
    .a(_00499_),
    .b(_01701_),
    .c(_01773_),
    .y(_03760_)
  );
  al_ao21 _09278_ (
    .a(_01701_),
    .b(_01773_),
    .c(\DFF_392.Q ),
    .y(_03761_)
  );
  al_nand3 _09279_ (
    .a(g35),
    .b(_03761_),
    .c(_03760_),
    .y(_03762_)
  );
  al_ao21ftf _09280_ (
    .a(g35),
    .b(\DFF_151.Q ),
    .c(_03762_),
    .y(\DFF_392.D )
  );
  al_nand3 _09281_ (
    .a(_03755_),
    .b(_01764_),
    .c(_01900_),
    .y(_03763_)
  );
  al_ao21ftf _09282_ (
    .a(g35),
    .b(\DFF_584.Q ),
    .c(_03763_),
    .y(\DFF_1273.D )
  );
  al_oai21 _09283_ (
    .a(\DFF_1320.Q ),
    .b(_01502_),
    .c(_01624_),
    .y(_03764_)
  );
  al_ao21ftf _09284_ (
    .a(g35),
    .b(\DFF_22.Q ),
    .c(_03764_),
    .y(\DFF_1320.D )
  );
  al_or2ft _09285_ (
    .a(\DFF_222.Q ),
    .b(_00365_),
    .y(_03765_)
  );
  al_inv _09286_ (
    .a(\DFF_356.Q ),
    .y(_03766_)
  );
  al_ao21ftf _09287_ (
    .a(_03766_),
    .b(_03725_),
    .c(_01626_),
    .y(_03767_)
  );
  al_and3ftt _09288_ (
    .a(_03725_),
    .b(_03766_),
    .c(_01626_),
    .y(_03768_)
  );
  al_aoi21 _09289_ (
    .a(_03765_),
    .b(_03767_),
    .c(_03768_),
    .y(\DFF_222.D )
  );
  al_nor2 _09290_ (
    .a(\DFF_8.Q ),
    .b(g35),
    .y(_03769_)
  );
  al_nor3ftt _09291_ (
    .a(\DFF_725.Q ),
    .b(_02132_),
    .c(_02134_),
    .y(_03770_)
  );
  al_nand3 _09292_ (
    .a(_03770_),
    .b(_01947_),
    .c(_01943_),
    .y(_03771_)
  );
  al_oai21ttf _09293_ (
    .a(_02132_),
    .b(_02134_),
    .c(\DFF_725.Q ),
    .y(_03772_)
  );
  al_and2 _09294_ (
    .a(g35),
    .b(_03772_),
    .y(_03773_)
  );
  al_aoi21 _09295_ (
    .a(_03773_),
    .b(_03771_),
    .c(_03769_),
    .y(\DFF_725.D )
  );
  al_nand3ftt _09296_ (
    .a(_00701_),
    .b(_00499_),
    .c(_02862_),
    .y(_03774_)
  );
  al_ao21ftt _09297_ (
    .a(_00701_),
    .b(_02862_),
    .c(\DFF_267.Q ),
    .y(_03775_)
  );
  al_nand3 _09298_ (
    .a(g35),
    .b(_03774_),
    .c(_03775_),
    .y(_03776_)
  );
  al_ao21ftf _09299_ (
    .a(g35),
    .b(\DFF_519.Q ),
    .c(_03776_),
    .y(\DFF_267.D )
  );
  al_mux2h _09300_ (
    .a(\DFF_618.Q ),
    .b(_01947_),
    .s(g35),
    .y(\DFF_57.D )
  );
  al_nand3 _09301_ (
    .a(_00499_),
    .b(_01105_),
    .c(_01764_),
    .y(_03777_)
  );
  al_ao21 _09302_ (
    .a(_01105_),
    .b(_01764_),
    .c(\DFF_464.Q ),
    .y(_03778_)
  );
  al_nand3 _09303_ (
    .a(g35),
    .b(_03778_),
    .c(_03777_),
    .y(_03779_)
  );
  al_ao21ftf _09304_ (
    .a(g35),
    .b(\DFF_345.Q ),
    .c(_03779_),
    .y(\DFF_464.D )
  );
  al_or3fft _09305_ (
    .a(g25259),
    .b(_00721_),
    .c(_00725_),
    .y(_03780_)
  );
  al_ao21 _09306_ (
    .a(g25259),
    .b(_00721_),
    .c(\DFF_864.Q ),
    .y(_03781_)
  );
  al_nand3 _09307_ (
    .a(g35),
    .b(_03781_),
    .c(_03780_),
    .y(_03782_)
  );
  al_ao21ftf _09308_ (
    .a(g35),
    .b(\DFF_564.Q ),
    .c(_03782_),
    .y(\DFF_864.D )
  );
  al_mux2l _09309_ (
    .a(\DFF_1289.Q ),
    .b(\DFF_1336.Q ),
    .s(g35),
    .y(\DFF_1289.D )
  );
  al_mux2l _09310_ (
    .a(\DFF_559.Q ),
    .b(\DFF_1134.Q ),
    .s(_01016_),
    .y(\DFF_1134.D )
  );
  al_mux2l _09311_ (
    .a(\DFF_1360.Q ),
    .b(\DFF_693.Q ),
    .s(_01403_),
    .y(\DFF_693.D )
  );
  al_nor2 _09312_ (
    .a(\DFF_834.Q ),
    .b(g35),
    .y(_03783_)
  );
  al_nand3ftt _09313_ (
    .a(_03235_),
    .b(\DFF_176.Q ),
    .c(_01948_),
    .y(_03784_)
  );
  al_aoi21ftf _09314_ (
    .a(\DFF_176.Q ),
    .b(_03235_),
    .c(g35),
    .y(_03785_)
  );
  al_aoi21 _09315_ (
    .a(_03785_),
    .b(_03784_),
    .c(_03783_),
    .y(\DFF_176.D )
  );
  al_nand3 _09316_ (
    .a(_00499_),
    .b(_02367_),
    .c(_02707_),
    .y(_03786_)
  );
  al_ao21 _09317_ (
    .a(_02707_),
    .b(_02367_),
    .c(\DFF_917.Q ),
    .y(_03787_)
  );
  al_nand3 _09318_ (
    .a(g35),
    .b(_03787_),
    .c(_03786_),
    .y(_03788_)
  );
  al_ao21ftf _09319_ (
    .a(g35),
    .b(\DFF_91.Q ),
    .c(_03788_),
    .y(\DFF_917.D )
  );
  al_mux2l _09320_ (
    .a(\DFF_1336.Q ),
    .b(\DFF_15.Q ),
    .s(g35),
    .y(\DFF_1336.D )
  );
  al_oa21ftf _09321_ (
    .a(\DFF_1223.Q ),
    .b(_00604_),
    .c(_01559_),
    .y(_03789_)
  );
  al_mux2h _09322_ (
    .a(\DFF_1288.Q ),
    .b(_03789_),
    .s(_03175_),
    .y(_03790_)
  );
  al_mux2h _09323_ (
    .a(\DFF_319.Q ),
    .b(_03790_),
    .s(g35),
    .y(\DFF_1288.D )
  );
  al_mux2l _09324_ (
    .a(\DFF_213.Q ),
    .b(\DFF_1332.Q ),
    .s(_01393_),
    .y(\DFF_1332.D )
  );
  al_nor3ftt _09325_ (
    .a(\DFF_217.Q ),
    .b(_01447_),
    .c(_01450_),
    .y(_03791_)
  );
  al_oai21ttf _09326_ (
    .a(_01447_),
    .b(_01450_),
    .c(\DFF_217.Q ),
    .y(_03792_)
  );
  al_and2 _09327_ (
    .a(g35),
    .b(_03792_),
    .y(_03793_)
  );
  al_ao21ttf _09328_ (
    .a(_03791_),
    .b(_01455_),
    .c(_03793_),
    .y(_03794_)
  );
  al_aoi21ftf _09329_ (
    .a(\DFF_762.Q ),
    .b(_00066_),
    .c(_03794_),
    .y(\DFF_217.D )
  );
  al_nand3 _09330_ (
    .a(_00499_),
    .b(_01312_),
    .c(_01409_),
    .y(_03795_)
  );
  al_ao21 _09331_ (
    .a(_01312_),
    .b(_01409_),
    .c(\DFF_950.Q ),
    .y(_03796_)
  );
  al_nand3 _09332_ (
    .a(g35),
    .b(_03796_),
    .c(_03795_),
    .y(_03797_)
  );
  al_ao21ftf _09333_ (
    .a(g35),
    .b(\DFF_1186.Q ),
    .c(_03797_),
    .y(\DFF_950.D )
  );
  al_nand3 _09334_ (
    .a(\DFF_1127.Q ),
    .b(_01809_),
    .c(_00721_),
    .y(_03798_)
  );
  al_aoi21ftf _09335_ (
    .a(\DFF_564.Q ),
    .b(_03798_),
    .c(g35),
    .y(_03799_)
  );
  al_oai21 _09336_ (
    .a(_00725_),
    .b(_03798_),
    .c(_03799_),
    .y(_03800_)
  );
  al_ao21ftf _09337_ (
    .a(g35),
    .b(\DFF_32.Q ),
    .c(_03800_),
    .y(\DFF_564.D )
  );
  al_nand3fft _09338_ (
    .a(_01413_),
    .b(\DFF_1141.Q ),
    .c(_01282_),
    .y(_03801_)
  );
  al_aoi21ftf _09339_ (
    .a(\DFF_1231.Q ),
    .b(_03801_),
    .c(g35),
    .y(_03802_)
  );
  al_oai21 _09340_ (
    .a(_01284_),
    .b(_03801_),
    .c(_03802_),
    .y(_03803_)
  );
  al_ao21ftf _09341_ (
    .a(g35),
    .b(\DFF_1096.Q ),
    .c(_03803_),
    .y(\DFF_1231.D )
  );
  al_nand3 _09342_ (
    .a(\DFF_589.Q ),
    .b(g35),
    .c(_00378_),
    .y(_03804_)
  );
  al_or2 _09343_ (
    .a(\DFF_688.Q ),
    .b(g35),
    .y(_03805_)
  );
  al_or3ftt _09344_ (
    .a(g35),
    .b(\DFF_589.Q ),
    .c(_00378_),
    .y(_03806_)
  );
  al_and3 _09345_ (
    .a(_03805_),
    .b(_03804_),
    .c(_03806_),
    .y(\DFF_589.D )
  );
  al_nand3 _09346_ (
    .a(\DFF_448.Q ),
    .b(\DFF_962.Q ),
    .c(g35),
    .y(_03807_)
  );
  al_oa21 _09347_ (
    .a(g35),
    .b(\DFF_843.Q ),
    .c(_03807_),
    .y(\DFF_962.D )
  );
  al_nand3 _09348_ (
    .a(_00499_),
    .b(_01409_),
    .c(_01840_),
    .y(_03808_)
  );
  al_ao21 _09349_ (
    .a(_01409_),
    .b(_01840_),
    .c(\DFF_773.Q ),
    .y(_03809_)
  );
  al_nand3 _09350_ (
    .a(g35),
    .b(_03809_),
    .c(_03808_),
    .y(_03810_)
  );
  al_ao21ftf _09351_ (
    .a(g35),
    .b(\DFF_923.Q ),
    .c(_03810_),
    .y(\DFF_773.D )
  );
  al_ao21ftf _09352_ (
    .a(\DFF_1107.Q ),
    .b(_01986_),
    .c(_01985_),
    .y(_03811_)
  );
  al_ao21ftf _09353_ (
    .a(g35),
    .b(\DFF_985.Q ),
    .c(_03811_),
    .y(\DFF_1107.D )
  );
  al_nand3 _09354_ (
    .a(\DFF_914.Q ),
    .b(\DFF_218.Q ),
    .c(_01983_),
    .y(_03812_)
  );
  al_ao21 _09355_ (
    .a(\DFF_847.Q ),
    .b(_01989_),
    .c(\DFF_914.Q ),
    .y(_03813_)
  );
  al_nand3 _09356_ (
    .a(_03812_),
    .b(_03813_),
    .c(_01984_),
    .y(_03814_)
  );
  al_ao21ftf _09357_ (
    .a(g35),
    .b(\DFF_847.Q ),
    .c(_03814_),
    .y(\DFF_914.D )
  );
  al_or2 _09358_ (
    .a(\DFF_847.Q ),
    .b(_01989_),
    .y(_03815_)
  );
  al_and3 _09359_ (
    .a(_03812_),
    .b(_03815_),
    .c(_01984_),
    .y(_03816_)
  );
  al_ao21ttf _09360_ (
    .a(\DFF_847.Q ),
    .b(_01989_),
    .c(_03816_),
    .y(_03817_)
  );
  al_ao21ftf _09361_ (
    .a(g35),
    .b(\DFF_218.Q ),
    .c(_03817_),
    .y(\DFF_847.D )
  );
  al_oa21ttf _09362_ (
    .a(\DFF_838.Q ),
    .b(\DFF_1048.Q ),
    .c(\DFF_851.Q ),
    .y(_03818_)
  );
  al_nand3 _09363_ (
    .a(_03818_),
    .b(_00898_),
    .c(_00894_),
    .y(_03819_)
  );
  al_nand3fft _09364_ (
    .a(\DFF_838.Q ),
    .b(\DFF_1048.Q ),
    .c(\DFF_851.Q ),
    .y(_03820_)
  );
  al_nand3 _09365_ (
    .a(g35),
    .b(_03820_),
    .c(_03819_),
    .y(_03821_)
  );
  al_aoi21ftf _09366_ (
    .a(\DFF_1048.Q ),
    .b(_00066_),
    .c(_03821_),
    .y(\DFF_851.D )
  );
  al_or2 _09367_ (
    .a(\DFF_113.Q ),
    .b(_03049_),
    .y(_03822_)
  );
  al_ao21 _09368_ (
    .a(_03047_),
    .b(_03822_),
    .c(_00066_),
    .y(_03823_)
  );
  al_and2 _09369_ (
    .a(\DFF_872.Q ),
    .b(_03823_),
    .y(\DFF_113.D )
  );
  al_oa21ftf _09370_ (
    .a(\DFF_48.Q ),
    .b(\DFF_756.Q ),
    .c(\DFF_1329.Q ),
    .y(_03824_)
  );
  al_or3 _09371_ (
    .a(\DFF_48.Q ),
    .b(\DFF_760.Q ),
    .c(\DFF_1329.Q ),
    .y(_03825_)
  );
  al_or2 _09372_ (
    .a(\DFF_1149.Q ),
    .b(_03825_),
    .y(_03826_)
  );
  al_aoi21ttf _09373_ (
    .a(\DFF_756.Q ),
    .b(_01431_),
    .c(_03826_),
    .y(_03827_)
  );
  al_ao21ftf _09374_ (
    .a(_03824_),
    .b(_02255_),
    .c(_03827_),
    .y(_03828_)
  );
  al_mux2h _09375_ (
    .a(\DFF_1149.Q ),
    .b(_03828_),
    .s(g35),
    .y(\DFF_532.D )
  );
  al_nor3ftt _09376_ (
    .a(\DFF_676.Q ),
    .b(_01998_),
    .c(_01994_),
    .y(_03829_)
  );
  al_nand3 _09377_ (
    .a(_02004_),
    .b(_02006_),
    .c(_03829_),
    .y(_03830_)
  );
  al_oai21ttf _09378_ (
    .a(_01998_),
    .b(_01994_),
    .c(\DFF_676.Q ),
    .y(_03831_)
  );
  al_nand3 _09379_ (
    .a(g35),
    .b(_03831_),
    .c(_03830_),
    .y(_03832_)
  );
  al_aoi21ftf _09380_ (
    .a(\DFF_394.Q ),
    .b(_00066_),
    .c(_03832_),
    .y(\DFF_676.D )
  );
  al_mux2l _09381_ (
    .a(\DFF_1042.Q ),
    .b(\DFF_238.Q ),
    .s(_01054_),
    .y(\DFF_238.D )
  );
  al_nor2 _09382_ (
    .a(\DFF_297.Q ),
    .b(g35),
    .y(_03833_)
  );
  al_and3 _09383_ (
    .a(_00604_),
    .b(_01394_),
    .c(_00425_),
    .y(_03834_)
  );
  al_nand3ftt _09384_ (
    .a(\DFF_297.Q ),
    .b(\DFF_681.Q ),
    .c(\DFF_379.Q ),
    .y(_03835_)
  );
  al_oai21ftf _09385_ (
    .a(\DFF_681.Q ),
    .b(\DFF_297.Q ),
    .c(\DFF_379.Q ),
    .y(_03836_)
  );
  al_nand3 _09386_ (
    .a(_03835_),
    .b(_03836_),
    .c(_03834_),
    .y(_03837_)
  );
  al_oa21ftf _09387_ (
    .a(\DFF_1337.Q ),
    .b(_03834_),
    .c(_00066_),
    .y(_03838_)
  );
  al_aoi21 _09388_ (
    .a(_03837_),
    .b(_03838_),
    .c(_03833_),
    .y(\DFF_1337.D )
  );
  al_and2 _09389_ (
    .a(\DFF_1242.Q ),
    .b(g35),
    .y(\DFF_1242.D )
  );
  al_aoi21ftf _09390_ (
    .a(\DFF_525.Q ),
    .b(_02024_),
    .c(_02027_),
    .y(_03839_)
  );
  al_ao21ftf _09391_ (
    .a(_02024_),
    .b(\DFF_525.Q ),
    .c(_03839_),
    .y(_03840_)
  );
  al_ao21ftf _09392_ (
    .a(g35),
    .b(\DFF_870.Q ),
    .c(_03840_),
    .y(\DFF_525.D )
  );
  al_nor2 _09393_ (
    .a(g35),
    .b(\DFF_1089.Q ),
    .y(_03841_)
  );
  al_nand3 _09394_ (
    .a(\DFF_1054.Q ),
    .b(_00721_),
    .c(_01707_),
    .y(_03842_)
  );
  al_oa21ftf _09395_ (
    .a(\DFF_1127.Q ),
    .b(_00721_),
    .c(_00066_),
    .y(_03843_)
  );
  al_aoi21 _09396_ (
    .a(_03843_),
    .b(_03842_),
    .c(_03841_),
    .y(\DFF_1127.D )
  );
  al_and2ft _09397_ (
    .a(g35),
    .b(\DFF_1143.Q ),
    .y(_03844_)
  );
  al_and3ftt _09398_ (
    .a(_00973_),
    .b(_00604_),
    .c(_02882_),
    .y(_03845_)
  );
  al_oai21ftt _09399_ (
    .a(\DFF_886.Q ),
    .b(\DFF_265.Q ),
    .c(\DFF_1181.Q ),
    .y(_03846_)
  );
  al_nand2ft _09400_ (
    .a(\DFF_1181.Q ),
    .b(_00329_),
    .y(_03847_)
  );
  al_nand3 _09401_ (
    .a(_03846_),
    .b(_03847_),
    .c(_03845_),
    .y(_03848_)
  );
  al_oa21ttf _09402_ (
    .a(\DFF_1254.Q ),
    .b(_03845_),
    .c(_00066_),
    .y(_03849_)
  );
  al_ao21 _09403_ (
    .a(_03848_),
    .b(_03849_),
    .c(_03844_),
    .y(\DFF_1254.D )
  );
  al_mux2l _09404_ (
    .a(\DFF_656.Q ),
    .b(\DFF_135.Q ),
    .s(_01054_),
    .y(\DFF_135.D )
  );
  al_mux2l _09405_ (
    .a(\DFF_689.Q ),
    .b(\DFF_1230.Q ),
    .s(_03057_),
    .y(_03850_)
  );
  al_mux2h _09406_ (
    .a(\DFF_1139.Q ),
    .b(_03850_),
    .s(g35),
    .y(\DFF_689.D )
  );
  al_oa21ftf _09407_ (
    .a(\DFF_768.Q ),
    .b(_02045_),
    .c(_00066_),
    .y(_03851_)
  );
  al_ao21ftf _09408_ (
    .a(\DFF_768.Q ),
    .b(_02045_),
    .c(_03851_),
    .y(_03852_)
  );
  al_aoi21ftf _09409_ (
    .a(\DFF_488.Q ),
    .b(_00066_),
    .c(_03852_),
    .y(\DFF_768.D )
  );
  al_ao21 _09410_ (
    .a(\DFF_953.Q ),
    .b(_00953_),
    .c(\DFF_1200.Q ),
    .y(_03853_)
  );
  al_nand3fft _09411_ (
    .a(_01837_),
    .b(_00954_),
    .c(_03853_),
    .y(_03854_)
  );
  al_ao21ftf _09412_ (
    .a(g35),
    .b(\DFF_953.Q ),
    .c(_03854_),
    .y(\DFF_1200.D )
  );
  al_ao21 _09413_ (
    .a(_02090_),
    .b(_02064_),
    .c(_00066_),
    .y(_03855_)
  );
  al_mux2l _09414_ (
    .a(\DFF_1342.Q ),
    .b(\DFF_1358.Q ),
    .s(_03855_),
    .y(\DFF_1358.D )
  );
  al_and2ft _09415_ (
    .a(g35),
    .b(\DFF_866.Q ),
    .y(_03856_)
  );
  al_ao21ftt _09416_ (
    .a(_00871_),
    .b(_01050_),
    .c(\DFF_902.Q ),
    .y(_03857_)
  );
  al_and2ft _09417_ (
    .a(_01597_),
    .b(_03857_),
    .y(_03858_)
  );
  al_ao21 _09418_ (
    .a(_03858_),
    .b(_01607_),
    .c(_03856_),
    .y(\DFF_902.D )
  );
  al_nand3fft _09419_ (
    .a(\DFF_271.Q ),
    .b(\DFF_522.Q ),
    .c(\DFF_54.Q ),
    .y(_03859_)
  );
  al_aoi21ftf _09420_ (
    .a(\DFF_1263.Q ),
    .b(_03859_),
    .c(g35),
    .y(_03860_)
  );
  al_ao21ftf _09421_ (
    .a(_03859_),
    .b(_00499_),
    .c(_03860_),
    .y(_03861_)
  );
  al_ao21ftf _09422_ (
    .a(g35),
    .b(\DFF_670.Q ),
    .c(_03861_),
    .y(\DFF_1263.D )
  );
  al_ao21 _09423_ (
    .a(g35),
    .b(\DFF_124.Q ),
    .c(\DFF_1372.Q ),
    .y(_03862_)
  );
  al_aoi21 _09424_ (
    .a(g35),
    .b(_02106_),
    .c(_03862_),
    .y(_03863_)
  );
  al_ao21ttf _09425_ (
    .a(_02090_),
    .b(_02064_),
    .c(\DFF_1409.Q ),
    .y(_03864_)
  );
  al_nand2 _09426_ (
    .a(\DFF_1372.Q ),
    .b(\DFF_124.Q ),
    .y(_03865_)
  );
  al_oa21ftf _09427_ (
    .a(_03865_),
    .b(_02106_),
    .c(_00066_),
    .y(_03866_)
  );
  al_aoi21 _09428_ (
    .a(_03864_),
    .b(_03866_),
    .c(_03863_),
    .y(\DFF_1409.D )
  );
  al_and2ft _09429_ (
    .a(g35),
    .b(\DFF_690.Q ),
    .y(_03867_)
  );
  al_nand2 _09430_ (
    .a(_01085_),
    .b(_01087_),
    .y(_03868_)
  );
  al_ao21ftf _09431_ (
    .a(_01090_),
    .b(\DFF_690.Q ),
    .c(_03868_),
    .y(_03869_)
  );
  al_ao21ttf _09432_ (
    .a(\DFF_1327.Q ),
    .b(_01101_),
    .c(_03869_),
    .y(_03870_)
  );
  al_oa21ftf _09433_ (
    .a(\DFF_1327.Q ),
    .b(_03869_),
    .c(_00066_),
    .y(_03871_)
  );
  al_ao21 _09434_ (
    .a(_03871_),
    .b(_03870_),
    .c(_03867_),
    .y(\DFF_1327.D )
  );
  al_mux2h _09435_ (
    .a(\DFF_1363.Q ),
    .b(_01934_),
    .s(g26801),
    .y(_03872_)
  );
  al_mux2h _09436_ (
    .a(\DFF_497.Q ),
    .b(_03872_),
    .s(g35),
    .y(\DFF_1363.D )
  );
  al_or3fft _09437_ (
    .a(_00335_),
    .b(_01889_),
    .c(_01892_),
    .y(_03873_)
  );
  al_ao21 _09438_ (
    .a(_00335_),
    .b(_01889_),
    .c(\DFF_1137.Q ),
    .y(_03874_)
  );
  al_nand3 _09439_ (
    .a(g35),
    .b(_03874_),
    .c(_03873_),
    .y(_03875_)
  );
  al_ao21ftf _09440_ (
    .a(g35),
    .b(\DFF_16.Q ),
    .c(_03875_),
    .y(\DFF_1137.D )
  );
  al_nand3ftt _09441_ (
    .a(_01151_),
    .b(_00439_),
    .c(_01363_),
    .y(_03876_)
  );
  al_ao21 _09442_ (
    .a(_00439_),
    .b(_01363_),
    .c(\DFF_862.Q ),
    .y(_03877_)
  );
  al_nand3 _09443_ (
    .a(g35),
    .b(_03876_),
    .c(_03877_),
    .y(_03878_)
  );
  al_ao21ftf _09444_ (
    .a(g35),
    .b(\DFF_465.Q ),
    .c(_03878_),
    .y(\DFF_862.D )
  );
  al_mux2l _09445_ (
    .a(\DFF_1045.Q ),
    .b(\DFF_292.Q ),
    .s(_01109_),
    .y(\DFF_292.D )
  );
  al_aoi21 _09446_ (
    .a(\DFF_664.Q ),
    .b(_01622_),
    .c(_00066_),
    .y(_03879_)
  );
  al_nand2ft _09447_ (
    .a(g35),
    .b(\DFF_664.Q ),
    .y(_03880_)
  );
  al_ao21ftf _09448_ (
    .a(\DFF_39.Q ),
    .b(_03879_),
    .c(_03880_),
    .y(\DFF_1214.D )
  );
  al_mux2l _09449_ (
    .a(\DFF_5.Q ),
    .b(\DFF_478.Q ),
    .s(g35),
    .y(\DFF_460.D )
  );
  al_nand3ftt _09450_ (
    .a(\DFF_68.Q ),
    .b(\DFF_598.Q ),
    .c(\DFF_1098.Q ),
    .y(_03881_)
  );
  al_aoi21ftf _09451_ (
    .a(\DFF_750.Q ),
    .b(_03881_),
    .c(g35),
    .y(_03882_)
  );
  al_ao21ftf _09452_ (
    .a(_03881_),
    .b(_00499_),
    .c(_03882_),
    .y(_03883_)
  );
  al_ao21ftf _09453_ (
    .a(g35),
    .b(\DFF_187.Q ),
    .c(_03883_),
    .y(\DFF_750.D )
  );
  al_nand3fft _09454_ (
    .a(\DFF_402.Q ),
    .b(_01614_),
    .c(_00641_),
    .y(_03884_)
  );
  al_aoi21ftf _09455_ (
    .a(\DFF_61.Q ),
    .b(_03884_),
    .c(g35),
    .y(_03885_)
  );
  al_ao21ftf _09456_ (
    .a(_03884_),
    .b(_01618_),
    .c(_03885_),
    .y(_03886_)
  );
  al_ao21ftf _09457_ (
    .a(g35),
    .b(\DFF_727.Q ),
    .c(_03886_),
    .y(\DFF_61.D )
  );
  al_and3ftt _09458_ (
    .a(\DFF_174.Q ),
    .b(\DFF_968.Q ),
    .c(\DFF_705.Q ),
    .y(_03887_)
  );
  al_and3ftt _09459_ (
    .a(\DFF_174.Q ),
    .b(\DFF_1422.Q ),
    .c(\DFF_103.Q ),
    .y(_03888_)
  );
  al_ao21 _09460_ (
    .a(\DFF_504.Q ),
    .b(_00431_),
    .c(_03888_),
    .y(_03889_)
  );
  al_and3ftt _09461_ (
    .a(\DFF_705.Q ),
    .b(\DFF_174.Q ),
    .c(\DFF_973.Q ),
    .y(_03890_)
  );
  al_nand3 _09462_ (
    .a(\DFF_1172.Q ),
    .b(\DFF_103.Q ),
    .c(\DFF_705.Q ),
    .y(_03891_)
  );
  al_nand3fft _09463_ (
    .a(\DFF_103.Q ),
    .b(\DFF_705.Q ),
    .c(\DFF_2.Q ),
    .y(_03892_)
  );
  al_and3ftt _09464_ (
    .a(_03890_),
    .b(_03891_),
    .c(_03892_),
    .y(_03893_)
  );
  al_nand3fft _09465_ (
    .a(_03887_),
    .b(_03889_),
    .c(_03893_),
    .y(_03894_)
  );
  al_mux2l _09466_ (
    .a(_03894_),
    .b(\DFF_772.Q ),
    .s(_02775_),
    .y(_03895_)
  );
  al_mux2h _09467_ (
    .a(\DFF_103.Q ),
    .b(_03895_),
    .s(g35),
    .y(\DFF_772.D )
  );
  al_nor2 _09468_ (
    .a(g35),
    .b(\DFF_1009.Q ),
    .y(_03896_)
  );
  al_nand3 _09469_ (
    .a(\DFF_111.Q ),
    .b(_01125_),
    .c(_01531_),
    .y(_03897_)
  );
  al_oa21ftf _09470_ (
    .a(\DFF_759.Q ),
    .b(_01125_),
    .c(_00066_),
    .y(_03898_)
  );
  al_aoi21 _09471_ (
    .a(_03898_),
    .b(_03897_),
    .c(_03896_),
    .y(\DFF_759.D )
  );
  al_nand3 _09472_ (
    .a(_00498_),
    .b(_00499_),
    .c(_01773_),
    .y(_03899_)
  );
  al_ao21 _09473_ (
    .a(_00498_),
    .b(_01773_),
    .c(\DFF_476.Q ),
    .y(_03900_)
  );
  al_nand3 _09474_ (
    .a(g35),
    .b(_03900_),
    .c(_03899_),
    .y(_03901_)
  );
  al_ao21ftf _09475_ (
    .a(g35),
    .b(\DFF_938.Q ),
    .c(_03901_),
    .y(\DFF_476.D )
  );
  al_and3ftt _09476_ (
    .a(\DFF_1148.Q ),
    .b(\DFF_717.Q ),
    .c(\DFF_327.Q ),
    .y(_03902_)
  );
  al_and3 _09477_ (
    .a(\DFF_193.Q ),
    .b(_03902_),
    .c(_01261_),
    .y(_03903_)
  );
  al_oa21ftf _09478_ (
    .a(_02795_),
    .b(_03903_),
    .c(_00066_),
    .y(_03904_)
  );
  al_ao21ftf _09479_ (
    .a(_02795_),
    .b(_03903_),
    .c(_03904_),
    .y(_03905_)
  );
  al_ao21ftf _09480_ (
    .a(g35),
    .b(\DFF_193.Q ),
    .c(_03905_),
    .y(\DFF_403.D )
  );
  al_nand3 _09481_ (
    .a(_00499_),
    .b(_00509_),
    .c(_01764_),
    .y(_03906_)
  );
  al_ao21 _09482_ (
    .a(_00509_),
    .b(_01764_),
    .c(\DFF_617.Q ),
    .y(_03907_)
  );
  al_nand3 _09483_ (
    .a(g35),
    .b(_03907_),
    .c(_03906_),
    .y(_03908_)
  );
  al_ao21ftf _09484_ (
    .a(g35),
    .b(\DFF_419.Q ),
    .c(_03908_),
    .y(\DFF_617.D )
  );
  al_mux2l _09485_ (
    .a(\DFF_580.Q ),
    .b(\DFF_1094.Q ),
    .s(_03693_),
    .y(\DFF_1094.D )
  );
  al_and2 _09486_ (
    .a(g35),
    .b(\DFF_663.Q ),
    .y(\DFF_929.D )
  );
  al_nand3fft _09487_ (
    .a(\DFF_1127.Q ),
    .b(_01810_),
    .c(_00721_),
    .y(_03909_)
  );
  al_aoi21ftf _09488_ (
    .a(\DFF_32.Q ),
    .b(_03909_),
    .c(g35),
    .y(_03910_)
  );
  al_oai21 _09489_ (
    .a(_00725_),
    .b(_03909_),
    .c(_03910_),
    .y(_03911_)
  );
  al_ao21ftf _09490_ (
    .a(g35),
    .b(\DFF_246.Q ),
    .c(_03911_),
    .y(\DFF_32.D )
  );
  al_oa21ftt _09491_ (
    .a(g35),
    .b(\DFF_1239.Q ),
    .c(\DFF_513.Q ),
    .y(\DFF_1405.D )
  );
  al_inv _09492_ (
    .a(_00758_),
    .y(_03912_)
  );
  al_nand3 _09493_ (
    .a(_03551_),
    .b(_00758_),
    .c(_02449_),
    .y(_03913_)
  );
  al_aoi21ftf _09494_ (
    .a(\DFF_562.Q ),
    .b(_03912_),
    .c(_03913_),
    .y(_03914_)
  );
  al_mux2h _09495_ (
    .a(\DFF_581.Q ),
    .b(_03914_),
    .s(g35),
    .y(\DFF_562.D )
  );
  al_nand3 _09496_ (
    .a(_00499_),
    .b(_01169_),
    .c(_02930_),
    .y(_03915_)
  );
  al_ao21 _09497_ (
    .a(_01169_),
    .b(_02930_),
    .c(\DFF_397.Q ),
    .y(_03916_)
  );
  al_nand3 _09498_ (
    .a(g35),
    .b(_03916_),
    .c(_03915_),
    .y(_03917_)
  );
  al_ao21ftf _09499_ (
    .a(g35),
    .b(\DFF_1011.Q ),
    .c(_03917_),
    .y(\DFF_397.D )
  );
  al_mux2l _09500_ (
    .a(\DFF_1042.Q ),
    .b(\DFF_1164.Q ),
    .s(_01053_),
    .y(_03918_)
  );
  al_and2 _09501_ (
    .a(g35),
    .b(_03918_),
    .y(\DFF_1042.D )
  );
  al_nand3ftt _09502_ (
    .a(_02806_),
    .b(_00426_),
    .c(_01394_),
    .y(_03919_)
  );
  al_ao21 _09503_ (
    .a(_00426_),
    .b(_01394_),
    .c(\DFF_1240.Q ),
    .y(_03920_)
  );
  al_nand3 _09504_ (
    .a(g35),
    .b(_03919_),
    .c(_03920_),
    .y(_03921_)
  );
  al_ao21ftf _09505_ (
    .a(g35),
    .b(\DFF_457.Q ),
    .c(_03921_),
    .y(\DFF_1240.D )
  );
  al_and2 _09506_ (
    .a(\DFF_1415.Q ),
    .b(\DFF_79.Q ),
    .y(_03922_)
  );
  al_nand3ftt _09507_ (
    .a(\DFF_79.Q ),
    .b(_01721_),
    .c(_01720_),
    .y(_03923_)
  );
  al_nand3fft _09508_ (
    .a(_00066_),
    .b(_03922_),
    .c(_03923_),
    .y(_03924_)
  );
  al_aoi21ftf _09509_ (
    .a(\DFF_813.Q ),
    .b(_00066_),
    .c(_03924_),
    .y(\DFF_1415.D )
  );
  al_aoi21 _09510_ (
    .a(\DFF_522.Q ),
    .b(g35),
    .c(\DFF_54.Q ),
    .y(_03925_)
  );
  al_ao21ftf _09511_ (
    .a(_01358_),
    .b(\DFF_522.Q ),
    .c(_01359_),
    .y(_03926_)
  );
  al_aoi21 _09512_ (
    .a(g35),
    .b(_03926_),
    .c(_03925_),
    .y(\DFF_522.D )
  );
  al_mux2l _09513_ (
    .a(\DFF_1376.Q ),
    .b(\DFF_77.Q ),
    .s(_01592_),
    .y(\DFF_77.D )
  );
  al_nand3ftt _09514_ (
    .a(_02030_),
    .b(_00499_),
    .c(_01045_),
    .y(_03927_)
  );
  al_ao21ftt _09515_ (
    .a(_02030_),
    .b(_01045_),
    .c(\DFF_1259.Q ),
    .y(_03928_)
  );
  al_nand3 _09516_ (
    .a(g35),
    .b(_03927_),
    .c(_03928_),
    .y(_03929_)
  );
  al_ao21ftf _09517_ (
    .a(g35),
    .b(\DFF_19.Q ),
    .c(_03929_),
    .y(\DFF_1259.D )
  );
  al_oai21 _09518_ (
    .a(\DFF_197.Q ),
    .b(\DFF_1074.Q ),
    .c(g35),
    .y(_03930_)
  );
  al_ao21ftf _09519_ (
    .a(g35),
    .b(\DFF_242.Q ),
    .c(_03930_),
    .y(\DFF_197.D )
  );
  al_mux2l _09520_ (
    .a(_01186_),
    .b(_01232_),
    .s(_01187_),
    .y(_03931_)
  );
  al_mux2h _09521_ (
    .a(\DFF_560.Q ),
    .b(_03931_),
    .s(g35),
    .y(\DFF_863.D )
  );
  al_nor2 _09522_ (
    .a(g35),
    .b(\DFF_1348.Q ),
    .y(_03932_)
  );
  al_nand2 _09523_ (
    .a(\DFF_1158.Q ),
    .b(\DFF_1169.Q ),
    .y(_03933_)
  );
  al_nand2 _09524_ (
    .a(\DFF_1294.Q ),
    .b(\DFF_971.Q ),
    .y(_03934_)
  );
  al_aoi21ttf _09525_ (
    .a(_03933_),
    .b(_03934_),
    .c(_00412_),
    .y(_03935_)
  );
  al_nand2ft _09526_ (
    .a(\DFF_878.Q ),
    .b(\DFF_952.Q ),
    .y(_03936_)
  );
  al_nand2 _09527_ (
    .a(\DFF_1185.Q ),
    .b(\DFF_1175.Q ),
    .y(_03937_)
  );
  al_nand2 _09528_ (
    .a(\DFF_378.Q ),
    .b(\DFF_780.Q ),
    .y(_03938_)
  );
  al_ao21 _09529_ (
    .a(_03937_),
    .b(_03938_),
    .c(_03936_),
    .y(_03939_)
  );
  al_and3fft _09530_ (
    .a(\DFF_952.Q ),
    .b(\DFF_878.Q ),
    .c(\DFF_836.Q ),
    .y(_03940_)
  );
  al_ao21 _09531_ (
    .a(\DFF_1120.Q ),
    .b(_03940_),
    .c(\DFF_198.Q ),
    .y(_03941_)
  );
  al_nand2ft _09532_ (
    .a(\DFF_952.Q ),
    .b(\DFF_878.Q ),
    .y(_03942_)
  );
  al_nand2 _09533_ (
    .a(\DFF_1024.Q ),
    .b(\DFF_1023.Q ),
    .y(_03943_)
  );
  al_nand2 _09534_ (
    .a(\DFF_610.Q ),
    .b(\DFF_163.Q ),
    .y(_03944_)
  );
  al_ao21 _09535_ (
    .a(_03943_),
    .b(_03944_),
    .c(_03942_),
    .y(_03945_)
  );
  al_and3ftt _09536_ (
    .a(_03941_),
    .b(_03939_),
    .c(_03945_),
    .y(_03946_)
  );
  al_nand3 _09537_ (
    .a(\DFF_617.Q ),
    .b(\DFF_780.Q ),
    .c(_00412_),
    .y(_03947_)
  );
  al_or3fft _09538_ (
    .a(\DFF_419.Q ),
    .b(\DFF_836.Q ),
    .c(_03942_),
    .y(_03948_)
  );
  al_and3 _09539_ (
    .a(\DFF_198.Q ),
    .b(_03948_),
    .c(_03947_),
    .y(_03949_)
  );
  al_nor2 _09540_ (
    .a(\DFF_952.Q ),
    .b(\DFF_878.Q ),
    .y(_03950_)
  );
  al_nand2 _09541_ (
    .a(\DFF_1174.Q ),
    .b(\DFF_163.Q ),
    .y(_03951_)
  );
  al_nand2 _09542_ (
    .a(\DFF_967.Q ),
    .b(\DFF_1023.Q ),
    .y(_03952_)
  );
  al_ao21ttf _09543_ (
    .a(_03951_),
    .b(_03952_),
    .c(_03950_),
    .y(_03953_)
  );
  al_nand2 _09544_ (
    .a(\DFF_957.Q ),
    .b(\DFF_971.Q ),
    .y(_03954_)
  );
  al_nand2 _09545_ (
    .a(\DFF_1158.Q ),
    .b(\DFF_1032.Q ),
    .y(_03955_)
  );
  al_ao21 _09546_ (
    .a(_03954_),
    .b(_03955_),
    .c(_03936_),
    .y(_03956_)
  );
  al_nand3 _09547_ (
    .a(_03953_),
    .b(_03956_),
    .c(_03949_),
    .y(_03957_)
  );
  al_ao21ftf _09548_ (
    .a(_03935_),
    .b(_03946_),
    .c(_03957_),
    .y(_03958_)
  );
  al_nand2 _09549_ (
    .a(\DFF_1348.Q ),
    .b(_02339_),
    .y(_03959_)
  );
  al_nor3fft _09550_ (
    .a(\DFF_1196.Q ),
    .b(\DFF_291.Q ),
    .c(_03936_),
    .y(_03960_)
  );
  al_nor3fft _09551_ (
    .a(\DFF_1248.Q ),
    .b(\DFF_779.Q ),
    .c(_03942_),
    .y(_03961_)
  );
  al_nor2 _09552_ (
    .a(\DFF_1158.Q ),
    .b(\DFF_198.Q ),
    .y(_03962_)
  );
  al_nand2 _09553_ (
    .a(\DFF_1158.Q ),
    .b(\DFF_198.Q ),
    .y(_03963_)
  );
  al_nand3 _09554_ (
    .a(\DFF_806.Q ),
    .b(\DFF_588.Q ),
    .c(_03950_),
    .y(_03964_)
  );
  al_and3ftt _09555_ (
    .a(_03962_),
    .b(_03963_),
    .c(_03964_),
    .y(_03965_)
  );
  al_nand3fft _09556_ (
    .a(_03960_),
    .b(_03961_),
    .c(_03965_),
    .y(_03966_)
  );
  al_and3 _09557_ (
    .a(\DFF_1196.Q ),
    .b(\DFF_345.Q ),
    .c(_00412_),
    .y(_03967_)
  );
  al_nand2ft _09558_ (
    .a(_03962_),
    .b(_03963_),
    .y(_03968_)
  );
  al_or3fft _09559_ (
    .a(\DFF_806.Q ),
    .b(\DFF_730.Q ),
    .c(_03942_),
    .y(_03969_)
  );
  al_and3 _09560_ (
    .a(\DFF_1248.Q ),
    .b(\DFF_464.Q ),
    .c(_03950_),
    .y(_03970_)
  );
  al_and3ftt _09561_ (
    .a(_03970_),
    .b(_03969_),
    .c(_03968_),
    .y(_03971_)
  );
  al_ao21ftf _09562_ (
    .a(_03967_),
    .b(_03971_),
    .c(_03966_),
    .y(_03972_)
  );
  al_nand3 _09563_ (
    .a(_03959_),
    .b(_03972_),
    .c(_03958_),
    .y(_03973_)
  );
  al_nand2 _09564_ (
    .a(_02338_),
    .b(_03973_),
    .y(_03974_)
  );
  al_oa21ftf _09565_ (
    .a(\DFF_714.Q ),
    .b(_02338_),
    .c(_00066_),
    .y(_03975_)
  );
  al_aoi21 _09566_ (
    .a(_03975_),
    .b(_03974_),
    .c(_03932_),
    .y(\DFF_714.D )
  );
  al_mux2h _09567_ (
    .a(\DFF_669.Q ),
    .b(_00309_),
    .s(\DFF_799.Q ),
    .y(_03976_)
  );
  al_mux2h _09568_ (
    .a(\DFF_736.Q ),
    .b(_03976_),
    .s(g35),
    .y(\DFF_669.D )
  );
  al_ao21 _09569_ (
    .a(\DFF_978.Q ),
    .b(g35),
    .c(_03315_),
    .y(_03977_)
  );
  al_and3 _09570_ (
    .a(\DFF_978.Q ),
    .b(g35),
    .c(_03315_),
    .y(_03978_)
  );
  al_and2ft _09571_ (
    .a(_03978_),
    .b(_03977_),
    .y(\DFF_978.D )
  );
  al_mux2l _09572_ (
    .a(\DFF_1164.Q ),
    .b(\DFF_1003.Q ),
    .s(_01557_),
    .y(_03979_)
  );
  al_mux2h _09573_ (
    .a(\DFF_346.Q ),
    .b(_03979_),
    .s(g35),
    .y(\DFF_1164.D )
  );
  al_nand3 _09574_ (
    .a(_00499_),
    .b(_01497_),
    .c(_02011_),
    .y(_03980_)
  );
  al_ao21 _09575_ (
    .a(_01497_),
    .b(_02011_),
    .c(\DFF_633.Q ),
    .y(_03981_)
  );
  al_nand3 _09576_ (
    .a(g35),
    .b(_03981_),
    .c(_03980_),
    .y(_03982_)
  );
  al_ao21ftf _09577_ (
    .a(g35),
    .b(\DFF_227.Q ),
    .c(_03982_),
    .y(\DFF_633.D )
  );
  al_or3fft _09578_ (
    .a(_01575_),
    .b(_01889_),
    .c(_01892_),
    .y(_03983_)
  );
  al_ao21 _09579_ (
    .a(_01575_),
    .b(_01889_),
    .c(\DFF_173.Q ),
    .y(_03984_)
  );
  al_nand3 _09580_ (
    .a(g35),
    .b(_03984_),
    .c(_03983_),
    .y(_03985_)
  );
  al_ao21ftf _09581_ (
    .a(g35),
    .b(\DFF_1137.Q ),
    .c(_03985_),
    .y(\DFF_173.D )
  );
  al_nand2 _09582_ (
    .a(\DFF_343.Q ),
    .b(_01123_),
    .y(_03986_)
  );
  al_oai21ftt _09583_ (
    .a(_03986_),
    .b(_01130_),
    .c(_01125_),
    .y(_03987_)
  );
  al_ao21 _09584_ (
    .a(\DFF_455.Q ),
    .b(_01126_),
    .c(_03987_),
    .y(_03988_)
  );
  al_nand3 _09585_ (
    .a(\DFF_455.Q ),
    .b(_01126_),
    .c(_03987_),
    .y(_03989_)
  );
  al_nand3 _09586_ (
    .a(g35),
    .b(_03989_),
    .c(_03988_),
    .y(_03990_)
  );
  al_aoi21ftf _09587_ (
    .a(\DFF_620.Q ),
    .b(_00066_),
    .c(_03990_),
    .y(\DFF_455.D )
  );
  al_and2 _09588_ (
    .a(\DFF_587.Q ),
    .b(g35),
    .y(\DFF_147.D )
  );
  al_nand3 _09589_ (
    .a(\DFF_434.Q ),
    .b(\DFF_891.Q ),
    .c(g35),
    .y(_03991_)
  );
  al_oa21 _09590_ (
    .a(g35),
    .b(\DFF_685.Q ),
    .c(_03991_),
    .y(\DFF_891.D )
  );
  al_mux2h _09591_ (
    .a(\DFF_1389.Q ),
    .b(_00868_),
    .s(g35),
    .y(\DFF_389.D )
  );
  al_nand2ft _09592_ (
    .a(\DFF_737.Q ),
    .b(\DFF_1087.Q ),
    .y(_03992_)
  );
  al_oai21ttf _09593_ (
    .a(\DFF_326.Q ),
    .b(\DFF_797.Q ),
    .c(_01501_),
    .y(_03993_)
  );
  al_or2 _09594_ (
    .a(\DFF_110.Q ),
    .b(\DFF_737.Q ),
    .y(_03994_)
  );
  al_ao21ttf _09595_ (
    .a(\DFF_797.Q ),
    .b(\DFF_110.Q ),
    .c(_03994_),
    .y(_03995_)
  );
  al_and3 _09596_ (
    .a(_03992_),
    .b(_03995_),
    .c(_03993_),
    .y(_03996_)
  );
  al_and3ftt _09597_ (
    .a(_01502_),
    .b(g35),
    .c(_03996_),
    .y(\DFF_30.D )
  );
  al_mux2l _09598_ (
    .a(\DFF_696.Q ),
    .b(\DFF_356.Q ),
    .s(_01626_),
    .y(\DFF_356.D )
  );
  al_and3ftt _09599_ (
    .a(\DFF_410.Q ),
    .b(_03755_),
    .c(_01923_),
    .y(\DFF_410.D )
  );
  al_mux2l _09600_ (
    .a(_01284_),
    .b(\DFF_1096.Q ),
    .s(_01858_),
    .y(_03997_)
  );
  al_mux2h _09601_ (
    .a(\DFF_1050.Q ),
    .b(_03997_),
    .s(g35),
    .y(\DFF_1096.D )
  );
  al_nand2 _09602_ (
    .a(\DFF_1306.Q ),
    .b(\DFF_632.Q ),
    .y(_03998_)
  );
  al_nor2 _09603_ (
    .a(\DFF_1306.Q ),
    .b(\DFF_632.Q ),
    .y(_03999_)
  );
  al_nand2ft _09604_ (
    .a(_03999_),
    .b(_03998_),
    .y(_04000_)
  );
  al_mux2l _09605_ (
    .a(\DFF_361.Q ),
    .b(_04000_),
    .s(_01958_),
    .y(_04001_)
  );
  al_mux2h _09606_ (
    .a(\DFF_632.Q ),
    .b(_04001_),
    .s(g35),
    .y(\DFF_361.D )
  );
  al_mux2l _09607_ (
    .a(\DFF_1278.Q ),
    .b(\DFF_1154.Q ),
    .s(_01429_),
    .y(\DFF_1154.D )
  );
  al_and2ft _09608_ (
    .a(g35),
    .b(\DFF_272.Q ),
    .y(_04002_)
  );
  al_and3ftt _09609_ (
    .a(_01888_),
    .b(_00604_),
    .c(_00334_),
    .y(_04003_)
  );
  al_oai21ftt _09610_ (
    .a(\DFF_18.Q ),
    .b(\DFF_500.Q ),
    .c(\DFF_1181.Q ),
    .y(_04004_)
  );
  al_nand2ft _09611_ (
    .a(\DFF_1181.Q ),
    .b(_00335_),
    .y(_04005_)
  );
  al_nand3 _09612_ (
    .a(_04004_),
    .b(_04005_),
    .c(_04003_),
    .y(_04006_)
  );
  al_oa21ftf _09613_ (
    .a(_03059_),
    .b(_04003_),
    .c(_00066_),
    .y(_04007_)
  );
  al_ao21 _09614_ (
    .a(_04006_),
    .b(_04007_),
    .c(_04002_),
    .y(\DFF_567.D )
  );
  al_ao21 _09615_ (
    .a(_00758_),
    .b(_02449_),
    .c(_00066_),
    .y(_04008_)
  );
  al_and3fft _09616_ (
    .a(_00066_),
    .b(_00758_),
    .c(_03551_),
    .y(_04009_)
  );
  al_aoi21 _09617_ (
    .a(_02452_),
    .b(_04008_),
    .c(_04009_),
    .y(\DFF_189.D )
  );
  al_oa21ttf _09618_ (
    .a(\DFF_1075.Q ),
    .b(_01890_),
    .c(_00066_),
    .y(_04010_)
  );
  al_ao21ttf _09619_ (
    .a(\DFF_1075.Q ),
    .b(_01890_),
    .c(_04010_),
    .y(_04011_)
  );
  al_ao21ftf _09620_ (
    .a(g35),
    .b(\DFF_814.Q ),
    .c(_04011_),
    .y(\DFF_1075.D )
  );
  al_nor2 _09621_ (
    .a(\DFF_475.Q ),
    .b(g35),
    .y(_04012_)
  );
  al_nor3ftt _09622_ (
    .a(\DFF_741.Q ),
    .b(_01631_),
    .c(_01628_),
    .y(_04013_)
  );
  al_nand3 _09623_ (
    .a(_04013_),
    .b(_01641_),
    .c(_01637_),
    .y(_04014_)
  );
  al_oai21ttf _09624_ (
    .a(_01631_),
    .b(_01628_),
    .c(\DFF_741.Q ),
    .y(_04015_)
  );
  al_and2 _09625_ (
    .a(g35),
    .b(_04015_),
    .y(_04016_)
  );
  al_aoi21 _09626_ (
    .a(_04016_),
    .b(_04014_),
    .c(_04012_),
    .y(\DFF_741.D )
  );
  al_nor2 _09627_ (
    .a(\DFF_95.Q ),
    .b(\DFF_858.Q ),
    .y(_04017_)
  );
  al_and3ftt _09628_ (
    .a(_01490_),
    .b(_04017_),
    .c(_01488_),
    .y(_04018_)
  );
  al_and3ftt _09629_ (
    .a(_01078_),
    .b(_04018_),
    .c(_01082_),
    .y(_04019_)
  );
  al_nand3 _09630_ (
    .a(_03525_),
    .b(_04019_),
    .c(_02840_),
    .y(_04020_)
  );
  al_aoi21ftf _09631_ (
    .a(\DFF_155.Q ),
    .b(_00066_),
    .c(_04020_),
    .y(\DFF_95.D )
  );
  al_nand2 _09632_ (
    .a(\DFF_745.Q ),
    .b(\DFF_802.Q ),
    .y(_04021_)
  );
  al_nor2 _09633_ (
    .a(\DFF_745.Q ),
    .b(\DFF_802.Q ),
    .y(_04022_)
  );
  al_and2ft _09634_ (
    .a(_04022_),
    .b(_04021_),
    .y(_04023_)
  );
  al_nand3 _09635_ (
    .a(g35),
    .b(_04023_),
    .c(_00935_),
    .y(_04024_)
  );
  al_ao21ftf _09636_ (
    .a(g35),
    .b(\DFF_802.Q ),
    .c(_04024_),
    .y(\DFF_745.D )
  );
  al_or2 _09637_ (
    .a(_01810_),
    .b(_00721_),
    .y(_04025_)
  );
  al_and2 _09638_ (
    .a(_01809_),
    .b(_00721_),
    .y(_04026_)
  );
  al_nand3 _09639_ (
    .a(_01796_),
    .b(_04026_),
    .c(_01707_),
    .y(_04027_)
  );
  al_aoi21 _09640_ (
    .a(_04025_),
    .b(_04027_),
    .c(_00066_),
    .y(\DFF_1054.D )
  );
  al_mux2l _09641_ (
    .a(\DFF_721.Q ),
    .b(\DFF_276.Q ),
    .s(g35),
    .y(\DFF_721.D )
  );
  al_and2 _09642_ (
    .a(g35),
    .b(\DFF_276.Q ),
    .y(\DFF_276.D )
  );
  al_and3fft _09643_ (
    .a(_01983_),
    .b(_02466_),
    .c(_01984_),
    .y(\DFF_935.D )
  );
  al_nand3ftt _09644_ (
    .a(_02030_),
    .b(_00499_),
    .c(_01070_),
    .y(_04028_)
  );
  al_ao21ftt _09645_ (
    .a(_02030_),
    .b(_01070_),
    .c(\DFF_12.Q ),
    .y(_04029_)
  );
  al_nand3 _09646_ (
    .a(g35),
    .b(_04028_),
    .c(_04029_),
    .y(_04030_)
  );
  al_ao21ftf _09647_ (
    .a(g35),
    .b(\DFF_982.Q ),
    .c(_04030_),
    .y(\DFF_12.D )
  );
  al_nand2 _09648_ (
    .a(\DFF_875.Q ),
    .b(\DFF_1215.Q ),
    .y(_04031_)
  );
  al_nor2 _09649_ (
    .a(\DFF_875.Q ),
    .b(\DFF_1215.Q ),
    .y(_04032_)
  );
  al_nand2ft _09650_ (
    .a(_04032_),
    .b(_04031_),
    .y(_04033_)
  );
  al_mux2l _09651_ (
    .a(\DFF_1079.Q ),
    .b(_04033_),
    .s(_01691_),
    .y(_04034_)
  );
  al_mux2h _09652_ (
    .a(\DFF_1215.Q ),
    .b(_04034_),
    .s(g35),
    .y(\DFF_1079.D )
  );
  al_or2ft _09653_ (
    .a(\DFF_400.Q ),
    .b(_00376_),
    .y(_04035_)
  );
  al_nand2ft _09654_ (
    .a(\DFF_400.Q ),
    .b(_00376_),
    .y(_04036_)
  );
  al_nand3 _09655_ (
    .a(g35),
    .b(_04036_),
    .c(_04035_),
    .y(_04037_)
  );
  al_aoi21ftf _09656_ (
    .a(\DFF_1203.Q ),
    .b(_00066_),
    .c(_04037_),
    .y(\DFF_400.D )
  );
  al_and2ft _09657_ (
    .a(g35),
    .b(\DFF_1347.Q ),
    .y(_04038_)
  );
  al_nand3 _09658_ (
    .a(_00587_),
    .b(_02064_),
    .c(_00389_),
    .y(_04039_)
  );
  al_ao21 _09659_ (
    .a(\DFF_1347.Q ),
    .b(_02064_),
    .c(\DFF_443.Q ),
    .y(_04040_)
  );
  al_nand3 _09660_ (
    .a(\DFF_1347.Q ),
    .b(\DFF_443.Q ),
    .c(_02064_),
    .y(_04041_)
  );
  al_and3 _09661_ (
    .a(g35),
    .b(_04041_),
    .c(_04040_),
    .y(_04042_)
  );
  al_ao21 _09662_ (
    .a(_04042_),
    .b(_04039_),
    .c(_04038_),
    .y(\DFF_443.D )
  );
  al_nor3ftt _09663_ (
    .a(\DFF_644.Q ),
    .b(_00499_),
    .c(_00373_),
    .y(_04043_)
  );
  al_oa21ftt _09664_ (
    .a(\DFF_644.Q ),
    .b(_00373_),
    .c(_00499_),
    .y(_04044_)
  );
  al_nor3ftt _09665_ (
    .a(g35),
    .b(_04043_),
    .c(_04044_),
    .y(\DFF_644.D )
  );
  al_ao21ftf _09666_ (
    .a(g35),
    .b(\DFF_1.Q ),
    .c(_03124_),
    .y(\DFF_865.D )
  );
  al_or3ftt _09667_ (
    .a(g73),
    .b(\DFF_439.Q ),
    .c(g72),
    .y(_04045_)
  );
  al_mux2l _09668_ (
    .a(_04045_),
    .b(\DFF_1022.Q ),
    .s(_01208_),
    .y(\DFF_226.D )
  );
  al_ao21 _09669_ (
    .a(_01690_),
    .b(_01689_),
    .c(_00066_),
    .y(_04046_)
  );
  al_mux2l _09670_ (
    .a(\DFF_875.Q ),
    .b(\DFF_1215.Q ),
    .s(_04046_),
    .y(\DFF_1215.D )
  );
  al_ao21 _09671_ (
    .a(\DFF_506.Q ),
    .b(_01185_),
    .c(\DFF_560.Q ),
    .y(_04047_)
  );
  al_nand3 _09672_ (
    .a(_02276_),
    .b(_01186_),
    .c(_04047_),
    .y(_04048_)
  );
  al_ao21ftf _09673_ (
    .a(g35),
    .b(\DFF_506.Q ),
    .c(_04048_),
    .y(\DFF_560.D )
  );
  al_nand3 _09674_ (
    .a(_00499_),
    .b(_00592_),
    .c(_02862_),
    .y(_04049_)
  );
  al_ao21 _09675_ (
    .a(_00592_),
    .b(_02862_),
    .c(\DFF_192.Q ),
    .y(_04050_)
  );
  al_nand3 _09676_ (
    .a(g35),
    .b(_04050_),
    .c(_04049_),
    .y(_04051_)
  );
  al_ao21ftf _09677_ (
    .a(g35),
    .b(\DFF_398.Q ),
    .c(_04051_),
    .y(\DFF_192.D )
  );
  al_nand2 _09678_ (
    .a(_02339_),
    .b(_02338_),
    .y(_04052_)
  );
  al_or3fft _09679_ (
    .a(\DFF_1278.Q ),
    .b(g35),
    .c(_04052_),
    .y(_04053_)
  );
  al_ao21ttf _09680_ (
    .a(_02339_),
    .b(_02338_),
    .c(_03704_),
    .y(_04054_)
  );
  al_or2 _09681_ (
    .a(\DFF_716.Q ),
    .b(g35),
    .y(_04055_)
  );
  al_and3 _09682_ (
    .a(_04055_),
    .b(_04054_),
    .c(_04053_),
    .y(\DFF_1278.D )
  );
  al_inv _09683_ (
    .a(\DFF_1308.Q ),
    .y(_04056_)
  );
  al_and3fft _09684_ (
    .a(\DFF_600.Q ),
    .b(_02196_),
    .c(_04056_),
    .y(_04057_)
  );
  al_or2ft _09685_ (
    .a(_04057_),
    .b(_03674_),
    .y(_04058_)
  );
  al_nand2ft _09686_ (
    .a(_04057_),
    .b(_03674_),
    .y(_04059_)
  );
  al_nand3 _09687_ (
    .a(g35),
    .b(_04059_),
    .c(_04058_),
    .y(_04060_)
  );
  al_aoi21ftf _09688_ (
    .a(\DFF_606.Q ),
    .b(_00066_),
    .c(_04060_),
    .y(\DFF_675.D )
  );
  al_mux2l _09689_ (
    .a(\DFF_347.Q ),
    .b(\DFF_423.Q ),
    .s(\DFF_286.Q ),
    .y(_04061_)
  );
  al_aoi21 _09690_ (
    .a(\DFF_517.Q ),
    .b(_04061_),
    .c(\DFF_229.Q ),
    .y(_04062_)
  );
  al_oai21 _09691_ (
    .a(\DFF_517.Q ),
    .b(_04061_),
    .c(_04062_),
    .y(_04063_)
  );
  al_ao21ttf _09692_ (
    .a(_03734_),
    .b(_04063_),
    .c(_00585_),
    .y(_04064_)
  );
  al_or2 _09693_ (
    .a(\DFF_229.Q ),
    .b(_00585_),
    .y(_04065_)
  );
  al_and3 _09694_ (
    .a(g35),
    .b(_04064_),
    .c(_04065_),
    .y(\DFF_229.D )
  );
  al_oa21ftt _09695_ (
    .a(\DFF_969.Q ),
    .b(\DFF_1113.Q ),
    .c(g35),
    .y(_04066_)
  );
  al_nand3fft _09696_ (
    .a(\DFF_975.Q ),
    .b(\DFF_969.Q ),
    .c(g35),
    .y(_04067_)
  );
  al_aoi21ttf _09697_ (
    .a(_04067_),
    .b(_04066_),
    .c(\DFF_907.Q ),
    .y(\DFF_3.D )
  );
  al_oai21ttf _09698_ (
    .a(_00575_),
    .b(_00756_),
    .c(_01963_),
    .y(_04068_)
  );
  al_aoi21ftf _09699_ (
    .a(\DFF_962.Q ),
    .b(_00066_),
    .c(_04068_),
    .y(\DFF_893.D )
  );
  al_mux2l _09700_ (
    .a(_00977_),
    .b(\DFF_273.Q ),
    .s(_02045_),
    .y(_04069_)
  );
  al_mux2h _09701_ (
    .a(\DFF_442.Q ),
    .b(_04069_),
    .s(g35),
    .y(\DFF_273.D )
  );
  al_and2ft _09702_ (
    .a(g35),
    .b(\DFF_381.Q ),
    .y(_04070_)
  );
  al_aoi21ftt _09703_ (
    .a(_01639_),
    .b(_01635_),
    .c(_03294_),
    .y(_04071_)
  );
  al_ao21ftf _09704_ (
    .a(_01638_),
    .b(_01634_),
    .c(_04071_),
    .y(_04072_)
  );
  al_ao21ftf _09705_ (
    .a(_01633_),
    .b(_01641_),
    .c(_04072_),
    .y(_04073_)
  );
  al_oa21ftf _09706_ (
    .a(\DFF_1334.Q ),
    .b(_04072_),
    .c(_00066_),
    .y(_04074_)
  );
  al_ao21 _09707_ (
    .a(_04073_),
    .b(_04074_),
    .c(_04070_),
    .y(\DFF_1334.D )
  );
  al_mux2l _09708_ (
    .a(\DFF_1313.Q ),
    .b(_00522_),
    .s(_02421_),
    .y(_04075_)
  );
  al_mux2h _09709_ (
    .a(\DFF_375.Q ),
    .b(_04075_),
    .s(g35),
    .y(\DFF_1313.D )
  );
  al_or2ft _09710_ (
    .a(\DFF_4.Q ),
    .b(_01914_),
    .y(_04076_)
  );
  al_ao21ftf _09711_ (
    .a(_00530_),
    .b(_01914_),
    .c(_04076_),
    .y(_04077_)
  );
  al_mux2h _09712_ (
    .a(\DFF_637.Q ),
    .b(_04077_),
    .s(g35),
    .y(\DFF_4.D )
  );
  al_nand3 _09713_ (
    .a(_00499_),
    .b(_02426_),
    .c(_02707_),
    .y(_04078_)
  );
  al_ao21 _09714_ (
    .a(_02426_),
    .b(_02707_),
    .c(\DFF_986.Q ),
    .y(_04079_)
  );
  al_nand3 _09715_ (
    .a(g35),
    .b(_04079_),
    .c(_04078_),
    .y(_04080_)
  );
  al_ao21ftf _09716_ (
    .a(g35),
    .b(\DFF_312.Q ),
    .c(_04080_),
    .y(\DFF_986.D )
  );
  al_ao21 _09717_ (
    .a(\DFF_20.Q ),
    .b(\DFF_104.Q ),
    .c(\DFF_916.Q ),
    .y(_04081_)
  );
  al_nand3ftt _09718_ (
    .a(_02170_),
    .b(_04081_),
    .c(_02804_),
    .y(_04082_)
  );
  al_ao21ftf _09719_ (
    .a(g35),
    .b(\DFF_20.Q ),
    .c(_04082_),
    .y(\DFF_916.D )
  );
  al_ao21ftf _09720_ (
    .a(g113),
    .b(_00342_),
    .c(\DFF_946.Q ),
    .y(_04083_)
  );
  al_aoi21ttf _09721_ (
    .a(\DFF_1111.Q ),
    .b(_00604_),
    .c(_04083_),
    .y(_04084_)
  );
  al_mux2h _09722_ (
    .a(\DFF_319.Q ),
    .b(_04084_),
    .s(_03269_),
    .y(_04085_)
  );
  al_mux2h _09723_ (
    .a(\DFF_931.Q ),
    .b(_04085_),
    .s(g35),
    .y(\DFF_319.D )
  );
  al_and2ft _09724_ (
    .a(g35),
    .b(\DFF_592.Q ),
    .y(_04086_)
  );
  al_and2 _09725_ (
    .a(_02133_),
    .b(_02135_),
    .y(_04087_)
  );
  al_ao21 _09726_ (
    .a(_04087_),
    .b(_01948_),
    .c(_02131_),
    .y(_04088_)
  );
  al_nand3 _09727_ (
    .a(_02131_),
    .b(_02133_),
    .c(_02135_),
    .y(_04089_)
  );
  al_and2 _09728_ (
    .a(g35),
    .b(_04089_),
    .y(_04090_)
  );
  al_ao21 _09729_ (
    .a(_04090_),
    .b(_04088_),
    .c(_04086_),
    .y(\DFF_521.D )
  );
  al_mux2l _09730_ (
    .a(\DFF_881.Q ),
    .b(\DFF_1035.Q ),
    .s(g35),
    .y(\DFF_881.D )
  );
  al_oai21ttf _09731_ (
    .a(\DFF_375.Q ),
    .b(_03125_),
    .c(_02422_),
    .y(_04091_)
  );
  al_ao21ftf _09732_ (
    .a(g35),
    .b(\DFF_1371.Q ),
    .c(_04091_),
    .y(\DFF_375.D )
  );
  al_oai21ftt _09733_ (
    .a(\DFF_1044.Q ),
    .b(\DFF_770.Q ),
    .c(g35),
    .y(_04092_)
  );
  al_ao21ftf _09734_ (
    .a(g35),
    .b(\DFF_1391.Q ),
    .c(_04092_),
    .y(\DFF_770.D )
  );
  al_ao21 _09735_ (
    .a(\DFF_1107.Q ),
    .b(_00466_),
    .c(\DFF_218.Q ),
    .y(_04093_)
  );
  al_nand3ftt _09736_ (
    .a(_01989_),
    .b(_04093_),
    .c(_01984_),
    .y(_04094_)
  );
  al_ao21ftf _09737_ (
    .a(g35),
    .b(\DFF_1176.Q ),
    .c(_04094_),
    .y(\DFF_218.D )
  );
  al_nand3 _09738_ (
    .a(_00499_),
    .b(_02029_),
    .c(_01046_),
    .y(_04095_)
  );
  al_ao21 _09739_ (
    .a(_02029_),
    .b(_01046_),
    .c(\DFF_1177.Q ),
    .y(_04096_)
  );
  al_nand3 _09740_ (
    .a(g35),
    .b(_04095_),
    .c(_04096_),
    .y(_04097_)
  );
  al_ao21ftf _09741_ (
    .a(g35),
    .b(\DFF_1244.Q ),
    .c(_04097_),
    .y(\DFF_1177.D )
  );
  al_nand3 _09742_ (
    .a(_00499_),
    .b(_01702_),
    .c(_01745_),
    .y(_04098_)
  );
  al_ao21 _09743_ (
    .a(_01745_),
    .b(_01702_),
    .c(\DFF_884.Q ),
    .y(_04099_)
  );
  al_nand3 _09744_ (
    .a(g35),
    .b(_04099_),
    .c(_04098_),
    .y(_04100_)
  );
  al_ao21ftf _09745_ (
    .a(g35),
    .b(\DFF_51.Q ),
    .c(_04100_),
    .y(\DFF_884.D )
  );
  al_ao21ttf _09746_ (
    .a(_02090_),
    .b(_02064_),
    .c(\DFF_1302.Q ),
    .y(_04101_)
  );
  al_nand2ft _09747_ (
    .a(\DFF_1342.Q ),
    .b(g35),
    .y(_04102_)
  );
  al_ao21ftf _09748_ (
    .a(_04102_),
    .b(\DFF_1358.Q ),
    .c(_03855_),
    .y(_04103_)
  );
  al_and3ftt _09749_ (
    .a(\DFF_1358.Q ),
    .b(_04102_),
    .c(_03855_),
    .y(_04104_)
  );
  al_aoi21 _09750_ (
    .a(_04101_),
    .b(_04103_),
    .c(_04104_),
    .y(\DFF_1302.D )
  );
  al_nand3 _09751_ (
    .a(_00499_),
    .b(_01312_),
    .c(_01976_),
    .y(_04105_)
  );
  al_ao21 _09752_ (
    .a(_01312_),
    .b(_01976_),
    .c(\DFF_1186.Q ),
    .y(_04106_)
  );
  al_nand3 _09753_ (
    .a(g35),
    .b(_04106_),
    .c(_04105_),
    .y(_04107_)
  );
  al_ao21ftf _09754_ (
    .a(g35),
    .b(\DFF_1325.Q ),
    .c(_04107_),
    .y(\DFF_1186.D )
  );
  al_ao21 _09755_ (
    .a(\DFF_99.Q ),
    .b(\DFF_1326.Q ),
    .c(\DFF_1029.Q ),
    .y(_04108_)
  );
  al_nand3ftt _09756_ (
    .a(_00466_),
    .b(_04108_),
    .c(_01984_),
    .y(_04109_)
  );
  al_ao21ftf _09757_ (
    .a(g35),
    .b(\DFF_1326.Q ),
    .c(_04109_),
    .y(\DFF_1029.D )
  );
  al_nand2 _09758_ (
    .a(\DFF_936.Q ),
    .b(_01481_),
    .y(_04110_)
  );
  al_or2 _09759_ (
    .a(\DFF_936.Q ),
    .b(_01481_),
    .y(_04111_)
  );
  al_nand3 _09760_ (
    .a(_04110_),
    .b(_04111_),
    .c(_03462_),
    .y(_04112_)
  );
  al_ao21ftf _09761_ (
    .a(g35),
    .b(\DFF_1237.Q ),
    .c(_04112_),
    .y(\DFF_936.D )
  );
  al_and2 _09762_ (
    .a(\DFF_130.Q ),
    .b(_02146_),
    .y(\DFF_160.D )
  );
  al_and2ft _09763_ (
    .a(\DFF_685.Q ),
    .b(g35),
    .y(_04113_)
  );
  al_nand3fft _09764_ (
    .a(\DFF_155.Q ),
    .b(\DFF_116.Q ),
    .c(_04113_),
    .y(_04114_)
  );
  al_aoi21ftf _09765_ (
    .a(g35),
    .b(_00270_),
    .c(_04114_),
    .y(\DFF_155.D )
  );
  al_or3 _09766_ (
    .a(\DFF_350.Q ),
    .b(g73),
    .c(g72),
    .y(_04115_)
  );
  al_mux2l _09767_ (
    .a(_04115_),
    .b(\DFF_1349.Q ),
    .s(_01208_),
    .y(\DFF_1362.D )
  );
  al_nor2 _09768_ (
    .a(\DFF_1015.Q ),
    .b(g35),
    .y(_04116_)
  );
  al_or2 _09769_ (
    .a(\DFF_1015.Q ),
    .b(_01999_),
    .y(_04117_)
  );
  al_aoi21ftf _09770_ (
    .a(_01997_),
    .b(_01995_),
    .c(_04117_),
    .y(_04118_)
  );
  al_nand3 _09771_ (
    .a(\DFF_260.Q ),
    .b(_02004_),
    .c(_04118_),
    .y(_04119_)
  );
  al_oa21ttf _09772_ (
    .a(\DFF_260.Q ),
    .b(_04118_),
    .c(_00066_),
    .y(_04120_)
  );
  al_aoi21 _09773_ (
    .a(_04119_),
    .b(_04120_),
    .c(_04116_),
    .y(\DFF_260.D )
  );
  al_mux2l _09774_ (
    .a(\DFF_900.Q ),
    .b(\DFF_866.Q ),
    .s(_01349_),
    .y(\DFF_866.D )
  );
  al_nand3 _09775_ (
    .a(_00499_),
    .b(_00591_),
    .c(_01467_),
    .y(_04121_)
  );
  al_ao21 _09776_ (
    .a(_00591_),
    .b(_01467_),
    .c(\DFF_336.Q ),
    .y(_04122_)
  );
  al_nand3 _09777_ (
    .a(g35),
    .b(_04121_),
    .c(_04122_),
    .y(_04123_)
  );
  al_ao21ftf _09778_ (
    .a(g35),
    .b(\DFF_949.Q ),
    .c(_04123_),
    .y(\DFF_336.D )
  );
  al_mux2l _09779_ (
    .a(\DFF_1018.Q ),
    .b(\DFF_388.Q ),
    .s(_01353_),
    .y(\DFF_388.D )
  );
  al_and3ftt _09780_ (
    .a(\DFF_871.Q ),
    .b(\DFF_1275.Q ),
    .c(g35),
    .y(\DFF_871.D )
  );
  al_mux2h _09781_ (
    .a(\DFF_466.Q ),
    .b(_02004_),
    .s(g35),
    .y(\DFF_1333.D )
  );
  al_mux2h _09782_ (
    .a(\DFF_1257.Q ),
    .b(_01041_),
    .s(g35),
    .y(\DFF_1113.D )
  );
  al_oa21ftt _09783_ (
    .a(g35),
    .b(\DFF_879.Q ),
    .c(\DFF_821.Q ),
    .y(\DFF_596.D )
  );
  al_mux2l _09784_ (
    .a(\DFF_1115.Q ),
    .b(\DFF_442.Q ),
    .s(_02190_),
    .y(\DFF_442.D )
  );
  al_and2ft _09785_ (
    .a(g35),
    .b(\DFF_833.Q ),
    .y(_04124_)
  );
  al_nand3 _09786_ (
    .a(_00587_),
    .b(_01956_),
    .c(_00398_),
    .y(_04125_)
  );
  al_ao21 _09787_ (
    .a(\DFF_833.Q ),
    .b(_01956_),
    .c(\DFF_429.Q ),
    .y(_04126_)
  );
  al_nand2 _09788_ (
    .a(_00399_),
    .b(_01956_),
    .y(_04127_)
  );
  al_and3 _09789_ (
    .a(g35),
    .b(_04127_),
    .c(_04126_),
    .y(_04128_)
  );
  al_ao21 _09790_ (
    .a(_04128_),
    .b(_04125_),
    .c(_04124_),
    .y(\DFF_429.D )
  );
  al_aoi21 _09791_ (
    .a(\DFF_724.Q ),
    .b(g35),
    .c(\DFF_268.Q ),
    .y(_04129_)
  );
  al_ao21ftf _09792_ (
    .a(_04129_),
    .b(_03453_),
    .c(_03452_),
    .y(\DFF_352.D )
  );
  al_nand2 _09793_ (
    .a(\DFF_1369.Q ),
    .b(\DFF_1184.Q ),
    .y(_04130_)
  );
  al_nor2 _09794_ (
    .a(\DFF_1369.Q ),
    .b(\DFF_1184.Q ),
    .y(_04131_)
  );
  al_nand2ft _09795_ (
    .a(_04131_),
    .b(_04130_),
    .y(_04132_)
  );
  al_mux2l _09796_ (
    .a(\DFF_520.Q ),
    .b(_04132_),
    .s(_02776_),
    .y(_04133_)
  );
  al_mux2h _09797_ (
    .a(\DFF_1369.Q ),
    .b(_04133_),
    .s(g35),
    .y(\DFF_520.D )
  );
  al_or2ft _09798_ (
    .a(g35),
    .b(_02278_),
    .y(_04134_)
  );
  al_mux2l _09799_ (
    .a(\DFF_167.Q ),
    .b(\DFF_182.Q ),
    .s(_04134_),
    .y(\DFF_182.D )
  );
  al_ao21ftf _09800_ (
    .a(_01622_),
    .b(_00767_),
    .c(_03879_),
    .y(_04135_)
  );
  al_ao21ftf _09801_ (
    .a(g35),
    .b(\DFF_290.Q ),
    .c(_04135_),
    .y(\DFF_664.D )
  );
  al_nand3ftt _09802_ (
    .a(_01768_),
    .b(_00499_),
    .c(_02930_),
    .y(_04136_)
  );
  al_ao21ftt _09803_ (
    .a(_01768_),
    .b(_02930_),
    .c(\DFF_579.Q ),
    .y(_04137_)
  );
  al_nand3 _09804_ (
    .a(g35),
    .b(_04136_),
    .c(_04137_),
    .y(_04138_)
  );
  al_ao21ftf _09805_ (
    .a(g35),
    .b(\DFF_916.Q ),
    .c(_04138_),
    .y(\DFF_579.D )
  );
  al_or3ftt _09806_ (
    .a(_01125_),
    .b(_00327_),
    .c(_01131_),
    .y(_04139_)
  );
  al_ao21ftt _09807_ (
    .a(_00327_),
    .b(_01125_),
    .c(\DFF_504.Q ),
    .y(_04140_)
  );
  al_nand3 _09808_ (
    .a(g35),
    .b(_04140_),
    .c(_04139_),
    .y(_04141_)
  );
  al_ao21ftf _09809_ (
    .a(g35),
    .b(\DFF_1422.Q ),
    .c(_04141_),
    .y(\DFF_504.D )
  );
  al_mux2l _09810_ (
    .a(\DFF_1195.Q ),
    .b(\DFF_87.Q ),
    .s(_02694_),
    .y(\DFF_87.D )
  );
  al_oai21ftt _09811_ (
    .a(g35),
    .b(_00758_),
    .c(\DFF_1082.Q ),
    .y(_04142_)
  );
  al_nand3 _09812_ (
    .a(\DFF_568.Q ),
    .b(g35),
    .c(_03552_),
    .y(_04143_)
  );
  al_and2ft _09813_ (
    .a(_04142_),
    .b(_04143_),
    .y(_04144_)
  );
  al_or2ft _09814_ (
    .a(_04142_),
    .b(_04143_),
    .y(_04145_)
  );
  al_nand2ft _09815_ (
    .a(_04144_),
    .b(_04145_),
    .y(\DFF_568.D )
  );
  al_ao21 _09816_ (
    .a(g35),
    .b(\DFF_87.Q ),
    .c(\DFF_546.Q ),
    .y(_04146_)
  );
  al_aoi21 _09817_ (
    .a(g35),
    .b(_00984_),
    .c(_04146_),
    .y(_04147_)
  );
  al_ao21ttf _09818_ (
    .a(_00983_),
    .b(_00585_),
    .c(\DFF_742.Q ),
    .y(_04148_)
  );
  al_nand2 _09819_ (
    .a(\DFF_546.Q ),
    .b(\DFF_87.Q ),
    .y(_04149_)
  );
  al_oa21ftf _09820_ (
    .a(_04149_),
    .b(_00984_),
    .c(_00066_),
    .y(_04150_)
  );
  al_aoi21 _09821_ (
    .a(_04148_),
    .b(_04150_),
    .c(_04147_),
    .y(\DFF_742.D )
  );
  al_oai21ttf _09822_ (
    .a(\DFF_1375.Q ),
    .b(_02360_),
    .c(_00066_),
    .y(_04151_)
  );
  al_or3fft _09823_ (
    .a(_00541_),
    .b(g35),
    .c(_00546_),
    .y(_04152_)
  );
  al_aoi21ftf _09824_ (
    .a(\DFF_984.Q ),
    .b(_00066_),
    .c(_04152_),
    .y(_04153_)
  );
  al_aoi21ftf _09825_ (
    .a(_04151_),
    .b(_01544_),
    .c(_04153_),
    .y(\DFF_552.D )
  );
  al_nand3 _09826_ (
    .a(_00499_),
    .b(_01408_),
    .c(_00567_),
    .y(_04154_)
  );
  al_ao21 _09827_ (
    .a(_01408_),
    .b(_00567_),
    .c(\DFF_497.Q ),
    .y(_04155_)
  );
  al_nand3 _09828_ (
    .a(g35),
    .b(_04154_),
    .c(_04155_),
    .y(_04156_)
  );
  al_ao21ftf _09829_ (
    .a(g35),
    .b(\DFF_1095.Q ),
    .c(_04156_),
    .y(\DFF_497.D )
  );
  al_nand2ft _09830_ (
    .a(\DFF_395.Q ),
    .b(_00519_),
    .y(_04157_)
  );
  al_aoi21ttf _09831_ (
    .a(_04157_),
    .b(_00529_),
    .c(_00526_),
    .y(_04158_)
  );
  al_or3fft _09832_ (
    .a(\DFF_795.Q ),
    .b(_04158_),
    .c(_01914_),
    .y(_04159_)
  );
  al_oai21ftf _09833_ (
    .a(\DFF_795.Q ),
    .b(_01914_),
    .c(_04158_),
    .y(_04160_)
  );
  al_ao21 _09834_ (
    .a(_04159_),
    .b(_04160_),
    .c(_00066_),
    .y(_04161_)
  );
  al_aoi21ftf _09835_ (
    .a(\DFF_1233.Q ),
    .b(_00066_),
    .c(_04161_),
    .y(\DFF_795.D )
  );
  al_oai21 _09836_ (
    .a(\DFF_758.Q ),
    .b(\DFF_127.Q ),
    .c(g35),
    .y(_04162_)
  );
  al_ao21ftf _09837_ (
    .a(g35),
    .b(\DFF_453.Q ),
    .c(_04162_),
    .y(\DFF_127.D )
  );
  al_nand3ftt _09838_ (
    .a(_02368_),
    .b(_00499_),
    .c(_00597_),
    .y(_04163_)
  );
  al_ao21ftt _09839_ (
    .a(_02368_),
    .b(_00597_),
    .c(\DFF_1350.Q ),
    .y(_04164_)
  );
  al_nand3 _09840_ (
    .a(g35),
    .b(_04163_),
    .c(_04164_),
    .y(_04165_)
  );
  al_ao21ftf _09841_ (
    .a(g35),
    .b(\DFF_590.Q ),
    .c(_04165_),
    .y(\DFF_1350.D )
  );
  al_ao21 _09842_ (
    .a(g35),
    .b(\DFF_482.Q ),
    .c(\DFF_490.Q ),
    .y(_04166_)
  );
  al_and3 _09843_ (
    .a(g35),
    .b(\DFF_482.Q ),
    .c(\DFF_490.Q ),
    .y(_04167_)
  );
  al_aoi21ttf _09844_ (
    .a(\DFF_1146.Q ),
    .b(\DFF_692.Q ),
    .c(g35),
    .y(_04168_)
  );
  al_oai21 _09845_ (
    .a(\DFF_1146.Q ),
    .b(\DFF_692.Q ),
    .c(_04168_),
    .y(_04169_)
  );
  al_ao21ftf _09846_ (
    .a(_04167_),
    .b(_04166_),
    .c(_04169_),
    .y(\DFF_1221.D )
  );
  al_ao21 _09847_ (
    .a(_01957_),
    .b(_01956_),
    .c(_00066_),
    .y(_04170_)
  );
  al_mux2l _09848_ (
    .a(\DFF_1306.Q ),
    .b(\DFF_632.Q ),
    .s(_04170_),
    .y(\DFF_632.D )
  );
  al_or3fft _09849_ (
    .a(\DFF_955.Q ),
    .b(g35),
    .c(_00809_),
    .y(_04171_)
  );
  al_ao21ttf _09850_ (
    .a(_00793_),
    .b(_00766_),
    .c(_01802_),
    .y(_04172_)
  );
  al_or2 _09851_ (
    .a(\DFF_778.Q ),
    .b(g35),
    .y(_04173_)
  );
  al_and3 _09852_ (
    .a(_04173_),
    .b(_04172_),
    .c(_04171_),
    .y(\DFF_955.D )
  );
  al_nor2 _09853_ (
    .a(\DFF_216.Q ),
    .b(\DFF_571.Q ),
    .y(_04174_)
  );
  al_nand2 _09854_ (
    .a(\DFF_216.Q ),
    .b(\DFF_571.Q ),
    .y(_04175_)
  );
  al_nand2ft _09855_ (
    .a(_04174_),
    .b(_04175_),
    .y(_04176_)
  );
  al_mux2l _09856_ (
    .a(_04176_),
    .b(\DFF_444.Q ),
    .s(_01914_),
    .y(_04177_)
  );
  al_mux2h _09857_ (
    .a(\DFF_216.Q ),
    .b(_04177_),
    .s(g35),
    .y(\DFF_444.D )
  );
  al_ao21 _09858_ (
    .a(\DFF_1189.Q ),
    .b(_00966_),
    .c(\DFF_614.Q ),
    .y(_04178_)
  );
  al_nand3 _09859_ (
    .a(_00967_),
    .b(_04178_),
    .c(_02741_),
    .y(_04179_)
  );
  al_ao21ftf _09860_ (
    .a(g35),
    .b(\DFF_1189.Q ),
    .c(_04179_),
    .y(\DFF_614.D )
  );
  al_mux2l _09861_ (
    .a(\DFF_571.Q ),
    .b(\DFF_216.Q ),
    .s(_02561_),
    .y(\DFF_216.D )
  );
  al_and2 _09862_ (
    .a(\DFF_965.Q ),
    .b(\DFF_549.Q ),
    .y(_04180_)
  );
  al_aoi21 _09863_ (
    .a(_04180_),
    .b(_01824_),
    .c(_00066_),
    .y(\DFF_440.D )
  );
  al_nand3 _09864_ (
    .a(\DFF_896.Q ),
    .b(g35),
    .c(_00941_),
    .y(_04181_)
  );
  al_aoi21 _09865_ (
    .a(\DFF_789.Q ),
    .b(_00952_),
    .c(_04181_),
    .y(_04182_)
  );
  al_ao21ftt _09866_ (
    .a(g35),
    .b(\DFF_789.Q ),
    .c(_00193_),
    .y(_04183_)
  );
  al_ao21 _09867_ (
    .a(_04183_),
    .b(_02375_),
    .c(_04182_),
    .y(\DFF_896.D )
  );
  al_nand2 _09868_ (
    .a(g35),
    .b(_02019_),
    .y(_04184_)
  );
  al_mux2l _09869_ (
    .a(\DFF_33.Q ),
    .b(\DFF_1226.Q ),
    .s(_04184_),
    .y(\DFF_1226.D )
  );
  al_nand2 _09870_ (
    .a(_02820_),
    .b(_00576_),
    .y(_04185_)
  );
  al_nand2 _09871_ (
    .a(\DFF_835.Q ),
    .b(\DFF_558.Q ),
    .y(_04186_)
  );
  al_nor2 _09872_ (
    .a(\DFF_835.Q ),
    .b(\DFF_558.Q ),
    .y(_04187_)
  );
  al_nand2ft _09873_ (
    .a(_04187_),
    .b(_04186_),
    .y(_04188_)
  );
  al_mux2l _09874_ (
    .a(\DFF_1031.Q ),
    .b(_04188_),
    .s(_04185_),
    .y(_04189_)
  );
  al_mux2h _09875_ (
    .a(\DFF_558.Q ),
    .b(_04189_),
    .s(g35),
    .y(\DFF_1031.D )
  );
  al_oa21ftt _09876_ (
    .a(g35),
    .b(\DFF_636.Q ),
    .c(\DFF_438.Q ),
    .y(_04190_)
  );
  al_aoi21ftf _09877_ (
    .a(\DFF_869.Q ),
    .b(g35),
    .c(_04190_),
    .y(_04191_)
  );
  al_or3fft _09878_ (
    .a(\DFF_459.Q ),
    .b(g35),
    .c(_04191_),
    .y(_04192_)
  );
  al_aoi21ftf _09879_ (
    .a(_00066_),
    .b(\DFF_459.Q ),
    .c(_04191_),
    .y(_04193_)
  );
  al_nand2ft _09880_ (
    .a(_04193_),
    .b(_04192_),
    .y(\DFF_459.D )
  );
  al_and2ft _09881_ (
    .a(g35),
    .b(\DFF_1060.Q ),
    .y(_04194_)
  );
  al_aoi21ftf _09882_ (
    .a(\DFF_1339.Q ),
    .b(_00489_),
    .c(_00495_),
    .y(_04195_)
  );
  al_ao21 _09883_ (
    .a(_00490_),
    .b(_04195_),
    .c(_04194_),
    .y(\DFF_1339.D )
  );
  al_nand3 _09884_ (
    .a(_01358_),
    .b(_02682_),
    .c(_01359_),
    .y(_04196_)
  );
  al_ao21ftf _09885_ (
    .a(g35),
    .b(\DFF_803.Q ),
    .c(_04196_),
    .y(\DFF_54.D )
  );
  al_mux2l _09886_ (
    .a(\DFF_1126.Q ),
    .b(\DFF_656.Q ),
    .s(_01054_),
    .y(\DFF_656.D )
  );
  al_mux2h _09887_ (
    .a(\DFF_1415.Q ),
    .b(_03440_),
    .s(g35),
    .y(\DFF_1345.D )
  );
  al_nand3 _09888_ (
    .a(_00499_),
    .b(_01114_),
    .c(_01467_),
    .y(_04197_)
  );
  al_ao21 _09889_ (
    .a(_01114_),
    .b(_01467_),
    .c(\DFF_471.Q ),
    .y(_04198_)
  );
  al_nand3 _09890_ (
    .a(g35),
    .b(_04198_),
    .c(_04197_),
    .y(_04199_)
  );
  al_ao21ftf _09891_ (
    .a(g35),
    .b(\DFF_1085.Q ),
    .c(_04199_),
    .y(\DFF_471.D )
  );
  al_and3ftt _09892_ (
    .a(\DFF_894.Q ),
    .b(\DFF_849.Q ),
    .c(_00461_),
    .y(_04200_)
  );
  al_or2 _09893_ (
    .a(\DFF_1006.Q ),
    .b(_04200_),
    .y(_04201_)
  );
  al_ao21ttf _09894_ (
    .a(_01221_),
    .b(_04201_),
    .c(_01226_),
    .y(_04202_)
  );
  al_ao21 _09895_ (
    .a(_04200_),
    .b(_01222_),
    .c(_00066_),
    .y(_04203_)
  );
  al_aoi21ftf _09896_ (
    .a(\DFF_837.Q ),
    .b(_04203_),
    .c(_04202_),
    .y(\DFF_1006.D )
  );
  al_nand3 _09897_ (
    .a(\DFF_119.Q ),
    .b(\DFF_751.Q ),
    .c(_01562_),
    .y(_04204_)
  );
  al_nand2ft _09898_ (
    .a(\DFF_119.Q ),
    .b(_01237_),
    .y(_04205_)
  );
  al_nand3 _09899_ (
    .a(_02276_),
    .b(_04205_),
    .c(_04204_),
    .y(_04206_)
  );
  al_ao21ftf _09900_ (
    .a(g35),
    .b(\DFF_751.Q ),
    .c(_04206_),
    .y(\DFF_119.D )
  );
  al_oai21ftf _09901_ (
    .a(\DFF_545.Q ),
    .b(\DFF_1228.Q ),
    .c(\DFF_366.Q ),
    .y(_04207_)
  );
  al_nand3ftt _09902_ (
    .a(\DFF_678.Q ),
    .b(g35),
    .c(_04207_),
    .y(_04208_)
  );
  al_ao21ftf _09903_ (
    .a(g35),
    .b(\DFF_1228.Q ),
    .c(_04208_),
    .y(\DFF_366.D )
  );
  al_oai21ttf _09904_ (
    .a(\DFF_1057.Q ),
    .b(_02870_),
    .c(_03245_),
    .y(_04209_)
  );
  al_ao21ftf _09905_ (
    .a(g35),
    .b(\DFF_90.Q ),
    .c(_04209_),
    .y(\DFF_1057.D )
  );
  al_nor2 _09906_ (
    .a(g35),
    .b(\DFF_1423.Q ),
    .y(_04210_)
  );
  al_oa21ftf _09907_ (
    .a(\DFF_1205.Q ),
    .b(_01689_),
    .c(_00066_),
    .y(_04211_)
  );
  al_aoi21 _09908_ (
    .a(_04211_),
    .b(_02528_),
    .c(_04210_),
    .y(\DFF_1205.D )
  );
  al_nand3 _09909_ (
    .a(_02192_),
    .b(_01702_),
    .c(_01894_),
    .y(_04212_)
  );
  al_ao21ftf _09910_ (
    .a(g35),
    .b(\DFF_958.Q ),
    .c(_04212_),
    .y(\DFF_289.D )
  );
  al_and2ft _09911_ (
    .a(g35),
    .b(\DFF_386.Q ),
    .y(_04213_)
  );
  al_nor2ft _09912_ (
    .a(_01087_),
    .b(_01090_),
    .y(_04214_)
  );
  al_ao21 _09913_ (
    .a(_04214_),
    .b(_01101_),
    .c(_01085_),
    .y(_04215_)
  );
  al_oa21ttf _09914_ (
    .a(_01090_),
    .b(_03868_),
    .c(_00066_),
    .y(_04216_)
  );
  al_ao21 _09915_ (
    .a(_04216_),
    .b(_04215_),
    .c(_04213_),
    .y(\DFF_690.D )
  );
  al_mux2l _09916_ (
    .a(\DFF_292.Q ),
    .b(\DFF_533.Q ),
    .s(_01109_),
    .y(\DFF_533.D )
  );
  al_and2ft _09917_ (
    .a(\DFF_1144.Q ),
    .b(\DFF_979.Q ),
    .y(_04217_)
  );
  al_mux2l _09918_ (
    .a(_04217_),
    .b(\DFF_1144.Q ),
    .s(_03659_),
    .y(_04218_)
  );
  al_mux2h _09919_ (
    .a(\DFF_486.Q ),
    .b(_04218_),
    .s(g35),
    .y(\DFF_1144.D )
  );
  al_nand2 _09920_ (
    .a(\DFF_452.Q ),
    .b(\DFF_417.D ),
    .y(_04219_)
  );
  al_oa21ttf _09921_ (
    .a(\DFF_894.Q ),
    .b(\DFF_849.Q ),
    .c(_01661_),
    .y(_04220_)
  );
  al_ao21ftf _09922_ (
    .a(_01224_),
    .b(\DFF_177.Q ),
    .c(_04220_),
    .y(_04221_)
  );
  al_ao21 _09923_ (
    .a(_04221_),
    .b(_04219_),
    .c(\DFF_62.Q ),
    .y(_04222_)
  );
  al_and3ftt _09924_ (
    .a(\DFF_894.Q ),
    .b(\DFF_849.Q ),
    .c(\DFF_677.Q ),
    .y(_04223_)
  );
  al_aoi21 _09925_ (
    .a(\DFF_1193.Q ),
    .b(_00455_),
    .c(_04223_),
    .y(_04224_)
  );
  al_nand3fft _09926_ (
    .a(\DFF_894.Q ),
    .b(\DFF_849.Q ),
    .c(\DFF_161.Q ),
    .y(_04225_)
  );
  al_nand3 _09927_ (
    .a(\DFF_894.Q ),
    .b(\DFF_849.Q ),
    .c(\DFF_1157.Q ),
    .y(_04226_)
  );
  al_and3 _09928_ (
    .a(_04225_),
    .b(_04226_),
    .c(_04224_),
    .y(_04227_)
  );
  al_nand2ft _09929_ (
    .a(\DFF_417.D ),
    .b(_04227_),
    .y(_04228_)
  );
  al_nand2ft _09930_ (
    .a(_04227_),
    .b(\DFF_417.D ),
    .y(_04229_)
  );
  al_nand3 _09931_ (
    .a(_00007_),
    .b(_04228_),
    .c(_04229_),
    .y(_04230_)
  );
  al_and3fft _09932_ (
    .a(_01730_),
    .b(_00461_),
    .c(_01660_),
    .y(_04231_)
  );
  al_nand3 _09933_ (
    .a(_04231_),
    .b(_04222_),
    .c(_04230_),
    .y(_04232_)
  );
  al_or2 _09934_ (
    .a(\DFF_635.Q ),
    .b(_01730_),
    .y(_04233_)
  );
  al_nand2 _09935_ (
    .a(\DFF_792.Q ),
    .b(\DFF_132.Q ),
    .y(_04234_)
  );
  al_aoi21ttf _09936_ (
    .a(\DFF_699.Q ),
    .b(\DFF_249.Q ),
    .c(_04234_),
    .y(_04235_)
  );
  al_nand2ft _09937_ (
    .a(\DFF_493.Q ),
    .b(\DFF_635.Q ),
    .y(_04236_)
  );
  al_ao21ftf _09938_ (
    .a(\DFF_1205.Q ),
    .b(\DFF_107.Q ),
    .c(_04236_),
    .y(_04237_)
  );
  al_nand3ftt _09939_ (
    .a(_04237_),
    .b(_04233_),
    .c(_04235_),
    .y(_04238_)
  );
  al_and3 _09940_ (
    .a(g35),
    .b(_04238_),
    .c(_04232_),
    .y(\DFF_1425.D )
  );
  al_nand3 _09941_ (
    .a(_00499_),
    .b(_02029_),
    .c(_02010_),
    .y(_04239_)
  );
  al_ao21 _09942_ (
    .a(_02010_),
    .b(_02029_),
    .c(\DFF_628.Q ),
    .y(_04240_)
  );
  al_nand3 _09943_ (
    .a(g35),
    .b(_04240_),
    .c(_04239_),
    .y(_04241_)
  );
  al_ao21ftf _09944_ (
    .a(g35),
    .b(\DFF_309.Q ),
    .c(_04241_),
    .y(\DFF_628.D )
  );
  al_or3ftt _09945_ (
    .a(g73),
    .b(\DFF_221.Q ),
    .c(g72),
    .y(_04242_)
  );
  al_mux2l _09946_ (
    .a(_04242_),
    .b(\DFF_624.Q ),
    .s(_01208_),
    .y(\DFF_268.D )
  );
  al_or2 _09947_ (
    .a(_01646_),
    .b(_01125_),
    .y(_04243_)
  );
  al_and2 _09948_ (
    .a(_01128_),
    .b(_01125_),
    .y(_04244_)
  );
  al_nand3 _09949_ (
    .a(_04244_),
    .b(_02686_),
    .c(_01531_),
    .y(_04245_)
  );
  al_aoi21 _09950_ (
    .a(_04243_),
    .b(_04245_),
    .c(_00066_),
    .y(\DFF_111.D )
  );
  al_and2 _09951_ (
    .a(\DFF_198.Q ),
    .b(g35),
    .y(_04246_)
  );
  al_aoi21ttf _09952_ (
    .a(_04246_),
    .b(_03028_),
    .c(\DFF_1130.Q ),
    .y(\DFF_683.D )
  );
  al_mux2l _09953_ (
    .a(\DFF_362.Q ),
    .b(\DFF_404.Q ),
    .s(_01557_),
    .y(_04247_)
  );
  al_mux2h _09954_ (
    .a(\DFF_648.Q ),
    .b(_04247_),
    .s(g35),
    .y(\DFF_362.D )
  );
  al_mux2h _09955_ (
    .a(\DFF_484.Q ),
    .b(_01934_),
    .s(_00376_),
    .y(_04248_)
  );
  al_mux2h _09956_ (
    .a(\DFF_298.Q ),
    .b(_04248_),
    .s(g35),
    .y(\DFF_484.D )
  );
  al_nand3ftt _09957_ (
    .a(\DFF_587.Q ),
    .b(\DFF_473.Q ),
    .c(\DFF_467.Q ),
    .y(_04249_)
  );
  al_aoi21ftf _09958_ (
    .a(\DFF_156.Q ),
    .b(_04249_),
    .c(g35),
    .y(_04250_)
  );
  al_ao21ftf _09959_ (
    .a(_04249_),
    .b(_00499_),
    .c(_04250_),
    .y(_04251_)
  );
  al_ao21ftf _09960_ (
    .a(g35),
    .b(\DFF_1317.Q ),
    .c(_04251_),
    .y(\DFF_156.D )
  );
  al_ao21ftf _09961_ (
    .a(_02803_),
    .b(\DFF_20.Q ),
    .c(_02804_),
    .y(_04252_)
  );
  al_aoi21 _09962_ (
    .a(\DFF_20.Q ),
    .b(g35),
    .c(\DFF_104.Q ),
    .y(_04253_)
  );
  al_aoi21 _09963_ (
    .a(g35),
    .b(_04252_),
    .c(_04253_),
    .y(\DFF_20.D )
  );
  al_nand2 _09964_ (
    .a(\DFF_727.Q ),
    .b(_00642_),
    .y(_04254_)
  );
  al_oai21 _09965_ (
    .a(_00642_),
    .b(_01618_),
    .c(_04254_),
    .y(_04255_)
  );
  al_mux2h _09966_ (
    .a(\DFF_682.Q ),
    .b(_04255_),
    .s(g35),
    .y(\DFF_727.D )
  );
  al_and3 _09967_ (
    .a(\DFF_63.Q ),
    .b(\DFF_358.Q ),
    .c(_00603_),
    .y(_04256_)
  );
  al_or2 _09968_ (
    .a(\DFF_718.Q ),
    .b(_04256_),
    .y(_04257_)
  );
  al_nand3 _09969_ (
    .a(_02227_),
    .b(_04257_),
    .c(_02228_),
    .y(_04258_)
  );
  al_ao21ftf _09970_ (
    .a(g35),
    .b(\DFF_63.Q ),
    .c(_04258_),
    .y(\DFF_718.D )
  );
  al_nand3ftt _09971_ (
    .a(\DFF_453.Q ),
    .b(\DFF_416.Q ),
    .c(g35),
    .y(_04259_)
  );
  al_oa21 _09972_ (
    .a(\DFF_1242.Q ),
    .b(g35),
    .c(_04259_),
    .y(\DFF_453.D )
  );
  al_nor2 _09973_ (
    .a(\DFF_725.Q ),
    .b(g35),
    .y(_04260_)
  );
  al_mux2h _09974_ (
    .a(_02132_),
    .b(_02134_),
    .s(\DFF_725.Q ),
    .y(_04261_)
  );
  al_nand3ftt _09975_ (
    .a(_04261_),
    .b(\DFF_592.Q ),
    .c(_01948_),
    .y(_04262_)
  );
  al_aoi21ftf _09976_ (
    .a(\DFF_592.Q ),
    .b(_04261_),
    .c(g35),
    .y(_04263_)
  );
  al_aoi21 _09977_ (
    .a(_04263_),
    .b(_04262_),
    .c(_04260_),
    .y(\DFF_592.D )
  );
  al_nand3ftt _09978_ (
    .a(_02368_),
    .b(_00499_),
    .c(_00691_),
    .y(_04264_)
  );
  al_ao21ftt _09979_ (
    .a(_02368_),
    .b(_00691_),
    .c(\DFF_340.Q ),
    .y(_04265_)
  );
  al_nand3 _09980_ (
    .a(g35),
    .b(_04264_),
    .c(_04265_),
    .y(_04266_)
  );
  al_ao21ftf _09981_ (
    .a(g35),
    .b(\DFF_587.Q ),
    .c(_04266_),
    .y(\DFF_340.D )
  );
  al_mux2l _09982_ (
    .a(\DFF_1301.Q ),
    .b(\DFF_994.Q ),
    .s(g35),
    .y(\DFF_1301.D )
  );
  al_ao21ttf _09983_ (
    .a(_00793_),
    .b(_00766_),
    .c(\DFF_778.Q ),
    .y(_04267_)
  );
  al_nand2ft _09984_ (
    .a(\DFF_589.Q ),
    .b(g35),
    .y(_04268_)
  );
  al_ao21ftf _09985_ (
    .a(_04268_),
    .b(\DFF_341.Q ),
    .c(_02727_),
    .y(_04269_)
  );
  al_and3ftt _09986_ (
    .a(\DFF_341.Q ),
    .b(_04268_),
    .c(_02727_),
    .y(_04270_)
  );
  al_aoi21 _09987_ (
    .a(_04267_),
    .b(_04269_),
    .c(_04270_),
    .y(\DFF_778.D )
  );
  al_mux2l _09988_ (
    .a(\DFF_1270.Q ),
    .b(\DFF_1067.Q ),
    .s(g35),
    .y(\DFF_1270.D )
  );
  al_nand3 _09989_ (
    .a(_00499_),
    .b(_02624_),
    .c(_01344_),
    .y(_04271_)
  );
  al_ao21 _09990_ (
    .a(_01344_),
    .b(_02624_),
    .c(\DFF_483.Q ),
    .y(_04272_)
  );
  al_nand3 _09991_ (
    .a(g35),
    .b(_04272_),
    .c(_04271_),
    .y(_04273_)
  );
  al_ao21ftf _09992_ (
    .a(g35),
    .b(\DFF_158.Q ),
    .c(_04273_),
    .y(\DFF_483.D )
  );
  al_inv _09993_ (
    .a(\DFF_297.Q ),
    .y(_04274_)
  );
  al_oa21ftf _09994_ (
    .a(_02654_),
    .b(_01394_),
    .c(_00066_),
    .y(_04275_)
  );
  al_ao21ttf _09995_ (
    .a(_04274_),
    .b(_02655_),
    .c(_04275_),
    .y(_04276_)
  );
  al_ao21ftf _09996_ (
    .a(g35),
    .b(\DFF_1337.Q ),
    .c(_04276_),
    .y(\DFF_681.D )
  );
  al_nand2 _09997_ (
    .a(\DFF_1189.Q ),
    .b(_00966_),
    .y(_04277_)
  );
  al_or2 _09998_ (
    .a(\DFF_1189.Q ),
    .b(_00966_),
    .y(_04278_)
  );
  al_nand3 _09999_ (
    .a(_04277_),
    .b(_04278_),
    .c(_02741_),
    .y(_04279_)
  );
  al_ao21ftf _10000_ (
    .a(g35),
    .b(\DFF_1159.Q ),
    .c(_04279_),
    .y(\DFF_1189.D )
  );
  al_or2 _10001_ (
    .a(_00066_),
    .b(_02655_),
    .y(_04280_)
  );
  al_and3fft _10002_ (
    .a(_00066_),
    .b(_01394_),
    .c(_04274_),
    .y(_04281_)
  );
  al_aoi21 _10003_ (
    .a(_02657_),
    .b(_04280_),
    .c(_04281_),
    .y(\DFF_297.D )
  );
  al_nand3 _10004_ (
    .a(_00499_),
    .b(_01840_),
    .c(_01976_),
    .y(_04282_)
  );
  al_ao21 _10005_ (
    .a(_01976_),
    .b(_01840_),
    .c(\DFF_923.Q ),
    .y(_04283_)
  );
  al_nand3 _10006_ (
    .a(g35),
    .b(_04283_),
    .c(_04282_),
    .y(_04284_)
  );
  al_ao21ftf _10007_ (
    .a(g35),
    .b(\DFF_638.Q ),
    .c(_04284_),
    .y(\DFF_923.D )
  );
  al_ao21 _10008_ (
    .a(\DFF_461.Q ),
    .b(_00459_),
    .c(\DFF_604.Q ),
    .y(_04285_)
  );
  al_aoi21ttf _10009_ (
    .a(\DFF_461.Q ),
    .b(_00460_),
    .c(_04285_),
    .y(_04286_)
  );
  al_and3ftt _10010_ (
    .a(_00460_),
    .b(_04286_),
    .c(_00745_),
    .y(_04287_)
  );
  al_mux2h _10011_ (
    .a(\DFF_461.Q ),
    .b(_04287_),
    .s(g35),
    .y(\DFF_604.D )
  );
  al_nor2 _10012_ (
    .a(\DFF_335.Q ),
    .b(g35),
    .y(_04288_)
  );
  al_or3fft _10013_ (
    .a(\DFF_381.Q ),
    .b(_01642_),
    .c(_04071_),
    .y(_04289_)
  );
  al_aoi21ftf _10014_ (
    .a(\DFF_381.Q ),
    .b(_04071_),
    .c(g35),
    .y(_04290_)
  );
  al_aoi21 _10015_ (
    .a(_04289_),
    .b(_04290_),
    .c(_04288_),
    .y(\DFF_381.D )
  );
  al_aoi21ftt _10016_ (
    .a(_00844_),
    .b(_00843_),
    .c(_00845_),
    .y(_04291_)
  );
  al_mux2h _10017_ (
    .a(\DFF_979.Q ),
    .b(_04291_),
    .s(g35),
    .y(\DFF_788.D )
  );
  al_and2 _10018_ (
    .a(\DFF_935.Q ),
    .b(_02146_),
    .y(\DFF_130.D )
  );
  al_mux2l _10019_ (
    .a(\DFF_435.Q ),
    .b(\DFF_1114.Q ),
    .s(_02454_),
    .y(\DFF_1114.D )
  );
  al_mux2l _10020_ (
    .a(\DFF_766.Q ),
    .b(\DFF_855.Q ),
    .s(g35),
    .y(\DFF_766.D )
  );
  al_nand3ftt _10021_ (
    .a(\DFF_749.Q ),
    .b(g91),
    .c(g35),
    .y(_04292_)
  );
  al_oa21 _10022_ (
    .a(g35),
    .b(\DFF_757.Q ),
    .c(_04292_),
    .y(\DFF_749.D )
  );
  al_ao21 _10023_ (
    .a(\DFF_438.Q ),
    .b(g35),
    .c(_02763_),
    .y(_04293_)
  );
  al_and3 _10024_ (
    .a(\DFF_438.Q ),
    .b(g35),
    .c(_02763_),
    .y(_04294_)
  );
  al_and2ft _10025_ (
    .a(_04294_),
    .b(_04293_),
    .y(\DFF_438.D )
  );
  al_nor2 _10026_ (
    .a(\DFF_671.Q ),
    .b(g35),
    .y(_04295_)
  );
  al_nand3 _10027_ (
    .a(\DFF_671.Q ),
    .b(_01150_),
    .c(_02593_),
    .y(_04296_)
  );
  al_oa21ftf _10028_ (
    .a(\DFF_996.Q ),
    .b(_01150_),
    .c(_00066_),
    .y(_04297_)
  );
  al_aoi21 _10029_ (
    .a(_04297_),
    .b(_04296_),
    .c(_04295_),
    .y(\DFF_996.D )
  );
  al_oa21ftf _10030_ (
    .a(_01999_),
    .b(_01995_),
    .c(_01997_),
    .y(_04298_)
  );
  al_nand3 _10031_ (
    .a(\DFF_1015.Q ),
    .b(_02004_),
    .c(_02006_),
    .y(_04299_)
  );
  al_nand3ftt _10032_ (
    .a(_01995_),
    .b(_01999_),
    .c(_04299_),
    .y(_04300_)
  );
  al_nand3fft _10033_ (
    .a(_00066_),
    .b(_04298_),
    .c(_04300_),
    .y(_04301_)
  );
  al_ao21ftf _10034_ (
    .a(g35),
    .b(\DFF_1246.Q ),
    .c(_04301_),
    .y(\DFF_1015.D )
  );
  al_mux2h _10035_ (
    .a(\DFF_1390.Q ),
    .b(_01348_),
    .s(g35),
    .y(_04302_)
  );
  al_nor3fft _10036_ (
    .a(\DFF_900.Q ),
    .b(g35),
    .c(_01348_),
    .y(_04303_)
  );
  al_ao21 _10037_ (
    .a(_04302_),
    .b(_01827_),
    .c(_04303_),
    .y(\DFF_900.D )
  );
  al_oa21ftf _10038_ (
    .a(_01873_),
    .b(_01870_),
    .c(_02581_),
    .y(_04304_)
  );
  al_nand3 _10039_ (
    .a(\DFF_518.Q ),
    .b(_01335_),
    .c(_01337_),
    .y(_04305_)
  );
  al_nand3ftt _10040_ (
    .a(_01870_),
    .b(_01873_),
    .c(_04305_),
    .y(_04306_)
  );
  al_nand3fft _10041_ (
    .a(_00066_),
    .b(_04304_),
    .c(_04306_),
    .y(_04307_)
  );
  al_ao21ftf _10042_ (
    .a(g35),
    .b(\DFF_665.Q ),
    .c(_04307_),
    .y(\DFF_518.D )
  );
  al_nand3 _10043_ (
    .a(_00499_),
    .b(_02113_),
    .c(_02682_),
    .y(_04308_)
  );
  al_ao21 _10044_ (
    .a(_02113_),
    .b(_02682_),
    .c(\DFF_1210.Q ),
    .y(_04309_)
  );
  al_nand3 _10045_ (
    .a(g35),
    .b(_04308_),
    .c(_04309_),
    .y(_04310_)
  );
  al_ao21ftf _10046_ (
    .a(g35),
    .b(\DFF_9.Q ),
    .c(_04310_),
    .y(\DFF_1210.D )
  );
  al_nand3ftt _10047_ (
    .a(\DFF_1014.Q ),
    .b(\DFF_686.Q ),
    .c(g35),
    .y(_04311_)
  );
  al_ao21ftf _10048_ (
    .a(g35),
    .b(\DFF_1014.Q ),
    .c(_04311_),
    .y(\DFF_240.D )
  );
  al_mux2l _10049_ (
    .a(\DFF_972.Q ),
    .b(\DFF_542.Q ),
    .s(_01174_),
    .y(\DFF_542.D )
  );
  al_mux2l _10050_ (
    .a(\DFF_430.Q ),
    .b(\DFF_11.Q ),
    .s(_01109_),
    .y(\DFF_11.D )
  );
  al_nand3 _10051_ (
    .a(_00499_),
    .b(_00706_),
    .c(_02682_),
    .y(_04312_)
  );
  al_ao21 _10052_ (
    .a(_00706_),
    .b(_02682_),
    .c(\DFF_1280.Q ),
    .y(_04313_)
  );
  al_nand3 _10053_ (
    .a(g35),
    .b(_04313_),
    .c(_04312_),
    .y(_04314_)
  );
  al_ao21ftf _10054_ (
    .a(g35),
    .b(\DFF_134.Q ),
    .c(_04314_),
    .y(\DFF_1280.D )
  );
  al_mux2l _10055_ (
    .a(\DFF_1193.Q ),
    .b(\DFF_677.Q ),
    .s(g35),
    .y(\DFF_1193.D )
  );
  al_nand2 _10056_ (
    .a(\DFF_1061.Q ),
    .b(\DFF_612.Q ),
    .y(_04315_)
  );
  al_oai21ttf _10057_ (
    .a(\DFF_824.Q ),
    .b(_04315_),
    .c(_00066_),
    .y(_04316_)
  );
  al_inv _10058_ (
    .a(\DFF_842.Q ),
    .y(_04317_)
  );
  al_mux2l _10059_ (
    .a(\DFF_956.Q ),
    .b(_04317_),
    .s(_04315_),
    .y(_04318_)
  );
  al_mux2l _10060_ (
    .a(\DFF_842.Q ),
    .b(_04318_),
    .s(_04316_),
    .y(\DFF_956.D )
  );
  al_and3ftt _10061_ (
    .a(_01122_),
    .b(_00604_),
    .c(_00326_),
    .y(_04319_)
  );
  al_or2 _10062_ (
    .a(\DFF_1009.Q ),
    .b(_04319_),
    .y(_04320_)
  );
  al_oai21ftt _10063_ (
    .a(\DFF_620.Q ),
    .b(\DFF_759.Q ),
    .c(\DFF_1181.Q ),
    .y(_04321_)
  );
  al_or3ftt _10064_ (
    .a(\DFF_620.Q ),
    .b(\DFF_759.Q ),
    .c(\DFF_1181.Q ),
    .y(_04322_)
  );
  al_nand3 _10065_ (
    .a(_04321_),
    .b(_04322_),
    .c(_04319_),
    .y(_04323_)
  );
  al_nand3 _10066_ (
    .a(g35),
    .b(_04323_),
    .c(_04320_),
    .y(_04324_)
  );
  al_ao21ftf _10067_ (
    .a(g35),
    .b(\DFF_111.Q ),
    .c(_04324_),
    .y(\DFF_1009.D )
  );
  al_nor2 _10068_ (
    .a(\DFF_265.Q ),
    .b(g35),
    .y(_04325_)
  );
  al_nand3 _10069_ (
    .a(\DFF_265.Q ),
    .b(_00974_),
    .c(_02883_),
    .y(_04326_)
  );
  al_oa21ftf _10070_ (
    .a(\DFF_886.Q ),
    .b(_00974_),
    .c(_00066_),
    .y(_04327_)
  );
  al_aoi21 _10071_ (
    .a(_04327_),
    .b(_04326_),
    .c(_04325_),
    .y(\DFF_886.D )
  );
  al_and2ft _10072_ (
    .a(\DFF_509.Q ),
    .b(g35),
    .y(\DFF_203.D )
  );
  al_ao21ftt _10073_ (
    .a(g35),
    .b(\DFF_1425.Q ),
    .c(\DFF_1425.D ),
    .y(\DFF_350.D )
  );
  al_nor3ftt _10074_ (
    .a(\DFF_826.Q ),
    .b(_00499_),
    .c(g26801),
    .y(_04328_)
  );
  al_oa21ftt _10075_ (
    .a(\DFF_826.Q ),
    .b(g26801),
    .c(_00499_),
    .y(_04329_)
  );
  al_nor3ftt _10076_ (
    .a(g35),
    .b(_04328_),
    .c(_04329_),
    .y(\DFF_826.D )
  );
  al_ao21 _10077_ (
    .a(g35),
    .b(\DFF_1055.Q ),
    .c(\DFF_694.Q ),
    .y(_04330_)
  );
  al_aoi21 _10078_ (
    .a(g35),
    .b(_04052_),
    .c(_04330_),
    .y(_04331_)
  );
  al_ao21ttf _10079_ (
    .a(_02339_),
    .b(_02338_),
    .c(\DFF_987.Q ),
    .y(_04332_)
  );
  al_nand2 _10080_ (
    .a(\DFF_694.Q ),
    .b(\DFF_1055.Q ),
    .y(_04333_)
  );
  al_oa21ftf _10081_ (
    .a(_04333_),
    .b(_04052_),
    .c(_00066_),
    .y(_04334_)
  );
  al_aoi21 _10082_ (
    .a(_04332_),
    .b(_04334_),
    .c(_04331_),
    .y(\DFF_987.D )
  );
  al_oa21ftt _10083_ (
    .a(\DFF_890.Q ),
    .b(\DFF_189.Q ),
    .c(\DFF_623.Q ),
    .y(_04335_)
  );
  al_ao21ttf _10084_ (
    .a(\DFF_727.Q ),
    .b(\DFF_562.Q ),
    .c(_04335_),
    .y(_04336_)
  );
  al_aoi21 _10085_ (
    .a(\DFF_61.Q ),
    .b(\DFF_189.Q ),
    .c(\DFF_623.Q ),
    .y(_04337_)
  );
  al_ao21ftf _10086_ (
    .a(\DFF_562.Q ),
    .b(\DFF_960.Q ),
    .c(_04337_),
    .y(_04338_)
  );
  al_and3ftt _10087_ (
    .a(\DFF_189.Q ),
    .b(\DFF_1097.Q ),
    .c(\DFF_562.Q ),
    .y(_04339_)
  );
  al_ao21 _10088_ (
    .a(\DFF_1380.Q ),
    .b(_00444_),
    .c(_04339_),
    .y(_04340_)
  );
  al_ao21 _10089_ (
    .a(_04338_),
    .b(_04336_),
    .c(_04340_),
    .y(_04341_)
  );
  al_mux2l _10090_ (
    .a(_04341_),
    .b(\DFF_1082.Q ),
    .s(_00758_),
    .y(_04342_)
  );
  al_mux2h _10091_ (
    .a(\DFF_562.Q ),
    .b(_04342_),
    .s(g35),
    .y(\DFF_1082.D )
  );
  al_nand3 _10092_ (
    .a(_00499_),
    .b(_00567_),
    .c(_01952_),
    .y(_04343_)
  );
  al_ao21 _10093_ (
    .a(_01952_),
    .b(_00567_),
    .c(\DFF_187.Q ),
    .y(_04344_)
  );
  al_nand3 _10094_ (
    .a(g35),
    .b(_04344_),
    .c(_04343_),
    .y(_04345_)
  );
  al_ao21ftf _10095_ (
    .a(g35),
    .b(\DFF_1212.Q ),
    .c(_04345_),
    .y(\DFF_187.D )
  );
  al_and3 _10096_ (
    .a(\DFF_720.Q ),
    .b(_02278_),
    .c(_01261_),
    .y(_04346_)
  );
  al_oa21ftf _10097_ (
    .a(_00636_),
    .b(_04346_),
    .c(_00066_),
    .y(_04347_)
  );
  al_ao21ftf _10098_ (
    .a(_00636_),
    .b(_04346_),
    .c(_04347_),
    .y(_04348_)
  );
  al_ao21ftf _10099_ (
    .a(g35),
    .b(\DFF_720.Q ),
    .c(_04348_),
    .y(\DFF_1323.D )
  );
  al_and2ft _10100_ (
    .a(g35),
    .b(\DFF_140.Q ),
    .y(_04349_)
  );
  al_or2 _10101_ (
    .a(\DFF_140.Q ),
    .b(_01448_),
    .y(_04350_)
  );
  al_aoi21ftf _10102_ (
    .a(_01445_),
    .b(_01451_),
    .c(_04350_),
    .y(_04351_)
  );
  al_ao21ftf _10103_ (
    .a(_01446_),
    .b(_01455_),
    .c(_04351_),
    .y(_04352_)
  );
  al_oa21ftf _10104_ (
    .a(\DFF_586.Q ),
    .b(_04351_),
    .c(_00066_),
    .y(_04353_)
  );
  al_ao21 _10105_ (
    .a(_04352_),
    .b(_04353_),
    .c(_04349_),
    .y(\DFF_586.D )
  );
  al_nand3 _10106_ (
    .a(_00499_),
    .b(_01170_),
    .c(_02625_),
    .y(_04354_)
  );
  al_ao21 _10107_ (
    .a(_01170_),
    .b(_02625_),
    .c(\DFF_1123.Q ),
    .y(_04355_)
  );
  al_nand3 _10108_ (
    .a(g35),
    .b(_04355_),
    .c(_04354_),
    .y(_04356_)
  );
  al_ao21ftf _10109_ (
    .a(g35),
    .b(\DFF_59.Q ),
    .c(_04356_),
    .y(\DFF_1123.D )
  );
  al_nand3 _10110_ (
    .a(_00499_),
    .b(_01772_),
    .c(_01744_),
    .y(_04357_)
  );
  al_ao21 _10111_ (
    .a(_01744_),
    .b(_01772_),
    .c(\DFF_1297.Q ),
    .y(_04358_)
  );
  al_nand3 _10112_ (
    .a(g35),
    .b(_04358_),
    .c(_04357_),
    .y(_04359_)
  );
  al_ao21ftf _10113_ (
    .a(g35),
    .b(\DFF_895.Q ),
    .c(_04359_),
    .y(\DFF_1297.D )
  );
  al_and2 _10114_ (
    .a(g35),
    .b(\DFF_1067.Q ),
    .y(\DFF_1067.D )
  );
  al_nor2 _10115_ (
    .a(g35),
    .b(\DFF_658.Q ),
    .y(_04360_)
  );
  al_nand3 _10116_ (
    .a(\DFF_769.Q ),
    .b(_01282_),
    .c(_02639_),
    .y(_04361_)
  );
  al_oa21ftf _10117_ (
    .a(\DFF_1141.Q ),
    .b(_01282_),
    .c(_00066_),
    .y(_04362_)
  );
  al_aoi21 _10118_ (
    .a(_04362_),
    .b(_04361_),
    .c(_04360_),
    .y(\DFF_1141.D )
  );
  al_nand2 _10119_ (
    .a(g35),
    .b(_00564_),
    .y(_04363_)
  );
  al_mux2l _10120_ (
    .a(\DFF_768.Q ),
    .b(\DFF_6.Q ),
    .s(_04363_),
    .y(\DFF_6.D )
  );
  al_nand2 _10121_ (
    .a(\DFF_963.Q ),
    .b(_01461_),
    .y(_04364_)
  );
  al_nand2 _10122_ (
    .a(\DFF_339.Q ),
    .b(\DFF_1241.Q ),
    .y(_04365_)
  );
  al_aoi21 _10123_ (
    .a(_04365_),
    .b(_04364_),
    .c(_01462_),
    .y(_04366_)
  );
  al_mux2h _10124_ (
    .a(\DFF_963.Q ),
    .b(_04366_),
    .s(g35),
    .y(\DFF_1241.D )
  );
  al_nand2 _10125_ (
    .a(\DFF_354.Q ),
    .b(g35),
    .y(_04367_)
  );
  al_aoi21ftt _10126_ (
    .a(\DFF_605.Q ),
    .b(_04367_),
    .c(_02283_),
    .y(\DFF_354.D )
  );
  al_or3ftt _10127_ (
    .a(_02157_),
    .b(\DFF_757.Q ),
    .c(_02152_),
    .y(_04368_)
  );
  al_mux2h _10128_ (
    .a(\DFF_223.Q ),
    .b(_04368_),
    .s(g35),
    .y(\DFF_757.D )
  );
  al_and2ft _10129_ (
    .a(g35),
    .b(\DFF_1132.Q ),
    .y(_04369_)
  );
  al_aoi21ttf _10130_ (
    .a(\DFF_1132.Q ),
    .b(_01338_),
    .c(_02583_),
    .y(_04370_)
  );
  al_ao21 _10131_ (
    .a(_04370_),
    .b(_02565_),
    .c(_02582_),
    .y(_04371_)
  );
  al_aoi21 _10132_ (
    .a(_02582_),
    .b(_04370_),
    .c(_00066_),
    .y(_04372_)
  );
  al_ao21 _10133_ (
    .a(_04372_),
    .b(_04371_),
    .c(_04369_),
    .y(\DFF_665.D )
  );
  al_ao21ftf _10134_ (
    .a(g35),
    .b(\DFF_576.Q ),
    .c(_01743_),
    .y(\DFF_125.D )
  );
  al_mux2l _10135_ (
    .a(\DFF_11.Q ),
    .b(\DFF_629.Q ),
    .s(_01109_),
    .y(\DFF_629.D )
  );
  al_aoi21 _10136_ (
    .a(\DFF_831.Q ),
    .b(g35),
    .c(\DFF_320.Q ),
    .y(_04373_)
  );
  al_and2 _10137_ (
    .a(g35),
    .b(\DFF_320.Q ),
    .y(_04374_)
  );
  al_aoi21 _10138_ (
    .a(\DFF_831.Q ),
    .b(_04374_),
    .c(_04373_),
    .y(\DFF_1384.D )
  );
  al_aoi21 _10139_ (
    .a(\DFF_833.Q ),
    .b(_01956_),
    .c(_00066_),
    .y(_04375_)
  );
  al_and2ft _10140_ (
    .a(g35),
    .b(\DFF_731.Q ),
    .y(_04376_)
  );
  al_ao21 _10141_ (
    .a(_01956_),
    .b(_04125_),
    .c(\DFF_833.Q ),
    .y(_04377_)
  );
  al_ao21 _10142_ (
    .a(_04375_),
    .b(_04377_),
    .c(_04376_),
    .y(\DFF_833.D )
  );
  al_aoi21 _10143_ (
    .a(\DFF_1184.Q ),
    .b(_01126_),
    .c(_00066_),
    .y(_04378_)
  );
  al_oai21 _10144_ (
    .a(\DFF_1184.Q ),
    .b(_01126_),
    .c(_04378_),
    .y(_04379_)
  );
  al_aoi21ftf _10145_ (
    .a(\DFF_1179.Q ),
    .b(_00066_),
    .c(_04379_),
    .y(\DFF_1184.D )
  );
  al_mux2l _10146_ (
    .a(\DFF_136.Q ),
    .b(\DFF_300.Q ),
    .s(_02170_),
    .y(\DFF_300.D )
  );
  al_oai21ftt _10147_ (
    .a(g35),
    .b(_02905_),
    .c(\DFF_1146.Q ),
    .y(_04380_)
  );
  al_ao21ftf _10148_ (
    .a(_00066_),
    .b(\DFF_613.Q ),
    .c(_04380_),
    .y(\DFF_482.D )
  );
  al_and3ftt _10149_ (
    .a(\DFF_925.Q ),
    .b(_02803_),
    .c(_03112_),
    .y(\DFF_925.D )
  );
  al_nand3fft _10150_ (
    .a(\DFF_1092.Q ),
    .b(\DFF_403.Q ),
    .c(_00516_),
    .y(_04381_)
  );
  al_ao21ftf _10151_ (
    .a(\DFF_1092.Q ),
    .b(_00516_),
    .c(\DFF_403.Q ),
    .y(_04382_)
  );
  al_nand3 _10152_ (
    .a(_03902_),
    .b(_04381_),
    .c(_04382_),
    .y(_04383_)
  );
  al_ao21 _10153_ (
    .a(_03902_),
    .b(_02800_),
    .c(\DFF_193.Q ),
    .y(_04384_)
  );
  al_nand3 _10154_ (
    .a(g35),
    .b(_04384_),
    .c(_04383_),
    .y(_04385_)
  );
  al_ao21ftf _10155_ (
    .a(_01259_),
    .b(_00066_),
    .c(_04385_),
    .y(\DFF_193.D )
  );
  al_and2 _10156_ (
    .a(g35),
    .b(\DFF_482.Q ),
    .y(_04386_)
  );
  al_or3fft _10157_ (
    .a(_00503_),
    .b(_04386_),
    .c(_00505_),
    .y(_04387_)
  );
  al_nand2ft _10158_ (
    .a(\DFF_1002.Q ),
    .b(_04387_),
    .y(\DFF_1146.D )
  );
  al_nand2ft _10159_ (
    .a(g35),
    .b(\DFF_198.Q ),
    .y(_04388_)
  );
  al_ao21ftf _10160_ (
    .a(\DFF_683.Q ),
    .b(_03029_),
    .c(_04388_),
    .y(\DFF_1130.D )
  );
  al_mux2l _10161_ (
    .a(\DFF_648.Q ),
    .b(\DFF_152.Q ),
    .s(_01557_),
    .y(_04389_)
  );
  al_mux2h _10162_ (
    .a(\DFF_496.Q ),
    .b(_04389_),
    .s(g35),
    .y(\DFF_648.D )
  );
  al_nand3fft _10163_ (
    .a(\DFF_1092.Q ),
    .b(\DFF_1323.Q ),
    .c(_00516_),
    .y(_04390_)
  );
  al_ao21ftf _10164_ (
    .a(\DFF_1092.Q ),
    .b(_00516_),
    .c(\DFF_1323.Q ),
    .y(_04391_)
  );
  al_nand3 _10165_ (
    .a(_02278_),
    .b(_04390_),
    .c(_04391_),
    .y(_04392_)
  );
  al_ao21 _10166_ (
    .a(_02278_),
    .b(_02800_),
    .c(\DFF_720.Q ),
    .y(_04393_)
  );
  al_nand3 _10167_ (
    .a(g35),
    .b(_04393_),
    .c(_04392_),
    .y(_04394_)
  );
  al_ao21ftf _10168_ (
    .a(_03613_),
    .b(_00066_),
    .c(_04394_),
    .y(\DFF_720.D )
  );
  al_nand3ftt _10169_ (
    .a(_00497_),
    .b(_00499_),
    .c(_01701_),
    .y(_04395_)
  );
  al_ao21ftt _10170_ (
    .a(_00497_),
    .b(_01701_),
    .c(\DFF_151.Q ),
    .y(_04396_)
  );
  al_nand3 _10171_ (
    .a(g35),
    .b(_04395_),
    .c(_04396_),
    .y(_04397_)
  );
  al_ao21ftf _10172_ (
    .a(g35),
    .b(\DFF_84.Q ),
    .c(_04397_),
    .y(\DFF_151.D )
  );
  al_nand3 _10173_ (
    .a(_00499_),
    .b(_00508_),
    .c(_01105_),
    .y(_04398_)
  );
  al_ao21 _10174_ (
    .a(_00508_),
    .b(_01105_),
    .c(\DFF_345.Q ),
    .y(_04399_)
  );
  al_nand3 _10175_ (
    .a(g35),
    .b(_04399_),
    .c(_04398_),
    .y(_04400_)
  );
  al_ao21ftf _10176_ (
    .a(g35),
    .b(\DFF_730.Q ),
    .c(_04400_),
    .y(\DFF_345.D )
  );
  al_nand3 _10177_ (
    .a(_00499_),
    .b(_01354_),
    .c(_02625_),
    .y(_04401_)
  );
  al_ao21 _10178_ (
    .a(_01354_),
    .b(_02625_),
    .c(\DFF_1307.Q ),
    .y(_04402_)
  );
  al_nand3 _10179_ (
    .a(g35),
    .b(_04402_),
    .c(_04401_),
    .y(_04403_)
  );
  al_ao21ftf _10180_ (
    .a(g35),
    .b(\DFF_904.Q ),
    .c(_04403_),
    .y(\DFF_1307.D )
  );
  al_and2ft _10181_ (
    .a(g35),
    .b(\DFF_1199.Q ),
    .y(_04404_)
  );
  al_nand2ft _10182_ (
    .a(\DFF_892.Q ),
    .b(_01990_),
    .y(_04405_)
  );
  al_aoi21ftf _10183_ (
    .a(_03812_),
    .b(_02036_),
    .c(_01984_),
    .y(_04406_)
  );
  al_ao21 _10184_ (
    .a(_04405_),
    .b(_04406_),
    .c(_04404_),
    .y(\DFF_892.D )
  );
  al_or3 _10185_ (
    .a(\DFF_541.Q ),
    .b(g73),
    .c(g72),
    .y(_04407_)
  );
  al_oai21ftt _10186_ (
    .a(\DFF_771.Q ),
    .b(g72),
    .c(g73),
    .y(_04408_)
  );
  al_oai21ftt _10187_ (
    .a(g72),
    .b(\DFF_648.Q ),
    .c(g35),
    .y(_04409_)
  );
  al_nand3ftt _10188_ (
    .a(_04409_),
    .b(_04407_),
    .c(_04408_),
    .y(_04410_)
  );
  al_ao21ftf _10189_ (
    .a(g35),
    .b(\DFF_357.Q ),
    .c(_04410_),
    .y(\DFF_143.D )
  );
  al_mux2l _10190_ (
    .a(\DFF_664.Q ),
    .b(\DFF_1298.Q ),
    .s(g35),
    .y(\DFF_1414.D )
  );
  al_oai21ftf _10191_ (
    .a(\DFF_74.Q ),
    .b(_02250_),
    .c(\DFF_50.Q ),
    .y(_04411_)
  );
  al_nand3fft _10192_ (
    .a(_01837_),
    .b(_00952_),
    .c(_04411_),
    .y(_04412_)
  );
  al_ao21ftf _10193_ (
    .a(g35),
    .b(\DFF_74.Q ),
    .c(_04412_),
    .y(\DFF_50.D )
  );
  al_mux2l _10194_ (
    .a(\DFF_1151.Q ),
    .b(\DFF_1282.Q ),
    .s(g35),
    .y(\DFF_1151.D )
  );
  al_ao21ftt _10195_ (
    .a(\DFF_425.Q ),
    .b(_00550_),
    .c(\DFF_534.Q ),
    .y(_04413_)
  );
  al_and2ft _10196_ (
    .a(g35),
    .b(\DFF_470.Q ),
    .y(_04414_)
  );
  al_ao21 _10197_ (
    .a(_00552_),
    .b(_04413_),
    .c(_04414_),
    .y(\DFF_534.D )
  );
  al_mux2l _10198_ (
    .a(\DFF_683.Q ),
    .b(\DFF_1130.Q ),
    .s(\DFF_952.Q ),
    .y(_04415_)
  );
  al_aoi21 _10199_ (
    .a(\DFF_878.Q ),
    .b(_04415_),
    .c(\DFF_782.Q ),
    .y(_04416_)
  );
  al_oai21 _10200_ (
    .a(\DFF_878.Q ),
    .b(_04415_),
    .c(_04416_),
    .y(_04417_)
  );
  al_ao21ttf _10201_ (
    .a(_00465_),
    .b(_04417_),
    .c(_02338_),
    .y(_04418_)
  );
  al_or2 _10202_ (
    .a(\DFF_782.Q ),
    .b(_02338_),
    .y(_04419_)
  );
  al_and3 _10203_ (
    .a(g35),
    .b(_04418_),
    .c(_04419_),
    .y(\DFF_782.D )
  );
  al_and2 _10204_ (
    .a(_01414_),
    .b(_01282_),
    .y(_04420_)
  );
  al_nor2 _10205_ (
    .a(_01413_),
    .b(_01282_),
    .y(_04421_)
  );
  al_ao21 _10206_ (
    .a(_04420_),
    .b(_02639_),
    .c(_04421_),
    .y(_04422_)
  );
  al_and3ftt _10207_ (
    .a(_00877_),
    .b(g35),
    .c(_04422_),
    .y(\DFF_769.D )
  );
  al_nor2 _10208_ (
    .a(g35),
    .b(\DFF_943.Q ),
    .y(_04423_)
  );
  al_nand3 _10209_ (
    .a(\DFF_209.Q ),
    .b(_00526_),
    .c(_02650_),
    .y(_04424_)
  );
  al_oa21ftf _10210_ (
    .a(\DFF_1010.Q ),
    .b(_00526_),
    .c(_00066_),
    .y(_04425_)
  );
  al_aoi21 _10211_ (
    .a(_04425_),
    .b(_04424_),
    .c(_04423_),
    .y(\DFF_1010.D )
  );
  al_ao21ftf _10212_ (
    .a(\DFF_597.Q ),
    .b(\DFF_1390.Q ),
    .c(_01175_),
    .y(_04426_)
  );
  al_ao21ftf _10213_ (
    .a(g35),
    .b(\DFF_1253.Q ),
    .c(_04426_),
    .y(\DFF_597.D )
  );
  al_nand3fft _10214_ (
    .a(\DFF_802.Q ),
    .b(_00066_),
    .c(_00935_),
    .y(_04427_)
  );
  al_ao21ftf _10215_ (
    .a(g35),
    .b(\DFF_128.Q ),
    .c(_04427_),
    .y(\DFF_802.D )
  );
  al_nor2 _10216_ (
    .a(\DFF_500.Q ),
    .b(g35),
    .y(_04428_)
  );
  al_nand3 _10217_ (
    .a(\DFF_500.Q ),
    .b(_01889_),
    .c(_03061_),
    .y(_04429_)
  );
  al_oa21ftf _10218_ (
    .a(\DFF_18.Q ),
    .b(_01889_),
    .c(_00066_),
    .y(_04430_)
  );
  al_aoi21 _10219_ (
    .a(_04430_),
    .b(_04429_),
    .c(_04428_),
    .y(\DFF_18.D )
  );
  al_nand3ftt _10220_ (
    .a(_03064_),
    .b(_02113_),
    .c(_00499_),
    .y(_04431_)
  );
  al_ao21ftt _10221_ (
    .a(_03064_),
    .b(_02113_),
    .c(\DFF_1208.Q ),
    .y(_04432_)
  );
  al_nand3 _10222_ (
    .a(g35),
    .b(_04431_),
    .c(_04432_),
    .y(_04433_)
  );
  al_ao21ftf _10223_ (
    .a(g35),
    .b(\DFF_1351.Q ),
    .c(_04433_),
    .y(\DFF_1208.D )
  );
  al_and2ft _10224_ (
    .a(g35),
    .b(\DFF_840.Q ),
    .y(_04434_)
  );
  al_ao21 _10225_ (
    .a(_02064_),
    .b(_04039_),
    .c(\DFF_1347.Q ),
    .y(_04435_)
  );
  al_aoi21 _10226_ (
    .a(\DFF_1347.Q ),
    .b(_02064_),
    .c(_00066_),
    .y(_04436_)
  );
  al_ao21 _10227_ (
    .a(_04436_),
    .b(_04435_),
    .c(_04434_),
    .y(\DFF_1347.D )
  );
  al_nand3 _10228_ (
    .a(_00499_),
    .b(_00591_),
    .c(_02871_),
    .y(_04437_)
  );
  al_ao21 _10229_ (
    .a(_02871_),
    .b(_00591_),
    .c(\DFF_854.Q ),
    .y(_04438_)
  );
  al_nand3 _10230_ (
    .a(g35),
    .b(_04438_),
    .c(_04437_),
    .y(_04439_)
  );
  al_ao21ftf _10231_ (
    .a(g35),
    .b(\DFF_17.Q ),
    .c(_04439_),
    .y(\DFF_854.D )
  );
  al_ao21ftt _10232_ (
    .a(_02788_),
    .b(_00549_),
    .c(\DFF_951.Q ),
    .y(_04440_)
  );
  al_ao21 _10233_ (
    .a(_04440_),
    .b(_02129_),
    .c(_01963_),
    .y(_04441_)
  );
  al_aoi21ftf _10234_ (
    .a(\DFF_428.Q ),
    .b(_00066_),
    .c(_04441_),
    .y(\DFF_951.D )
  );
  al_nor2 _10235_ (
    .a(g35),
    .b(\DFF_253.Q ),
    .y(_04442_)
  );
  al_oa21ftf _10236_ (
    .a(\DFF_857.Q ),
    .b(_00585_),
    .c(_00066_),
    .y(_04443_)
  );
  al_aoi21 _10237_ (
    .a(_04443_),
    .b(_02417_),
    .c(_04442_),
    .y(\DFF_857.D )
  );
  al_oai21ftf _10238_ (
    .a(\DFF_678.Q ),
    .b(\DFF_458.Q ),
    .c(\DFF_1065.Q ),
    .y(_04444_)
  );
  al_nand3ftt _10239_ (
    .a(\DFF_545.Q ),
    .b(g35),
    .c(_04444_),
    .y(_04445_)
  );
  al_ao21ftf _10240_ (
    .a(g35),
    .b(\DFF_458.Q ),
    .c(_04445_),
    .y(\DFF_1065.D )
  );
  al_mux2l _10241_ (
    .a(\DFF_198.Q ),
    .b(\DFF_732.Q ),
    .s(g35),
    .y(\DFF_371.D )
  );
  al_nand3 _10242_ (
    .a(_00499_),
    .b(_01114_),
    .c(_02871_),
    .y(_04446_)
  );
  al_ao21 _10243_ (
    .a(_01114_),
    .b(_02871_),
    .c(\DFF_920.Q ),
    .y(_04447_)
  );
  al_nand3 _10244_ (
    .a(g35),
    .b(_04447_),
    .c(_04446_),
    .y(_04448_)
  );
  al_ao21ftf _10245_ (
    .a(g35),
    .b(\DFF_241.Q ),
    .c(_04448_),
    .y(\DFF_920.D )
  );
  al_and2ft _10246_ (
    .a(g35),
    .b(\DFF_40.Q ),
    .y(_04449_)
  );
  al_and2 _10247_ (
    .a(_01295_),
    .b(_01296_),
    .y(_04450_)
  );
  al_ao21 _10248_ (
    .a(_04450_),
    .b(_00899_),
    .c(_01294_),
    .y(_04451_)
  );
  al_nand3 _10249_ (
    .a(_01294_),
    .b(_01295_),
    .c(_01296_),
    .y(_04452_)
  );
  al_and2 _10250_ (
    .a(g35),
    .b(_04452_),
    .y(_04453_)
  );
  al_ao21 _10251_ (
    .a(_04453_),
    .b(_04451_),
    .c(_04449_),
    .y(\DFF_712.D )
  );
  al_mux2h _10252_ (
    .a(\DFF_1334.Q ),
    .b(_01641_),
    .s(g35),
    .y(\DFF_548.D )
  );
  al_ao21ftf _10253_ (
    .a(_01460_),
    .b(\DFF_149.Q ),
    .c(_03727_),
    .y(_04454_)
  );
  al_nand3 _10254_ (
    .a(g35),
    .b(_01464_),
    .c(_04454_),
    .y(_04455_)
  );
  al_ao21ftf _10255_ (
    .a(g35),
    .b(\DFF_859.Q ),
    .c(_04455_),
    .y(\DFF_149.D )
  );
  al_oai21 _10256_ (
    .a(_01744_),
    .b(_01773_),
    .c(_03698_),
    .y(_04456_)
  );
  al_ao21ftf _10257_ (
    .a(g35),
    .b(\DFF_244.Q ),
    .c(_04456_),
    .y(\DFF_958.D )
  );
  al_mux2l _10258_ (
    .a(\DFF_677.Q ),
    .b(\DFF_1157.Q ),
    .s(g35),
    .y(\DFF_677.D )
  );
  al_ao21 _10259_ (
    .a(\DFF_94.Q ),
    .b(g35),
    .c(\DFF_880.Q ),
    .y(_04457_)
  );
  al_nand3 _10260_ (
    .a(\DFF_880.Q ),
    .b(\DFF_94.Q ),
    .c(g35),
    .y(_04458_)
  );
  al_and3ftt _10261_ (
    .a(_02714_),
    .b(_04457_),
    .c(_04458_),
    .y(\DFF_94.D )
  );
  al_oa21ttf _10262_ (
    .a(g35),
    .b(\DFF_1041.Q ),
    .c(_04374_),
    .y(\DFF_831.D )
  );
  al_mux2l _10263_ (
    .a(\DFF_822.Q ),
    .b(\DFF_167.Q ),
    .s(_04134_),
    .y(\DFF_167.D )
  );
  al_nand2 _10264_ (
    .a(\DFF_339.Q ),
    .b(\DFF_963.Q ),
    .y(_04459_)
  );
  al_aoi21ftf _10265_ (
    .a(_01461_),
    .b(_04459_),
    .c(_04364_),
    .y(_04460_)
  );
  al_mux2h _10266_ (
    .a(\DFF_94.Q ),
    .b(_04460_),
    .s(g35),
    .y(\DFF_963.D )
  );
  al_ao21ftt _10267_ (
    .a(g35),
    .b(\DFF_456.Q ),
    .c(_03562_),
    .y(_04461_)
  );
  al_mux2l _10268_ (
    .a(_04461_),
    .b(\DFF_1211.Q ),
    .s(_03339_),
    .y(\DFF_1211.D )
  );
  al_and2 _10269_ (
    .a(\DFF_141.Q ),
    .b(g35),
    .y(_04462_)
  );
  al_aoi21ttf _10270_ (
    .a(_04462_),
    .b(_02913_),
    .c(\DFF_1400.Q ),
    .y(\DFF_1285.D )
  );
  al_nand3fft _10271_ (
    .a(\DFF_500.Q ),
    .b(_01885_),
    .c(_01889_),
    .y(_04463_)
  );
  al_aoi21ftf _10272_ (
    .a(\DFF_41.Q ),
    .b(_04463_),
    .c(g35),
    .y(_04464_)
  );
  al_oai21 _10273_ (
    .a(_01892_),
    .b(_04463_),
    .c(_04464_),
    .y(_04465_)
  );
  al_ao21ftf _10274_ (
    .a(g35),
    .b(\DFF_1258.Q ),
    .c(_04465_),
    .y(\DFF_41.D )
  );
  al_nand3 _10275_ (
    .a(\DFF_694.Q ),
    .b(_04052_),
    .c(_03974_),
    .y(_04466_)
  );
  al_ao21 _10276_ (
    .a(\DFF_694.Q ),
    .b(_04052_),
    .c(_03974_),
    .y(_04467_)
  );
  al_nand3 _10277_ (
    .a(g35),
    .b(_04466_),
    .c(_04467_),
    .y(_04468_)
  );
  al_aoi21ftf _10278_ (
    .a(\DFF_1055.Q ),
    .b(_00066_),
    .c(_04468_),
    .y(\DFF_694.D )
  );
  al_ao21ftf _10279_ (
    .a(g35),
    .b(\DFF_701.Q ),
    .c(_02615_),
    .y(_04469_)
  );
  al_oa21 _10280_ (
    .a(\DFF_701.Q ),
    .b(\DFF_939.Q ),
    .c(_04469_),
    .y(\DFF_939.D )
  );
  al_nor2 _10281_ (
    .a(\DFF_1344.Q ),
    .b(g35),
    .y(_04470_)
  );
  al_nand3 _10282_ (
    .a(_00604_),
    .b(_01056_),
    .c(_00452_),
    .y(_04471_)
  );
  al_oai21ftf _10283_ (
    .a(\DFF_794.Q ),
    .b(\DFF_1344.Q ),
    .c(\DFF_379.Q ),
    .y(_04472_)
  );
  al_nand3ftt _10284_ (
    .a(\DFF_1344.Q ),
    .b(\DFF_794.Q ),
    .c(\DFF_379.Q ),
    .y(_04473_)
  );
  al_or3fft _10285_ (
    .a(_04472_),
    .b(_04473_),
    .c(_04471_),
    .y(_04474_)
  );
  al_aoi21 _10286_ (
    .a(\DFF_342.Q ),
    .b(_04471_),
    .c(_00066_),
    .y(_04475_)
  );
  al_aoi21 _10287_ (
    .a(_04474_),
    .b(_04475_),
    .c(_04470_),
    .y(\DFF_342.D )
  );
  al_nand2ft _10288_ (
    .a(g35),
    .b(\DFF_141.Q ),
    .y(_04476_)
  );
  al_ao21ftf _10289_ (
    .a(\DFF_1285.Q ),
    .b(_02914_),
    .c(_04476_),
    .y(\DFF_1400.D )
  );
  al_or3ftt _10290_ (
    .a(\DFF_473.Q ),
    .b(\DFF_587.Q ),
    .c(\DFF_467.Q ),
    .y(_04477_)
  );
  al_aoi21ftf _10291_ (
    .a(\DFF_590.Q ),
    .b(_04477_),
    .c(g35),
    .y(_04478_)
  );
  al_ao21ftf _10292_ (
    .a(_04477_),
    .b(_00499_),
    .c(_04478_),
    .y(_04479_)
  );
  al_ao21ftf _10293_ (
    .a(g35),
    .b(\DFF_947.Q ),
    .c(_04479_),
    .y(\DFF_590.D )
  );
  al_ao21 _10294_ (
    .a(\DFF_358.Q ),
    .b(_00603_),
    .c(\DFF_63.Q ),
    .y(_04480_)
  );
  al_nand3ftt _10295_ (
    .a(_04256_),
    .b(_04480_),
    .c(_02228_),
    .y(_04481_)
  );
  al_ao21ftf _10296_ (
    .a(g35),
    .b(\DFF_358.Q ),
    .c(_04481_),
    .y(\DFF_63.D )
  );
  al_ao21 _10297_ (
    .a(\DFF_1275.Q ),
    .b(_02533_),
    .c(\DFF_1008.Q ),
    .y(_04482_)
  );
  al_and3 _10298_ (
    .a(_02535_),
    .b(_02534_),
    .c(_04482_),
    .y(\DFF_1008.D )
  );
  al_mux2l _10299_ (
    .a(\DFF_330.Q ),
    .b(\DFF_282.Q ),
    .s(_01193_),
    .y(_04483_)
  );
  al_mux2h _10300_ (
    .a(\DFF_247.Q ),
    .b(_04483_),
    .s(g35),
    .y(\DFF_330.D )
  );
  al_and2ft _10301_ (
    .a(g35),
    .b(\DFF_1028.Q ),
    .y(_04484_)
  );
  al_nand3 _10302_ (
    .a(_00817_),
    .b(_00563_),
    .c(_00815_),
    .y(_04485_)
  );
  al_oa21ftf _10303_ (
    .a(_00560_),
    .b(_00563_),
    .c(_00066_),
    .y(_04486_)
  );
  al_ao21 _10304_ (
    .a(_04486_),
    .b(_04485_),
    .c(_04484_),
    .y(\DFF_148.D )
  );
  al_mux2l _10305_ (
    .a(\DFF_1188.Q ),
    .b(\DFF_251.Q ),
    .s(\DFF_139.Q ),
    .y(_04487_)
  );
  al_aoi21 _10306_ (
    .a(\DFF_118.Q ),
    .b(_04487_),
    .c(\DFF_837.Q ),
    .y(_04488_)
  );
  al_oai21 _10307_ (
    .a(\DFF_118.Q ),
    .b(_04487_),
    .c(_04488_),
    .y(_04489_)
  );
  al_ao21ttf _10308_ (
    .a(_04200_),
    .b(_04489_),
    .c(_01663_),
    .y(_04490_)
  );
  al_or2 _10309_ (
    .a(\DFF_837.Q ),
    .b(_01663_),
    .y(_04491_)
  );
  al_and3 _10310_ (
    .a(g35),
    .b(_04490_),
    .c(_04491_),
    .y(\DFF_837.D )
  );
  al_or3fft _10311_ (
    .a(\DFF_446.Q ),
    .b(g35),
    .c(_02019_),
    .y(_04492_)
  );
  al_or2 _10312_ (
    .a(g35),
    .b(\DFF_583.Q ),
    .y(_04493_)
  );
  al_nand3fft _10313_ (
    .a(\DFF_446.Q ),
    .b(_00066_),
    .c(_02019_),
    .y(_04494_)
  );
  al_and3 _10314_ (
    .a(_04493_),
    .b(_04494_),
    .c(_04492_),
    .y(\DFF_446.D )
  );
  al_nand3 _10315_ (
    .a(\DFF_157.Q ),
    .b(g35),
    .c(_00941_),
    .y(_04495_)
  );
  al_mux2l _10316_ (
    .a(_00242_),
    .b(_04495_),
    .s(_02248_),
    .y(_04496_)
  );
  al_ao21ftf _10317_ (
    .a(g35),
    .b(\DFF_328.Q ),
    .c(_04496_),
    .y(\DFF_157.D )
  );
  al_oa21ftf _10318_ (
    .a(_03304_),
    .b(_00576_),
    .c(_00066_),
    .y(_04497_)
  );
  al_ao21ttf _10319_ (
    .a(_00448_),
    .b(_00578_),
    .c(_04497_),
    .y(_04498_)
  );
  al_ao21ftf _10320_ (
    .a(g35),
    .b(\DFF_462.Q ),
    .c(_04498_),
    .y(\DFF_1091.D )
  );
  al_ao21ftt _10321_ (
    .a(_00100_),
    .b(_01183_),
    .c(_01190_),
    .y(_04499_)
  );
  al_or3fft _10322_ (
    .a(g35),
    .b(_04499_),
    .c(_02551_),
    .y(_04500_)
  );
  al_ao21ftf _10323_ (
    .a(g35),
    .b(\DFF_162.Q ),
    .c(_04500_),
    .y(\DFF_1090.D )
  );
  al_nand3ftt _10324_ (
    .a(_03064_),
    .b(_00499_),
    .c(_00706_),
    .y(_04501_)
  );
  al_ao21ftt _10325_ (
    .a(_03064_),
    .b(_00706_),
    .c(\DFF_1197.Q ),
    .y(_04502_)
  );
  al_nand3 _10326_ (
    .a(g35),
    .b(_04501_),
    .c(_04502_),
    .y(_04503_)
  );
  al_ao21ftf _10327_ (
    .a(g35),
    .b(\DFF_645.Q ),
    .c(_04503_),
    .y(\DFF_1197.D )
  );
  al_nand3ftt _10328_ (
    .a(\DFF_932.Q ),
    .b(g35),
    .c(_00516_),
    .y(_04504_)
  );
  al_aoi21ftf _10329_ (
    .a(\DFF_323.Q ),
    .b(_00066_),
    .c(_04504_),
    .y(\DFF_932.D )
  );
  al_mux2l _10330_ (
    .a(\DFF_1315.Q ),
    .b(\DFF_1108.Q ),
    .s(_01174_),
    .y(\DFF_1108.D )
  );
  al_ao21 _10331_ (
    .a(_03181_),
    .b(_00550_),
    .c(\DFF_946.Q ),
    .y(_04505_)
  );
  al_and2ft _10332_ (
    .a(g35),
    .b(\DFF_1223.Q ),
    .y(_04506_)
  );
  al_ao21 _10333_ (
    .a(_00552_),
    .b(_04505_),
    .c(_04506_),
    .y(\DFF_946.D )
  );
  al_inv _10334_ (
    .a(\DFF_408.Q ),
    .y(_04507_)
  );
  al_and2ft _10335_ (
    .a(\DFF_171.Q ),
    .b(\DFF_990.Q ),
    .y(_04508_)
  );
  al_nand2ft _10336_ (
    .a(\DFF_990.Q ),
    .b(\DFF_171.Q ),
    .y(_04509_)
  );
  al_nand2ft _10337_ (
    .a(_04508_),
    .b(_04509_),
    .y(_04510_)
  );
  al_and3fft _10338_ (
    .a(_00960_),
    .b(_01696_),
    .c(_04510_),
    .y(_04511_)
  );
  al_ao21 _10339_ (
    .a(g35),
    .b(_04511_),
    .c(_04507_),
    .y(_04512_)
  );
  al_and3 _10340_ (
    .a(_04507_),
    .b(g35),
    .c(_04511_),
    .y(_04513_)
  );
  al_nand2ft _10341_ (
    .a(_04513_),
    .b(_04512_),
    .y(\DFF_937.D )
  );
  al_mux2h _10342_ (
    .a(\DFF_729.Q ),
    .b(_01934_),
    .s(_00365_),
    .y(_04514_)
  );
  al_mux2h _10343_ (
    .a(\DFF_1210.Q ),
    .b(_04514_),
    .s(g35),
    .y(\DFF_729.D )
  );
  al_ao21 _10344_ (
    .a(_01576_),
    .b(_00550_),
    .c(\DFF_1223.Q ),
    .y(_04515_)
  );
  al_and2ft _10345_ (
    .a(g35),
    .b(\DFF_1036.Q ),
    .y(_04516_)
  );
  al_ao21 _10346_ (
    .a(_00552_),
    .b(_04515_),
    .c(_04516_),
    .y(\DFF_1223.D )
  );
  al_mux2l _10347_ (
    .a(\DFF_824.Q ),
    .b(_04317_),
    .s(_04315_),
    .y(_04517_)
  );
  al_mux2h _10348_ (
    .a(\DFF_258.Q ),
    .b(_04517_),
    .s(g35),
    .y(\DFF_824.D )
  );
  al_and2 _10349_ (
    .a(\DFF_1068.Q ),
    .b(g35),
    .y(\DFF_861.D )
  );
  al_nor2 _10350_ (
    .a(_00066_),
    .b(_02775_),
    .y(_04518_)
  );
  al_nand2ft _10351_ (
    .a(\DFF_174.Q ),
    .b(_03179_),
    .y(_04519_)
  );
  al_mux2h _10352_ (
    .a(\DFF_1063.Q ),
    .b(_04519_),
    .s(g35),
    .y(_04520_)
  );
  al_aoi21ftf _10353_ (
    .a(\DFF_103.Q ),
    .b(_04518_),
    .c(_04520_),
    .y(\DFF_103.D )
  );
  al_nand3 _10354_ (
    .a(_00499_),
    .b(_02113_),
    .c(_00705_),
    .y(_04521_)
  );
  al_ao21 _10355_ (
    .a(_00705_),
    .b(_02113_),
    .c(\DFF_9.Q ),
    .y(_04522_)
  );
  al_nand3 _10356_ (
    .a(g35),
    .b(_04522_),
    .c(_04521_),
    .y(_04523_)
  );
  al_ao21ftf _10357_ (
    .a(g35),
    .b(\DFF_640.Q ),
    .c(_04523_),
    .y(\DFF_9.D )
  );
  al_nand2ft _10358_ (
    .a(\DFF_395.Q ),
    .b(_00638_),
    .y(_04524_)
  );
  al_aoi21ttf _10359_ (
    .a(_04524_),
    .b(_01617_),
    .c(_00641_),
    .y(_04525_)
  );
  al_nand3 _10360_ (
    .a(\DFF_820.Q ),
    .b(_00642_),
    .c(_04525_),
    .y(_04526_)
  );
  al_ao21 _10361_ (
    .a(\DFF_820.Q ),
    .b(_00642_),
    .c(_04525_),
    .y(_04527_)
  );
  al_ao21 _10362_ (
    .a(_04526_),
    .b(_04527_),
    .c(_00066_),
    .y(_04528_)
  );
  al_aoi21ftf _10363_ (
    .a(\DFF_505.Q ),
    .b(_00066_),
    .c(_04528_),
    .y(\DFF_820.D )
  );
  al_oai21ftf _10364_ (
    .a(\DFF_376.Q ),
    .b(\DFF_365.Q ),
    .c(\DFF_329.Q ),
    .y(_04529_)
  );
  al_nand3ftt _10365_ (
    .a(\DFF_85.Q ),
    .b(g35),
    .c(_04529_),
    .y(_04530_)
  );
  al_ao21ftf _10366_ (
    .a(g35),
    .b(\DFF_365.Q ),
    .c(_04530_),
    .y(\DFF_329.D )
  );
  al_and2ft _10367_ (
    .a(g35),
    .b(\DFF_1170.Q ),
    .y(_04531_)
  );
  al_nor2ft _10368_ (
    .a(_01448_),
    .b(_01451_),
    .y(_04532_)
  );
  al_ao21ftf _10369_ (
    .a(_01445_),
    .b(_01455_),
    .c(_04532_),
    .y(_04533_)
  );
  al_oa21ftf _10370_ (
    .a(\DFF_140.Q ),
    .b(_04532_),
    .c(_00066_),
    .y(_04534_)
  );
  al_ao21 _10371_ (
    .a(_04533_),
    .b(_04534_),
    .c(_04531_),
    .y(\DFF_140.D )
  );
  al_or3fft _10372_ (
    .a(_00324_),
    .b(_01150_),
    .c(_01153_),
    .y(_04535_)
  );
  al_ao21 _10373_ (
    .a(_00324_),
    .b(_01150_),
    .c(\DFF_809.Q ),
    .y(_04536_)
  );
  al_nand3 _10374_ (
    .a(g35),
    .b(_04536_),
    .c(_04535_),
    .y(_04537_)
  );
  al_ao21ftf _10375_ (
    .a(g35),
    .b(\DFF_924.Q ),
    .c(_04537_),
    .y(\DFF_809.D )
  );
  al_or3fft _10376_ (
    .a(_00364_),
    .b(_01832_),
    .c(_00851_),
    .y(_04538_)
  );
  al_nand3fft _10377_ (
    .a(\DFF_434.Q ),
    .b(_00066_),
    .c(_04538_),
    .y(_04539_)
  );
  al_ao21ftf _10378_ (
    .a(g35),
    .b(\DFF_1204.Q ),
    .c(_04539_),
    .y(\DFF_685.D )
  );
  al_nand2 _10379_ (
    .a(\DFF_1075.Q ),
    .b(\DFF_882.Q ),
    .y(_04540_)
  );
  al_nor2 _10380_ (
    .a(\DFF_1075.Q ),
    .b(\DFF_882.Q ),
    .y(_04541_)
  );
  al_nand2ft _10381_ (
    .a(_04541_),
    .b(_04540_),
    .y(_04542_)
  );
  al_mux2l _10382_ (
    .a(\DFF_1163.Q ),
    .b(_04542_),
    .s(_00547_),
    .y(_04543_)
  );
  al_mux2h _10383_ (
    .a(\DFF_882.Q ),
    .b(_04543_),
    .s(g35),
    .y(\DFF_1163.D )
  );
  al_mux2l _10384_ (
    .a(g6744),
    .b(\DFF_760.Q ),
    .s(g35),
    .y(\DFF_48.D )
  );
  al_or2 _10385_ (
    .a(_00514_),
    .b(_00526_),
    .y(_04544_)
  );
  al_and3 _10386_ (
    .a(_00513_),
    .b(_02806_),
    .c(_00526_),
    .y(_04545_)
  );
  al_nand2 _10387_ (
    .a(_04545_),
    .b(_02650_),
    .y(_04546_)
  );
  al_aoi21 _10388_ (
    .a(_04544_),
    .b(_04546_),
    .c(_00066_),
    .y(\DFF_209.D )
  );
  al_mux2l _10389_ (
    .a(\DFF_855.Q ),
    .b(\DFF_721.Q ),
    .s(g35),
    .y(\DFF_855.D )
  );
  al_or3ftt _10390_ (
    .a(g44),
    .b(\DFF_349.Q ),
    .c(\DFF_852.Q ),
    .y(_04547_)
  );
  al_mux2h _10391_ (
    .a(\DFF_899.Q ),
    .b(_04547_),
    .s(g35),
    .y(\DFF_852.D )
  );
  al_nand2ft _10392_ (
    .a(\DFF_1014.Q ),
    .b(g35),
    .y(_04548_)
  );
  al_ao21ftf _10393_ (
    .a(g35),
    .b(\DFF_532.Q ),
    .c(_04548_),
    .y(\DFF_686.D )
  );
  al_ao21ftf _10394_ (
    .a(_00940_),
    .b(_00954_),
    .c(_03206_),
    .y(_04549_)
  );
  al_nand3 _10395_ (
    .a(_01175_),
    .b(_03207_),
    .c(_04549_),
    .y(_04550_)
  );
  al_ao21ftf _10396_ (
    .a(g35),
    .b(\DFF_661.Q ),
    .c(_04550_),
    .y(\DFF_21.D )
  );
  al_inv _10397_ (
    .a(\DFF_334.Q ),
    .y(_04551_)
  );
  al_and3fft _10398_ (
    .a(\DFF_327.Q ),
    .b(_02533_),
    .c(_04551_),
    .y(_04552_)
  );
  al_oa21ttf _10399_ (
    .a(_04552_),
    .b(_04511_),
    .c(_00066_),
    .y(_04553_)
  );
  al_ao21ttf _10400_ (
    .a(_04511_),
    .b(_04552_),
    .c(_04553_),
    .y(_04554_)
  );
  al_ao21ftf _10401_ (
    .a(g35),
    .b(\DFF_67.Q ),
    .c(_04554_),
    .y(\DFF_60.D )
  );
  al_and3 _10402_ (
    .a(\DFF_215.Q ),
    .b(\DFF_1190.Q ),
    .c(\DFF_73.Q ),
    .y(_04555_)
  );
  al_or2ft _10403_ (
    .a(\DFF_210.Q ),
    .b(_04555_),
    .y(_04556_)
  );
  al_nand2ft _10404_ (
    .a(\DFF_210.Q ),
    .b(_04555_),
    .y(_04557_)
  );
  al_nand3 _10405_ (
    .a(g35),
    .b(_04557_),
    .c(_04556_),
    .y(_04558_)
  );
  al_aoi21ftf _10406_ (
    .a(\DFF_215.Q ),
    .b(_00066_),
    .c(_04558_),
    .y(\DFF_210.D )
  );
  al_mux2l _10407_ (
    .a(\DFF_1005.Q ),
    .b(\DFF_838.Q ),
    .s(g35),
    .y(\DFF_86.D )
  );
  al_oai21ftf _10408_ (
    .a(g35),
    .b(_03179_),
    .c(\DFF_705.Q ),
    .y(_04559_)
  );
  al_aoi21ftf _10409_ (
    .a(\DFF_174.Q ),
    .b(_04518_),
    .c(_04559_),
    .y(\DFF_174.D )
  );
  al_oa21ftt _10410_ (
    .a(g35),
    .b(_00745_),
    .c(\DFF_107.Q ),
    .y(\DFF_699.D )
  );
  al_nand3 _10411_ (
    .a(\DFF_1281.Q ),
    .b(g35),
    .c(_02440_),
    .y(_04560_)
  );
  al_and3ftt _10412_ (
    .a(_01063_),
    .b(\DFF_1069.Q ),
    .c(_04560_),
    .y(_04561_)
  );
  al_ao21ftt _10413_ (
    .a(_01063_),
    .b(\DFF_1069.Q ),
    .c(_04560_),
    .y(_04562_)
  );
  al_nand2ft _10414_ (
    .a(_04561_),
    .b(_04562_),
    .y(\DFF_1281.D )
  );
  al_aoi21ftf _10415_ (
    .a(\DFF_1299.Q ),
    .b(_00392_),
    .c(\DFF_436.Q ),
    .y(g34839)
  );
  al_nand3 _10416_ (
    .a(_00210_),
    .b(_00201_),
    .c(_00197_),
    .y(\DFF_206.D )
  );
  al_buf _10417_ (
    .a(\DFF_1305.Q ),
    .y(\DFF_530.D )
  );
  al_buf _10418_ (
    .a(\DFF_126.Q ),
    .y(\DFF_448.D )
  );
  al_buf _10419_ (
    .a(\DFF_615.Q ),
    .y(\DFF_184.D )
  );
  al_buf _10420_ (
    .a(\DFF_934.Q ),
    .y(\DFF_961.D )
  );
  al_nand3 _10421_ (
    .a(_00116_),
    .b(_00106_),
    .c(_00099_),
    .y(\DFF_514.D )
  );
  al_nand2 _10422_ (
    .a(_00180_),
    .b(_00164_),
    .y(\DFF_1322.D )
  );
  al_nand3 _10423_ (
    .a(_00258_),
    .b(_00249_),
    .c(_00266_),
    .y(\DFF_150.D )
  );
  al_nand2 _10424_ (
    .a(_00302_),
    .b(_00304_),
    .y(\DFF_621.D )
  );
  al_buf _10425_ (
    .a(\DFF_908.Q ),
    .y(\DFF_1099.D )
  );
  al_nand2 _10426_ (
    .a(_00238_),
    .b(_00223_),
    .y(\DFF_420.D )
  );
  al_nand3fft _10427_ (
    .a(_00130_),
    .b(_00142_),
    .c(_00152_),
    .y(\DFF_1012.D )
  );
  al_buf _10428_ (
    .a(\DFF_1329.Q ),
    .y(\DFF_1149.D )
  );
  al_buf _10429_ (
    .a(\DFF_527.Q ),
    .y(\DFF_434.D )
  );
  al_and2 _10430_ (
    .a(g35),
    .b(g125),
    .y(\DFF_527.D )
  );
  al_and2 _10431_ (
    .a(g113),
    .b(g35),
    .y(\DFF_672.D )
  );
  al_nand2 _10432_ (
    .a(_00276_),
    .b(_00295_),
    .y(\DFF_829.D )
  );
  al_buf _10433_ (
    .a(\DFF_1411.Q ),
    .y(g12832)
  );
  al_nand3 _10434_ (
    .a(_00070_),
    .b(_00092_),
    .c(_00053_),
    .y(\DFF_477.D )
  );
  al_dffl _10435_ (
    .clk(CK),
    .d(\DFF_0.D ),
    .q(\DFF_0.Q )
  );
  al_dffl _10436_ (
    .clk(CK),
    .d(\DFF_1.D ),
    .q(\DFF_1.Q )
  );
  al_dffl _10437_ (
    .clk(CK),
    .d(\DFF_2.D ),
    .q(\DFF_2.Q )
  );
  al_dffl _10438_ (
    .clk(CK),
    .d(\DFF_3.D ),
    .q(\DFF_3.Q )
  );
  al_dffl _10439_ (
    .clk(CK),
    .d(\DFF_4.D ),
    .q(\DFF_4.Q )
  );
  al_dffl _10440_ (
    .clk(CK),
    .d(\DFF_5.D ),
    .q(\DFF_5.Q )
  );
  al_dffl _10441_ (
    .clk(CK),
    .d(\DFF_6.D ),
    .q(\DFF_6.Q )
  );
  al_dffl _10442_ (
    .clk(CK),
    .d(\DFF_752.D ),
    .q(\DFF_752.Q )
  );
  al_dffl _10443_ (
    .clk(CK),
    .d(\DFF_752.Q ),
    .q(\DFF_109.Q )
  );
  al_dffl _10444_ (
    .clk(CK),
    .d(\DFF_109.Q ),
    .q(\DFF_7.Q )
  );
  al_dffl _10445_ (
    .clk(CK),
    .d(\DFF_8.D ),
    .q(\DFF_8.Q )
  );
  al_dffl _10446_ (
    .clk(CK),
    .d(\DFF_9.D ),
    .q(\DFF_9.Q )
  );
  al_dffl _10447_ (
    .clk(CK),
    .d(\DFF_10.D ),
    .q(\DFF_10.Q )
  );
  al_dffl _10448_ (
    .clk(CK),
    .d(\DFF_11.D ),
    .q(\DFF_11.Q )
  );
  al_dffl _10449_ (
    .clk(CK),
    .d(\DFF_12.D ),
    .q(\DFF_12.Q )
  );
  al_dffl _10450_ (
    .clk(CK),
    .d(\DFF_13.D ),
    .q(\DFF_13.Q )
  );
  al_dffl _10451_ (
    .clk(CK),
    .d(\DFF_14.D ),
    .q(\DFF_14.Q )
  );
  al_dffl _10452_ (
    .clk(CK),
    .d(\DFF_15.D ),
    .q(\DFF_15.Q )
  );
  al_dffl _10453_ (
    .clk(CK),
    .d(\DFF_16.D ),
    .q(\DFF_16.Q )
  );
  al_dffl _10454_ (
    .clk(CK),
    .d(\DFF_17.D ),
    .q(\DFF_17.Q )
  );
  al_dffl _10455_ (
    .clk(CK),
    .d(\DFF_18.D ),
    .q(\DFF_18.Q )
  );
  al_dffl _10456_ (
    .clk(CK),
    .d(\DFF_19.D ),
    .q(\DFF_19.Q )
  );
  al_dffl _10457_ (
    .clk(CK),
    .d(\DFF_20.D ),
    .q(\DFF_20.Q )
  );
  al_dffl _10458_ (
    .clk(CK),
    .d(\DFF_21.D ),
    .q(\DFF_21.Q )
  );
  al_dffl _10459_ (
    .clk(CK),
    .d(\DFF_30.D ),
    .q(\DFF_30.Q )
  );
  al_dffl _10460_ (
    .clk(CK),
    .d(\DFF_30.Q ),
    .q(\DFF_326.Q )
  );
  al_dffl _10461_ (
    .clk(CK),
    .d(\DFF_326.Q ),
    .q(\DFF_797.Q )
  );
  al_dffl _10462_ (
    .clk(CK),
    .d(\DFF_797.Q ),
    .q(\DFF_110.Q )
  );
  al_dffl _10463_ (
    .clk(CK),
    .d(\DFF_110.Q ),
    .q(\DFF_737.Q )
  );
  al_dffl _10464_ (
    .clk(CK),
    .d(\DFF_737.Q ),
    .q(\DFF_1087.Q )
  );
  al_dffl _10465_ (
    .clk(CK),
    .d(\DFF_1087.Q ),
    .q(\DFF_848.Q )
  );
  al_dffl _10466_ (
    .clk(CK),
    .d(\DFF_848.Q ),
    .q(\DFF_1102.Q )
  );
  al_dffl _10467_ (
    .clk(CK),
    .d(\DFF_1102.Q ),
    .q(\DFF_279.Q )
  );
  al_dffl _10468_ (
    .clk(CK),
    .d(\DFF_279.Q ),
    .q(\DFF_22.Q )
  );
  al_dffl _10469_ (
    .clk(CK),
    .d(\DFF_23.D ),
    .q(\DFF_23.Q )
  );
  al_dffl _10470_ (
    .clk(CK),
    .d(\DFF_24.D ),
    .q(\DFF_24.Q )
  );
  al_dffl _10471_ (
    .clk(CK),
    .d(\DFF_25.D ),
    .q(\DFF_25.Q )
  );
  al_dffl _10472_ (
    .clk(CK),
    .d(\DFF_26.D ),
    .q(\DFF_26.Q )
  );
  al_dffl _10473_ (
    .clk(CK),
    .d(\DFF_27.D ),
    .q(\DFF_27.Q )
  );
  al_dffl _10474_ (
    .clk(CK),
    .d(\DFF_28.D ),
    .q(\DFF_28.Q )
  );
  al_dffl _10475_ (
    .clk(CK),
    .d(\DFF_29.D ),
    .q(\DFF_29.Q )
  );
  al_dffl _10476_ (
    .clk(CK),
    .d(\DFF_389.D ),
    .q(\DFF_389.Q )
  );
  al_dffl _10477_ (
    .clk(CK),
    .d(\DFF_389.Q ),
    .q(\DFF_1286.Q )
  );
  al_dffl _10478_ (
    .clk(CK),
    .d(\DFF_1286.Q ),
    .q(\DFF_485.Q )
  );
  al_dffl _10479_ (
    .clk(CK),
    .d(\DFF_485.Q ),
    .q(\DFF_992.Q )
  );
  al_dffl _10480_ (
    .clk(CK),
    .d(\DFF_992.Q ),
    .q(\DFF_885.Q )
  );
  al_dffl _10481_ (
    .clk(CK),
    .d(\DFF_885.Q ),
    .q(\DFF_418.Q )
  );
  al_dffl _10482_ (
    .clk(CK),
    .d(\DFF_418.Q ),
    .q(\DFF_944.Q )
  );
  al_dffl _10483_ (
    .clk(CK),
    .d(\DFF_944.Q ),
    .q(\DFF_1338.Q )
  );
  al_dffl _10484_ (
    .clk(CK),
    .d(\DFF_1338.Q ),
    .q(\DFF_31.Q )
  );
  al_dffl _10485_ (
    .clk(CK),
    .d(\DFF_32.D ),
    .q(\DFF_32.Q )
  );
  al_dffl _10486_ (
    .clk(CK),
    .d(\DFF_33.D ),
    .q(\DFF_33.Q )
  );
  al_dffl _10487_ (
    .clk(CK),
    .d(\DFF_1420.D ),
    .q(\DFF_1420.Q )
  );
  al_dffl _10488_ (
    .clk(CK),
    .d(\DFF_1420.Q ),
    .q(\DFF_468.Q )
  );
  al_dffl _10489_ (
    .clk(CK),
    .d(\DFF_468.Q ),
    .q(\DFF_942.Q )
  );
  al_dffl _10490_ (
    .clk(CK),
    .d(\DFF_942.Q ),
    .q(\DFF_220.Q )
  );
  al_dffl _10491_ (
    .clk(CK),
    .d(\DFF_220.Q ),
    .q(\DFF_81.Q )
  );
  al_dffl _10492_ (
    .clk(CK),
    .d(\DFF_81.Q ),
    .q(\DFF_34.Q )
  );
  al_dffl _10493_ (
    .clk(CK),
    .d(\DFF_35.D ),
    .q(\DFF_35.Q )
  );
  al_dffl _10494_ (
    .clk(CK),
    .d(\DFF_36.D ),
    .q(\DFF_36.Q )
  );
  al_dffl _10495_ (
    .clk(CK),
    .d(\DFF_37.D ),
    .q(\DFF_37.Q )
  );
  al_dffl _10496_ (
    .clk(CK),
    .d(\DFF_1362.Q ),
    .q(\DFF_528.Q )
  );
  al_dffl _10497_ (
    .clk(CK),
    .d(\DFF_528.Q ),
    .q(\DFF_38.Q )
  );
  al_dffl _10498_ (
    .clk(CK),
    .d(\DFF_39.D ),
    .q(\DFF_39.Q )
  );
  al_dffl _10499_ (
    .clk(CK),
    .d(\DFF_40.D ),
    .q(\DFF_40.Q )
  );
  al_dffl _10500_ (
    .clk(CK),
    .d(\DFF_41.D ),
    .q(\DFF_41.Q )
  );
  al_dffl _10501_ (
    .clk(CK),
    .d(\DFF_42.D ),
    .q(\DFF_42.Q )
  );
  al_dffl _10502_ (
    .clk(CK),
    .d(\DFF_43.D ),
    .q(\DFF_43.Q )
  );
  al_dffl _10503_ (
    .clk(CK),
    .d(\DFF_44.D ),
    .q(\DFF_44.Q )
  );
  al_dffl _10504_ (
    .clk(CK),
    .d(\DFF_45.D ),
    .q(\DFF_45.Q )
  );
  al_dffl _10505_ (
    .clk(CK),
    .d(\DFF_46.D ),
    .q(\DFF_46.Q )
  );
  al_dffl _10506_ (
    .clk(CK),
    .d(\DFF_47.D ),
    .q(\DFF_47.Q )
  );
  al_dffl _10507_ (
    .clk(CK),
    .d(\DFF_48.D ),
    .q(\DFF_48.Q )
  );
  al_dffl _10508_ (
    .clk(CK),
    .d(\DFF_49.D ),
    .q(\DFF_49.Q )
  );
  al_dffl _10509_ (
    .clk(CK),
    .d(\DFF_50.D ),
    .q(\DFF_50.Q )
  );
  al_dffl _10510_ (
    .clk(CK),
    .d(\DFF_51.D ),
    .q(\DFF_51.Q )
  );
  al_dffl _10511_ (
    .clk(CK),
    .d(\DFF_52.D ),
    .q(\DFF_52.Q )
  );
  al_dffl _10512_ (
    .clk(CK),
    .d(\DFF_554.D ),
    .q(\DFF_554.Q )
  );
  al_dffl _10513_ (
    .clk(CK),
    .d(\DFF_554.Q ),
    .q(\DFF_188.Q )
  );
  al_dffl _10514_ (
    .clk(CK),
    .d(\DFF_188.Q ),
    .q(\DFF_474.Q )
  );
  al_dffl _10515_ (
    .clk(CK),
    .d(\DFF_474.Q ),
    .q(\DFF_315.Q )
  );
  al_dffl _10516_ (
    .clk(CK),
    .d(\DFF_315.Q ),
    .q(\DFF_123.Q )
  );
  al_dffl _10517_ (
    .clk(CK),
    .d(\DFF_123.Q ),
    .q(\DFF_1119.Q )
  );
  al_dffl _10518_ (
    .clk(CK),
    .d(\DFF_1119.Q ),
    .q(\DFF_970.Q )
  );
  al_dffl _10519_ (
    .clk(CK),
    .d(\DFF_970.Q ),
    .q(\DFF_905.Q )
  );
  al_dffl _10520_ (
    .clk(CK),
    .d(\DFF_905.Q ),
    .q(\DFF_898.Q )
  );
  al_dffl _10521_ (
    .clk(CK),
    .d(\DFF_898.Q ),
    .q(\DFF_53.Q )
  );
  al_dffl _10522_ (
    .clk(CK),
    .d(\DFF_54.D ),
    .q(\DFF_54.Q )
  );
  al_dffl _10523_ (
    .clk(CK),
    .d(\DFF_55.D ),
    .q(\DFF_55.Q )
  );
  al_dffl _10524_ (
    .clk(CK),
    .d(\DFF_56.D ),
    .q(\DFF_56.Q )
  );
  al_dffl _10525_ (
    .clk(CK),
    .d(\DFF_57.D ),
    .q(\DFF_57.Q )
  );
  al_dffl _10526_ (
    .clk(CK),
    .d(\DFF_58.D ),
    .q(\DFF_58.Q )
  );
  al_dffl _10527_ (
    .clk(CK),
    .d(\DFF_59.D ),
    .q(\DFF_59.Q )
  );
  al_dffl _10528_ (
    .clk(CK),
    .d(\DFF_60.D ),
    .q(\DFF_60.Q )
  );
  al_dffl _10529_ (
    .clk(CK),
    .d(\DFF_61.D ),
    .q(\DFF_61.Q )
  );
  al_dffl _10530_ (
    .clk(CK),
    .d(\DFF_62.D ),
    .q(\DFF_62.Q )
  );
  al_dffl _10531_ (
    .clk(CK),
    .d(\DFF_63.D ),
    .q(\DFF_63.Q )
  );
  al_dffl _10532_ (
    .clk(CK),
    .d(\DFF_64.D ),
    .q(\DFF_64.Q )
  );
  al_dffl _10533_ (
    .clk(CK),
    .d(\DFF_65.D ),
    .q(\DFF_65.Q )
  );
  al_dffl _10534_ (
    .clk(CK),
    .d(\DFF_66.D ),
    .q(\DFF_66.Q )
  );
  al_dffl _10535_ (
    .clk(CK),
    .d(\DFF_67.D ),
    .q(\DFF_67.Q )
  );
  al_dffl _10536_ (
    .clk(CK),
    .d(\DFF_68.D ),
    .q(\DFF_68.Q )
  );
  al_dffl _10537_ (
    .clk(CK),
    .d(\DFF_69.D ),
    .q(\DFF_69.Q )
  );
  al_dffl _10538_ (
    .clk(CK),
    .d(\DFF_70.D ),
    .q(\DFF_70.Q )
  );
  al_dffl _10539_ (
    .clk(CK),
    .d(\DFF_71.D ),
    .q(\DFF_71.Q )
  );
  al_dffl _10540_ (
    .clk(CK),
    .d(\DFF_72.D ),
    .q(\DFF_72.Q )
  );
  al_dffl _10541_ (
    .clk(CK),
    .d(\DFF_73.D ),
    .q(\DFF_73.Q )
  );
  al_dffl _10542_ (
    .clk(CK),
    .d(\DFF_74.D ),
    .q(\DFF_74.Q )
  );
  al_dffl _10543_ (
    .clk(CK),
    .d(\DFF_75.D ),
    .q(\DFF_75.Q )
  );
  al_dffl _10544_ (
    .clk(CK),
    .d(\DFF_819.D ),
    .q(\DFF_819.Q )
  );
  al_dffl _10545_ (
    .clk(CK),
    .d(\DFF_819.Q ),
    .q(\DFF_529.Q )
  );
  al_dffl _10546_ (
    .clk(CK),
    .d(\DFF_529.Q ),
    .q(\DFF_1038.Q )
  );
  al_dffl _10547_ (
    .clk(CK),
    .d(\DFF_1038.Q ),
    .q(\DFF_1293.Q )
  );
  al_dffl _10548_ (
    .clk(CK),
    .d(\DFF_1293.Q ),
    .q(\DFF_1354.Q )
  );
  al_dffl _10549_ (
    .clk(CK),
    .d(\DFF_1354.Q ),
    .q(\DFF_1155.Q )
  );
  al_dffl _10550_ (
    .clk(CK),
    .d(\DFF_1155.Q ),
    .q(\DFF_856.Q )
  );
  al_dffl _10551_ (
    .clk(CK),
    .d(\DFF_856.Q ),
    .q(\DFF_76.Q )
  );
  al_dffl _10552_ (
    .clk(CK),
    .d(\DFF_77.D ),
    .q(\DFF_77.Q )
  );
  al_dffl _10553_ (
    .clk(CK),
    .d(\DFF_78.D ),
    .q(\DFF_78.Q )
  );
  al_dffl _10554_ (
    .clk(CK),
    .d(\DFF_79.D ),
    .q(\DFF_79.Q )
  );
  al_dffl _10555_ (
    .clk(CK),
    .d(\DFF_80.D ),
    .q(\DFF_80.Q )
  );
  al_dffl _10556_ (
    .clk(CK),
    .d(\DFF_82.D ),
    .q(\DFF_82.Q )
  );
  al_dffl _10557_ (
    .clk(CK),
    .d(\DFF_83.D ),
    .q(\DFF_83.Q )
  );
  al_dffl _10558_ (
    .clk(CK),
    .d(\DFF_84.D ),
    .q(\DFF_84.Q )
  );
  al_dffl _10559_ (
    .clk(CK),
    .d(\DFF_85.D ),
    .q(\DFF_85.Q )
  );
  al_dffl _10560_ (
    .clk(CK),
    .d(\DFF_86.D ),
    .q(\DFF_86.Q )
  );
  al_dffl _10561_ (
    .clk(CK),
    .d(\DFF_87.D ),
    .q(\DFF_87.Q )
  );
  al_dffl _10562_ (
    .clk(CK),
    .d(\DFF_88.D ),
    .q(\DFF_88.Q )
  );
  al_dffl _10563_ (
    .clk(CK),
    .d(\DFF_89.D ),
    .q(\DFF_89.Q )
  );
  al_dffl _10564_ (
    .clk(CK),
    .d(\DFF_90.D ),
    .q(\DFF_90.Q )
  );
  al_dffl _10565_ (
    .clk(CK),
    .d(\DFF_91.D ),
    .q(\DFF_91.Q )
  );
  al_dffl _10566_ (
    .clk(CK),
    .d(\DFF_92.D ),
    .q(\DFF_92.Q )
  );
  al_dffl _10567_ (
    .clk(CK),
    .d(\DFF_93.D ),
    .q(\DFF_93.Q )
  );
  al_dffl _10568_ (
    .clk(CK),
    .d(\DFF_94.D ),
    .q(\DFF_94.Q )
  );
  al_dffl _10569_ (
    .clk(CK),
    .d(\DFF_95.D ),
    .q(\DFF_95.Q )
  );
  al_dffl _10570_ (
    .clk(CK),
    .d(\DFF_96.D ),
    .q(\DFF_96.Q )
  );
  al_dffl _10571_ (
    .clk(CK),
    .d(\DFF_97.D ),
    .q(\DFF_97.Q )
  );
  al_dffl _10572_ (
    .clk(CK),
    .d(\DFF_98.D ),
    .q(\DFF_98.Q )
  );
  al_dffl _10573_ (
    .clk(CK),
    .d(\DFF_99.D ),
    .q(\DFF_99.Q )
  );
  al_dffl _10574_ (
    .clk(CK),
    .d(\DFF_100.D ),
    .q(\DFF_100.Q )
  );
  al_dffl _10575_ (
    .clk(CK),
    .d(\DFF_46.Q ),
    .q(\DFF_1335.Q )
  );
  al_dffl _10576_ (
    .clk(CK),
    .d(\DFF_1335.Q ),
    .q(\DFF_117.Q )
  );
  al_dffl _10577_ (
    .clk(CK),
    .d(\DFF_117.Q ),
    .q(\DFF_263.Q )
  );
  al_dffl _10578_ (
    .clk(CK),
    .d(\DFF_263.Q ),
    .q(\DFF_101.Q )
  );
  al_dffl _10579_ (
    .clk(CK),
    .d(\DFF_102.D ),
    .q(\DFF_102.Q )
  );
  al_dffl _10580_ (
    .clk(CK),
    .d(\DFF_103.D ),
    .q(\DFF_103.Q )
  );
  al_dffl _10581_ (
    .clk(CK),
    .d(\DFF_104.D ),
    .q(\DFF_104.Q )
  );
  al_dffl _10582_ (
    .clk(CK),
    .d(\DFF_105.D ),
    .q(\DFF_105.Q )
  );
  al_dffl _10583_ (
    .clk(CK),
    .d(\DFF_106.D ),
    .q(\DFF_106.Q )
  );
  al_dffl _10584_ (
    .clk(CK),
    .d(\DFF_107.D ),
    .q(\DFF_107.Q )
  );
  al_dffl _10585_ (
    .clk(CK),
    .d(\DFF_108.D ),
    .q(\DFF_108.Q )
  );
  al_dffl _10586_ (
    .clk(CK),
    .d(\DFF_111.D ),
    .q(\DFF_111.Q )
  );
  al_dffl _10587_ (
    .clk(CK),
    .d(\DFF_112.D ),
    .q(\DFF_112.Q )
  );
  al_dffl _10588_ (
    .clk(CK),
    .d(\DFF_113.D ),
    .q(\DFF_113.Q )
  );
  al_dffl _10589_ (
    .clk(CK),
    .d(\DFF_114.D ),
    .q(\DFF_114.Q )
  );
  al_dffl _10590_ (
    .clk(CK),
    .d(\DFF_115.D ),
    .q(\DFF_115.Q )
  );
  al_dffl _10591_ (
    .clk(CK),
    .d(\DFF_116.D ),
    .q(\DFF_116.Q )
  );
  al_dffl _10592_ (
    .clk(CK),
    .d(\DFF_118.D ),
    .q(\DFF_118.Q )
  );
  al_dffl _10593_ (
    .clk(CK),
    .d(\DFF_119.D ),
    .q(\DFF_119.Q )
  );
  al_dffl _10594_ (
    .clk(CK),
    .d(\DFF_120.D ),
    .q(\DFF_120.Q )
  );
  al_dffl _10595_ (
    .clk(CK),
    .d(\DFF_121.D ),
    .q(\DFF_121.Q )
  );
  al_dffl _10596_ (
    .clk(CK),
    .d(\DFF_122.D ),
    .q(\DFF_122.Q )
  );
  al_dffl _10597_ (
    .clk(CK),
    .d(\DFF_124.D ),
    .q(\DFF_124.Q )
  );
  al_dffl _10598_ (
    .clk(CK),
    .d(\DFF_125.D ),
    .q(\DFF_125.Q )
  );
  al_dffl _10599_ (
    .clk(CK),
    .d(\DFF_126.D ),
    .q(\DFF_126.Q )
  );
  al_dffl _10600_ (
    .clk(CK),
    .d(\DFF_127.D ),
    .q(\DFF_127.Q )
  );
  al_dffl _10601_ (
    .clk(CK),
    .d(\DFF_128.D ),
    .q(\DFF_128.Q )
  );
  al_dffl _10602_ (
    .clk(CK),
    .d(\DFF_129.D ),
    .q(\DFF_129.Q )
  );
  al_dffl _10603_ (
    .clk(CK),
    .d(\DFF_130.D ),
    .q(\DFF_130.Q )
  );
  al_dffl _10604_ (
    .clk(CK),
    .d(\DFF_131.D ),
    .q(\DFF_131.Q )
  );
  al_dffl _10605_ (
    .clk(CK),
    .d(\DFF_132.D ),
    .q(\DFF_132.Q )
  );
  al_dffl _10606_ (
    .clk(CK),
    .d(\DFF_133.D ),
    .q(\DFF_133.Q )
  );
  al_dffl _10607_ (
    .clk(CK),
    .d(\DFF_134.D ),
    .q(\DFF_134.Q )
  );
  al_dffl _10608_ (
    .clk(CK),
    .d(\DFF_135.D ),
    .q(\DFF_135.Q )
  );
  al_dffl _10609_ (
    .clk(CK),
    .d(\DFF_136.D ),
    .q(\DFF_136.Q )
  );
  al_dffl _10610_ (
    .clk(CK),
    .d(\DFF_137.D ),
    .q(\DFF_137.Q )
  );
  al_dffl _10611_ (
    .clk(CK),
    .d(\DFF_138.D ),
    .q(\DFF_138.Q )
  );
  al_dffl _10612_ (
    .clk(CK),
    .d(\DFF_139.D ),
    .q(\DFF_139.Q )
  );
  al_dffl _10613_ (
    .clk(CK),
    .d(\DFF_140.D ),
    .q(\DFF_140.Q )
  );
  al_dffl _10614_ (
    .clk(CK),
    .d(\DFF_141.D ),
    .q(\DFF_141.Q )
  );
  al_dffl _10615_ (
    .clk(CK),
    .d(\DFF_142.D ),
    .q(\DFF_142.Q )
  );
  al_dffl _10616_ (
    .clk(CK),
    .d(\DFF_143.D ),
    .q(\DFF_143.Q )
  );
  al_dffl _10617_ (
    .clk(CK),
    .d(\DFF_144.D ),
    .q(\DFF_144.Q )
  );
  al_dffl _10618_ (
    .clk(CK),
    .d(\DFF_145.D ),
    .q(\DFF_145.Q )
  );
  al_dffl _10619_ (
    .clk(CK),
    .d(\DFF_422.D ),
    .q(\DFF_422.Q )
  );
  al_dffl _10620_ (
    .clk(CK),
    .d(\DFF_422.Q ),
    .q(\DFF_146.Q )
  );
  al_dffl _10621_ (
    .clk(CK),
    .d(\DFF_147.D ),
    .q(\DFF_147.Q )
  );
  al_dffl _10622_ (
    .clk(CK),
    .d(\DFF_148.D ),
    .q(\DFF_148.Q )
  );
  al_dffl _10623_ (
    .clk(CK),
    .d(\DFF_149.D ),
    .q(\DFF_149.Q )
  );
  al_dffl _10624_ (
    .clk(CK),
    .d(\DFF_150.D ),
    .q(\DFF_150.Q )
  );
  al_dffl _10625_ (
    .clk(CK),
    .d(\DFF_151.D ),
    .q(\DFF_151.Q )
  );
  al_dffl _10626_ (
    .clk(CK),
    .d(\DFF_585.D ),
    .q(\DFF_585.Q )
  );
  al_dffl _10627_ (
    .clk(CK),
    .d(\DFF_585.Q ),
    .q(\DFF_561.Q )
  );
  al_dffl _10628_ (
    .clk(CK),
    .d(\DFF_561.Q ),
    .q(\DFF_1106.Q )
  );
  al_dffl _10629_ (
    .clk(CK),
    .d(\DFF_1106.Q ),
    .q(\DFF_152.Q )
  );
  al_dffl _10630_ (
    .clk(CK),
    .d(\DFF_153.D ),
    .q(\DFF_153.Q )
  );
  al_dffl _10631_ (
    .clk(CK),
    .d(\DFF_154.D ),
    .q(\DFF_154.Q )
  );
  al_dffl _10632_ (
    .clk(CK),
    .d(\DFF_155.D ),
    .q(\DFF_155.Q )
  );
  al_dffl _10633_ (
    .clk(CK),
    .d(\DFF_156.D ),
    .q(\DFF_156.Q )
  );
  al_dffl _10634_ (
    .clk(CK),
    .d(\DFF_157.D ),
    .q(\DFF_157.Q )
  );
  al_dffl _10635_ (
    .clk(CK),
    .d(\DFF_158.D ),
    .q(\DFF_158.Q )
  );
  al_dffl _10636_ (
    .clk(CK),
    .d(\DFF_159.D ),
    .q(\DFF_159.Q )
  );
  al_dffl _10637_ (
    .clk(CK),
    .d(\DFF_160.D ),
    .q(\DFF_160.Q )
  );
  al_dffl _10638_ (
    .clk(CK),
    .d(\DFF_161.D ),
    .q(\DFF_161.Q )
  );
  al_dffl _10639_ (
    .clk(CK),
    .d(\DFF_162.D ),
    .q(\DFF_162.Q )
  );
  al_dffl _10640_ (
    .clk(CK),
    .d(\DFF_1158.D ),
    .q(\DFF_1158.Q )
  );
  al_dffl _10641_ (
    .clk(CK),
    .d(\DFF_1158.Q ),
    .q(\DFF_806.Q )
  );
  al_dffl _10642_ (
    .clk(CK),
    .d(\DFF_806.Q ),
    .q(\DFF_1196.Q )
  );
  al_dffl _10643_ (
    .clk(CK),
    .d(\DFF_1196.Q ),
    .q(\DFF_1248.Q )
  );
  al_dffl _10644_ (
    .clk(CK),
    .d(\DFF_1248.Q ),
    .q(\DFF_1185.Q )
  );
  al_dffl _10645_ (
    .clk(CK),
    .d(\DFF_1185.Q ),
    .q(\DFF_163.Q )
  );
  al_dffl _10646_ (
    .clk(CK),
    .d(\DFF_164.D ),
    .q(\DFF_164.Q )
  );
  al_dffl _10647_ (
    .clk(CK),
    .d(\DFF_165.D ),
    .q(\DFF_165.Q )
  );
  al_dffl _10648_ (
    .clk(CK),
    .d(\DFF_317.D ),
    .q(\DFF_317.Q )
  );
  al_dffl _10649_ (
    .clk(CK),
    .d(\DFF_317.Q ),
    .q(\DFF_166.Q )
  );
  al_dffl _10650_ (
    .clk(CK),
    .d(\DFF_167.D ),
    .q(\DFF_167.Q )
  );
  al_dffl _10651_ (
    .clk(CK),
    .d(\DFF_371.D ),
    .q(\DFF_371.Q )
  );
  al_dffl _10652_ (
    .clk(CK),
    .d(\DFF_371.Q ),
    .q(\DFF_168.Q )
  );
  al_dffl _10653_ (
    .clk(CK),
    .d(\DFF_169.D ),
    .q(\DFF_169.Q )
  );
  al_dffl _10654_ (
    .clk(CK),
    .d(\DFF_170.D ),
    .q(\DFF_170.Q )
  );
  al_dffl _10655_ (
    .clk(CK),
    .d(\DFF_1072.D ),
    .q(\DFF_1072.Q )
  );
  al_dffl _10656_ (
    .clk(CK),
    .d(\DFF_1072.Q ),
    .q(\DFF_171.Q )
  );
  al_dffl _10657_ (
    .clk(CK),
    .d(\DFF_172.D ),
    .q(\DFF_172.Q )
  );
  al_dffl _10658_ (
    .clk(CK),
    .d(\DFF_173.D ),
    .q(\DFF_173.Q )
  );
  al_dffl _10659_ (
    .clk(CK),
    .d(\DFF_174.D ),
    .q(\DFF_174.Q )
  );
  al_dffl _10660_ (
    .clk(CK),
    .d(\DFF_175.D ),
    .q(\DFF_175.Q )
  );
  al_dffl _10661_ (
    .clk(CK),
    .d(\DFF_176.D ),
    .q(\DFF_176.Q )
  );
  al_dffl _10662_ (
    .clk(CK),
    .d(\DFF_177.D ),
    .q(\DFF_177.Q )
  );
  al_dffl _10663_ (
    .clk(CK),
    .d(\DFF_178.D ),
    .q(\DFF_178.Q )
  );
  al_dffl _10664_ (
    .clk(CK),
    .d(\DFF_179.D ),
    .q(\DFF_179.Q )
  );
  al_dffl _10665_ (
    .clk(CK),
    .d(\DFF_180.D ),
    .q(\DFF_180.Q )
  );
  al_dffl _10666_ (
    .clk(CK),
    .d(\DFF_1001.D ),
    .q(\DFF_1001.Q )
  );
  al_dffl _10667_ (
    .clk(CK),
    .d(\DFF_1001.Q ),
    .q(\DFF_401.Q )
  );
  al_dffl _10668_ (
    .clk(CK),
    .d(\DFF_401.Q ),
    .q(\DFF_305.Q )
  );
  al_dffl _10669_ (
    .clk(CK),
    .d(\DFF_305.Q ),
    .q(\DFF_181.Q )
  );
  al_dffl _10670_ (
    .clk(CK),
    .d(\DFF_182.D ),
    .q(\DFF_182.Q )
  );
  al_dffl _10671_ (
    .clk(CK),
    .d(\DFF_183.D ),
    .q(\DFF_183.Q )
  );
  al_dffl _10672_ (
    .clk(CK),
    .d(\DFF_184.D ),
    .q(\DFF_184.Q )
  );
  al_dffl _10673_ (
    .clk(CK),
    .d(\DFF_185.D ),
    .q(\DFF_185.Q )
  );
  al_dffl _10674_ (
    .clk(CK),
    .d(\DFF_186.D ),
    .q(\DFF_186.Q )
  );
  al_dffl _10675_ (
    .clk(CK),
    .d(\DFF_187.D ),
    .q(\DFF_187.Q )
  );
  al_dffl _10676_ (
    .clk(CK),
    .d(\DFF_189.D ),
    .q(\DFF_189.Q )
  );
  al_dffl _10677_ (
    .clk(CK),
    .d(\DFF_190.D ),
    .q(\DFF_190.Q )
  );
  al_dffl _10678_ (
    .clk(CK),
    .d(\DFF_191.D ),
    .q(\DFF_191.Q )
  );
  al_dffl _10679_ (
    .clk(CK),
    .d(\DFF_192.D ),
    .q(\DFF_192.Q )
  );
  al_dffl _10680_ (
    .clk(CK),
    .d(\DFF_193.D ),
    .q(\DFF_193.Q )
  );
  al_dffl _10681_ (
    .clk(CK),
    .d(\DFF_194.D ),
    .q(\DFF_194.Q )
  );
  al_dffl _10682_ (
    .clk(CK),
    .d(\DFF_195.D ),
    .q(\DFF_195.Q )
  );
  al_dffl _10683_ (
    .clk(CK),
    .d(\DFF_196.D ),
    .q(\DFF_196.Q )
  );
  al_dffl _10684_ (
    .clk(CK),
    .d(\DFF_197.D ),
    .q(\DFF_197.Q )
  );
  al_dffl _10685_ (
    .clk(CK),
    .d(\DFF_198.D ),
    .q(\DFF_198.Q )
  );
  al_dffl _10686_ (
    .clk(CK),
    .d(\DFF_199.D ),
    .q(\DFF_199.Q )
  );
  al_dffl _10687_ (
    .clk(CK),
    .d(\DFF_200.D ),
    .q(\DFF_200.Q )
  );
  al_dffl _10688_ (
    .clk(CK),
    .d(\DFF_201.D ),
    .q(\DFF_201.Q )
  );
  al_dffl _10689_ (
    .clk(CK),
    .d(\DFF_202.D ),
    .q(\DFF_202.Q )
  );
  al_dffl _10690_ (
    .clk(CK),
    .d(\DFF_203.D ),
    .q(\DFF_203.Q )
  );
  al_dffl _10691_ (
    .clk(CK),
    .d(\DFF_204.D ),
    .q(\DFF_204.Q )
  );
  al_dffl _10692_ (
    .clk(CK),
    .d(\DFF_205.D ),
    .q(\DFF_205.Q )
  );
  al_dffl _10693_ (
    .clk(CK),
    .d(\DFF_206.D ),
    .q(\DFF_206.Q )
  );
  al_dffl _10694_ (
    .clk(CK),
    .d(\DFF_207.D ),
    .q(\DFF_207.Q )
  );
  al_dffl _10695_ (
    .clk(CK),
    .d(\DFF_208.D ),
    .q(\DFF_208.Q )
  );
  al_dffl _10696_ (
    .clk(CK),
    .d(\DFF_209.D ),
    .q(\DFF_209.Q )
  );
  al_dffl _10697_ (
    .clk(CK),
    .d(\DFF_210.D ),
    .q(\DFF_210.Q )
  );
  al_dffl _10698_ (
    .clk(CK),
    .d(\DFF_211.D ),
    .q(\DFF_211.Q )
  );
  al_dffl _10699_ (
    .clk(CK),
    .d(\DFF_212.D ),
    .q(\DFF_212.Q )
  );
  al_dffl _10700_ (
    .clk(CK),
    .d(\DFF_213.D ),
    .q(\DFF_213.Q )
  );
  al_dffl _10701_ (
    .clk(CK),
    .d(\DFF_214.D ),
    .q(\DFF_214.Q )
  );
  al_dffl _10702_ (
    .clk(CK),
    .d(\DFF_215.D ),
    .q(\DFF_215.Q )
  );
  al_dffl _10703_ (
    .clk(CK),
    .d(\DFF_216.D ),
    .q(\DFF_216.Q )
  );
  al_dffl _10704_ (
    .clk(CK),
    .d(\DFF_217.D ),
    .q(\DFF_217.Q )
  );
  al_dffl _10705_ (
    .clk(CK),
    .d(\DFF_218.D ),
    .q(\DFF_218.Q )
  );
  al_dffl _10706_ (
    .clk(CK),
    .d(\DFF_219.D ),
    .q(\DFF_219.Q )
  );
  al_dffl _10707_ (
    .clk(CK),
    .d(\DFF_221.D ),
    .q(\DFF_221.Q )
  );
  al_dffl _10708_ (
    .clk(CK),
    .d(\DFF_222.D ),
    .q(\DFF_222.Q )
  );
  al_dffl _10709_ (
    .clk(CK),
    .d(\DFF_223.D ),
    .q(\DFF_223.Q )
  );
  al_dffl _10710_ (
    .clk(CK),
    .d(\DFF_224.D ),
    .q(\DFF_224.Q )
  );
  al_dffl _10711_ (
    .clk(CK),
    .d(\DFF_225.D ),
    .q(\DFF_225.Q )
  );
  al_dffl _10712_ (
    .clk(CK),
    .d(\DFF_226.D ),
    .q(\DFF_226.Q )
  );
  al_dffl _10713_ (
    .clk(CK),
    .d(\DFF_227.D ),
    .q(\DFF_227.Q )
  );
  al_dffl _10714_ (
    .clk(CK),
    .d(\DFF_228.D ),
    .q(\DFF_228.Q )
  );
  al_dffl _10715_ (
    .clk(CK),
    .d(\DFF_229.D ),
    .q(\DFF_229.Q )
  );
  al_dffl _10716_ (
    .clk(CK),
    .d(\DFF_230.D ),
    .q(\DFF_230.Q )
  );
  al_dffl _10717_ (
    .clk(CK),
    .d(\DFF_231.D ),
    .q(\DFF_231.Q )
  );
  al_dffl _10718_ (
    .clk(CK),
    .d(\DFF_232.D ),
    .q(\DFF_232.Q )
  );
  al_dffl _10719_ (
    .clk(CK),
    .d(\DFF_233.D ),
    .q(\DFF_233.Q )
  );
  al_dffl _10720_ (
    .clk(CK),
    .d(\DFF_234.D ),
    .q(\DFF_234.Q )
  );
  al_dffl _10721_ (
    .clk(CK),
    .d(\DFF_85.Q ),
    .q(\DFF_235.Q )
  );
  al_dffl _10722_ (
    .clk(CK),
    .d(\DFF_236.D ),
    .q(\DFF_236.Q )
  );
  al_dffl _10723_ (
    .clk(CK),
    .d(\DFF_237.D ),
    .q(\DFF_237.Q )
  );
  al_dffl _10724_ (
    .clk(CK),
    .d(\DFF_238.D ),
    .q(\DFF_238.Q )
  );
  al_dffl _10725_ (
    .clk(CK),
    .d(\DFF_239.D ),
    .q(\DFF_239.Q )
  );
  al_dffl _10726_ (
    .clk(CK),
    .d(\DFF_240.D ),
    .q(\DFF_240.Q )
  );
  al_dffl _10727_ (
    .clk(CK),
    .d(\DFF_241.D ),
    .q(\DFF_241.Q )
  );
  al_dffl _10728_ (
    .clk(CK),
    .d(\DFF_242.D ),
    .q(\DFF_242.Q )
  );
  al_dffl _10729_ (
    .clk(CK),
    .d(\DFF_243.D ),
    .q(\DFF_243.Q )
  );
  al_dffl _10730_ (
    .clk(CK),
    .d(\DFF_244.D ),
    .q(\DFF_244.Q )
  );
  al_dffl _10731_ (
    .clk(CK),
    .d(\DFF_245.D ),
    .q(\DFF_245.Q )
  );
  al_dffl _10732_ (
    .clk(CK),
    .d(\DFF_246.D ),
    .q(\DFF_246.Q )
  );
  al_dffl _10733_ (
    .clk(CK),
    .d(\DFF_247.D ),
    .q(\DFF_247.Q )
  );
  al_dffl _10734_ (
    .clk(CK),
    .d(\DFF_248.D ),
    .q(\DFF_248.Q )
  );
  al_dffl _10735_ (
    .clk(CK),
    .d(\DFF_249.D ),
    .q(\DFF_249.Q )
  );
  al_dffl _10736_ (
    .clk(CK),
    .d(\DFF_250.D ),
    .q(\DFF_250.Q )
  );
  al_dffl _10737_ (
    .clk(CK),
    .d(\DFF_251.D ),
    .q(\DFF_251.Q )
  );
  al_dffl _10738_ (
    .clk(CK),
    .d(\DFF_252.D ),
    .q(\DFF_252.Q )
  );
  al_dffl _10739_ (
    .clk(CK),
    .d(\DFF_253.D ),
    .q(\DFF_253.Q )
  );
  al_dffl _10740_ (
    .clk(CK),
    .d(\DFF_254.D ),
    .q(\DFF_254.Q )
  );
  al_dffl _10741_ (
    .clk(CK),
    .d(\DFF_255.D ),
    .q(\DFF_255.Q )
  );
  al_dffl _10742_ (
    .clk(CK),
    .d(\DFF_515.D ),
    .q(\DFF_515.Q )
  );
  al_dffl _10743_ (
    .clk(CK),
    .d(\DFF_515.Q ),
    .q(\DFF_1081.Q )
  );
  al_dffl _10744_ (
    .clk(CK),
    .d(\DFF_1081.Q ),
    .q(\DFF_256.Q )
  );
  al_dffl _10745_ (
    .clk(CK),
    .d(\DFF_257.D ),
    .q(\DFF_257.Q )
  );
  al_dffl _10746_ (
    .clk(CK),
    .d(\DFF_258.D ),
    .q(\DFF_258.Q )
  );
  al_dffl _10747_ (
    .clk(CK),
    .d(\DFF_259.D ),
    .q(\DFF_259.Q )
  );
  al_dffl _10748_ (
    .clk(CK),
    .d(\DFF_260.D ),
    .q(\DFF_260.Q )
  );
  al_dffl _10749_ (
    .clk(CK),
    .d(\DFF_261.D ),
    .q(\DFF_261.Q )
  );
  al_dffl _10750_ (
    .clk(CK),
    .d(\DFF_264.D ),
    .q(\DFF_264.Q )
  );
  al_dffl _10751_ (
    .clk(CK),
    .d(\DFF_265.D ),
    .q(\DFF_265.Q )
  );
  al_dffl _10752_ (
    .clk(CK),
    .d(\DFF_266.D ),
    .q(\DFF_266.Q )
  );
  al_dffl _10753_ (
    .clk(CK),
    .d(\DFF_267.D ),
    .q(\DFF_267.Q )
  );
  al_dffl _10754_ (
    .clk(CK),
    .d(\DFF_268.D ),
    .q(\DFF_268.Q )
  );
  al_dffl _10755_ (
    .clk(CK),
    .d(\DFF_269.D ),
    .q(\DFF_269.Q )
  );
  al_dffl _10756_ (
    .clk(CK),
    .d(\DFF_270.D ),
    .q(\DFF_270.Q )
  );
  al_dffl _10757_ (
    .clk(CK),
    .d(\DFF_271.D ),
    .q(\DFF_271.Q )
  );
  al_dffl _10758_ (
    .clk(CK),
    .d(\DFF_272.D ),
    .q(\DFF_272.Q )
  );
  al_dffl _10759_ (
    .clk(CK),
    .d(\DFF_273.D ),
    .q(\DFF_273.Q )
  );
  al_dffl _10760_ (
    .clk(CK),
    .d(\DFF_274.D ),
    .q(\DFF_274.Q )
  );
  al_dffl _10761_ (
    .clk(CK),
    .d(\DFF_275.D ),
    .q(\DFF_275.Q )
  );
  al_dffl _10762_ (
    .clk(CK),
    .d(\DFF_276.D ),
    .q(\DFF_276.Q )
  );
  al_dffl _10763_ (
    .clk(CK),
    .d(\DFF_277.D ),
    .q(\DFF_277.Q )
  );
  al_dffl _10764_ (
    .clk(CK),
    .d(\DFF_278.D ),
    .q(\DFF_278.Q )
  );
  al_dffl _10765_ (
    .clk(CK),
    .d(\DFF_280.D ),
    .q(\DFF_280.Q )
  );
  al_dffl _10766_ (
    .clk(CK),
    .d(\DFF_165.Q ),
    .q(\DFF_655.Q )
  );
  al_dffl _10767_ (
    .clk(CK),
    .d(\DFF_655.Q ),
    .q(\DFF_927.Q )
  );
  al_dffl _10768_ (
    .clk(CK),
    .d(\DFF_927.Q ),
    .q(\DFF_906.Q )
  );
  al_dffl _10769_ (
    .clk(CK),
    .d(\DFF_906.Q ),
    .q(\DFF_566.Q )
  );
  al_dffl _10770_ (
    .clk(CK),
    .d(\DFF_566.Q ),
    .q(\DFF_616.Q )
  );
  al_dffl _10771_ (
    .clk(CK),
    .d(\DFF_616.Q ),
    .q(\DFF_765.Q )
  );
  al_dffl _10772_ (
    .clk(CK),
    .d(\DFF_765.Q ),
    .q(\DFF_537.Q )
  );
  al_dffl _10773_ (
    .clk(CK),
    .d(\DFF_537.Q ),
    .q(\DFF_360.Q )
  );
  al_dffl _10774_ (
    .clk(CK),
    .d(\DFF_360.Q ),
    .q(\DFF_281.Q )
  );
  al_dffl _10775_ (
    .clk(CK),
    .d(\DFF_282.D ),
    .q(\DFF_282.Q )
  );
  al_dffl _10776_ (
    .clk(CK),
    .d(\DFF_283.D ),
    .q(\DFF_283.Q )
  );
  al_dffl _10777_ (
    .clk(CK),
    .d(\DFF_284.D ),
    .q(\DFF_284.Q )
  );
  al_dffl _10778_ (
    .clk(CK),
    .d(\DFF_285.D ),
    .q(\DFF_285.Q )
  );
  al_dffl _10779_ (
    .clk(CK),
    .d(\DFF_286.D ),
    .q(\DFF_286.Q )
  );
  al_dffl _10780_ (
    .clk(CK),
    .d(\DFF_287.D ),
    .q(\DFF_287.Q )
  );
  al_dffl _10781_ (
    .clk(CK),
    .d(\DFF_288.D ),
    .q(\DFF_288.Q )
  );
  al_dffl _10782_ (
    .clk(CK),
    .d(\DFF_289.D ),
    .q(\DFF_289.Q )
  );
  al_dffl _10783_ (
    .clk(CK),
    .d(\DFF_34.Q ),
    .q(\DFF_873.Q )
  );
  al_dffl _10784_ (
    .clk(CK),
    .d(\DFF_873.Q ),
    .q(\DFF_369.Q )
  );
  al_dffl _10785_ (
    .clk(CK),
    .d(\DFF_369.Q ),
    .q(\DFF_1300.Q )
  );
  al_dffl _10786_ (
    .clk(CK),
    .d(\DFF_1300.Q ),
    .q(\DFF_290.Q )
  );
  al_dffl _10787_ (
    .clk(CK),
    .d(\DFF_291.D ),
    .q(\DFF_291.Q )
  );
  al_dffl _10788_ (
    .clk(CK),
    .d(\DFF_292.D ),
    .q(\DFF_292.Q )
  );
  al_dffl _10789_ (
    .clk(CK),
    .d(\DFF_293.D ),
    .q(\DFF_293.Q )
  );
  al_dffl _10790_ (
    .clk(CK),
    .d(\DFF_294.D ),
    .q(\DFF_294.Q )
  );
  al_dffl _10791_ (
    .clk(CK),
    .d(\DFF_711.D ),
    .q(\DFF_711.Q )
  );
  al_dffl _10792_ (
    .clk(CK),
    .d(\DFF_711.Q ),
    .q(\DFF_643.Q )
  );
  al_dffl _10793_ (
    .clk(CK),
    .d(\DFF_643.Q ),
    .q(\DFF_1122.Q )
  );
  al_dffl _10794_ (
    .clk(CK),
    .d(\DFF_1122.Q ),
    .q(\DFF_295.Q )
  );
  al_dffl _10795_ (
    .clk(CK),
    .d(\DFF_296.D ),
    .q(\DFF_296.Q )
  );
  al_dffl _10796_ (
    .clk(CK),
    .d(\DFF_297.D ),
    .q(\DFF_297.Q )
  );
  al_dffl _10797_ (
    .clk(CK),
    .d(\DFF_298.D ),
    .q(\DFF_298.Q )
  );
  al_dffl _10798_ (
    .clk(CK),
    .d(\DFF_147.Q ),
    .q(\DFF_299.Q )
  );
  al_dffl _10799_ (
    .clk(CK),
    .d(\DFF_300.D ),
    .q(\DFF_300.Q )
  );
  al_dffl _10800_ (
    .clk(CK),
    .d(\DFF_301.D ),
    .q(\DFF_301.Q )
  );
  al_dffl _10801_ (
    .clk(CK),
    .d(\DFF_302.D ),
    .q(\DFF_302.Q )
  );
  al_dffl _10802_ (
    .clk(CK),
    .d(\DFF_303.D ),
    .q(\DFF_303.Q )
  );
  al_dffl _10803_ (
    .clk(CK),
    .d(\DFF_304.D ),
    .q(\DFF_304.Q )
  );
  al_dffl _10804_ (
    .clk(CK),
    .d(\DFF_306.D ),
    .q(\DFF_306.Q )
  );
  al_dffl _10805_ (
    .clk(CK),
    .d(\DFF_307.D ),
    .q(\DFF_307.Q )
  );
  al_dffl _10806_ (
    .clk(CK),
    .d(\DFF_308.D ),
    .q(\DFF_308.Q )
  );
  al_dffl _10807_ (
    .clk(CK),
    .d(\DFF_309.D ),
    .q(\DFF_309.Q )
  );
  al_dffl _10808_ (
    .clk(CK),
    .d(\DFF_310.D ),
    .q(\DFF_310.Q )
  );
  al_dffl _10809_ (
    .clk(CK),
    .d(\DFF_311.D ),
    .q(\DFF_311.Q )
  );
  al_dffl _10810_ (
    .clk(CK),
    .d(\DFF_312.D ),
    .q(\DFF_312.Q )
  );
  al_dffl _10811_ (
    .clk(CK),
    .d(\DFF_313.D ),
    .q(\DFF_313.Q )
  );
  al_dffl _10812_ (
    .clk(CK),
    .d(\DFF_314.D ),
    .q(\DFF_314.Q )
  );
  al_dffl _10813_ (
    .clk(CK),
    .d(\DFF_316.D ),
    .q(\DFF_316.Q )
  );
  al_dffl _10814_ (
    .clk(CK),
    .d(\DFF_318.D ),
    .q(\DFF_318.Q )
  );
  al_dffl _10815_ (
    .clk(CK),
    .d(\DFF_319.D ),
    .q(\DFF_319.Q )
  );
  al_dffl _10816_ (
    .clk(CK),
    .d(\DFF_831.D ),
    .q(\DFF_831.Q )
  );
  al_dffl _10817_ (
    .clk(CK),
    .d(\DFF_831.Q ),
    .q(\DFF_320.Q )
  );
  al_dffl _10818_ (
    .clk(CK),
    .d(\DFF_321.D ),
    .q(\DFF_321.Q )
  );
  al_dffl _10819_ (
    .clk(CK),
    .d(\DFF_322.D ),
    .q(\DFF_322.Q )
  );
  al_dffl _10820_ (
    .clk(CK),
    .d(\DFF_323.D ),
    .q(\DFF_323.Q )
  );
  al_dffl _10821_ (
    .clk(CK),
    .d(\DFF_324.D ),
    .q(\DFF_324.Q )
  );
  al_dffl _10822_ (
    .clk(CK),
    .d(\DFF_739.D ),
    .q(\DFF_739.Q )
  );
  al_dffl _10823_ (
    .clk(CK),
    .d(\DFF_739.Q ),
    .q(\DFF_325.Q )
  );
  al_dffl _10824_ (
    .clk(CK),
    .d(\DFF_937.D ),
    .q(\DFF_937.Q )
  );
  al_dffl _10825_ (
    .clk(CK),
    .d(\DFF_937.Q ),
    .q(\DFF_327.Q )
  );
  al_dffl _10826_ (
    .clk(CK),
    .d(\DFF_328.D ),
    .q(\DFF_328.Q )
  );
  al_dffl _10827_ (
    .clk(CK),
    .d(\DFF_329.D ),
    .q(\DFF_329.Q )
  );
  al_dffl _10828_ (
    .clk(CK),
    .d(\DFF_330.D ),
    .q(\DFF_330.Q )
  );
  al_dffl _10829_ (
    .clk(CK),
    .d(\DFF_331.D ),
    .q(\DFF_331.Q )
  );
  al_dffl _10830_ (
    .clk(CK),
    .d(\DFF_332.D ),
    .q(\DFF_332.Q )
  );
  al_dffl _10831_ (
    .clk(CK),
    .d(\DFF_333.D ),
    .q(\DFF_333.Q )
  );
  al_dffl _10832_ (
    .clk(CK),
    .d(\DFF_60.Q ),
    .q(\DFF_334.Q )
  );
  al_dffl _10833_ (
    .clk(CK),
    .d(\DFF_335.D ),
    .q(\DFF_335.Q )
  );
  al_dffl _10834_ (
    .clk(CK),
    .d(\DFF_336.D ),
    .q(\DFF_336.Q )
  );
  al_dffl _10835_ (
    .clk(CK),
    .d(\DFF_337.D ),
    .q(\DFF_337.Q )
  );
  al_dffl _10836_ (
    .clk(CK),
    .d(\DFF_338.D ),
    .q(\DFF_338.Q )
  );
  al_dffl _10837_ (
    .clk(CK),
    .d(\DFF_339.D ),
    .q(\DFF_339.Q )
  );
  al_dffl _10838_ (
    .clk(CK),
    .d(\DFF_340.D ),
    .q(\DFF_340.Q )
  );
  al_dffl _10839_ (
    .clk(CK),
    .d(\DFF_341.D ),
    .q(\DFF_341.Q )
  );
  al_dffl _10840_ (
    .clk(CK),
    .d(\DFF_342.D ),
    .q(\DFF_342.Q )
  );
  al_dffl _10841_ (
    .clk(CK),
    .d(\DFF_343.D ),
    .q(\DFF_343.Q )
  );
  al_dffl _10842_ (
    .clk(CK),
    .d(\DFF_344.D ),
    .q(\DFF_344.Q )
  );
  al_dffl _10843_ (
    .clk(CK),
    .d(\DFF_345.D ),
    .q(\DFF_345.Q )
  );
  al_dffl _10844_ (
    .clk(CK),
    .d(\DFF_346.D ),
    .q(\DFF_346.Q )
  );
  al_dffl _10845_ (
    .clk(CK),
    .d(\DFF_347.D ),
    .q(\DFF_347.Q )
  );
  al_dffl _10846_ (
    .clk(CK),
    .d(\DFF_348.D ),
    .q(\DFF_348.Q )
  );
  al_dffl _10847_ (
    .clk(CK),
    .d(\DFF_349.D ),
    .q(\DFF_349.Q )
  );
  al_dffl _10848_ (
    .clk(CK),
    .d(\DFF_350.D ),
    .q(\DFF_350.Q )
  );
  al_dffl _10849_ (
    .clk(CK),
    .d(\DFF_351.D ),
    .q(\DFF_351.Q )
  );
  al_dffl _10850_ (
    .clk(CK),
    .d(\DFF_352.D ),
    .q(\DFF_352.Q )
  );
  al_dffl _10851_ (
    .clk(CK),
    .d(\DFF_353.D ),
    .q(\DFF_353.Q )
  );
  al_dffl _10852_ (
    .clk(CK),
    .d(\DFF_354.D ),
    .q(\DFF_354.Q )
  );
  al_dffl _10853_ (
    .clk(CK),
    .d(\DFF_355.D ),
    .q(\DFF_355.Q )
  );
  al_dffl _10854_ (
    .clk(CK),
    .d(\DFF_356.D ),
    .q(\DFF_356.Q )
  );
  al_dffl _10855_ (
    .clk(CK),
    .d(\DFF_357.D ),
    .q(\DFF_357.Q )
  );
  al_dffl _10856_ (
    .clk(CK),
    .d(\DFF_358.D ),
    .q(\DFF_358.Q )
  );
  al_dffl _10857_ (
    .clk(CK),
    .d(\DFF_359.D ),
    .q(\DFF_359.Q )
  );
  al_dffl _10858_ (
    .clk(CK),
    .d(\DFF_361.D ),
    .q(\DFF_361.Q )
  );
  al_dffl _10859_ (
    .clk(CK),
    .d(\DFF_362.D ),
    .q(\DFF_362.Q )
  );
  al_dffl _10860_ (
    .clk(CK),
    .d(\DFF_363.D ),
    .q(\DFF_363.Q )
  );
  al_dffl _10861_ (
    .clk(CK),
    .d(\DFF_364.D ),
    .q(\DFF_364.Q )
  );
  al_dffl _10862_ (
    .clk(CK),
    .d(\DFF_376.D ),
    .q(\DFF_376.Q )
  );
  al_dffl _10863_ (
    .clk(CK),
    .d(\DFF_376.Q ),
    .q(\DFF_365.Q )
  );
  al_dffl _10864_ (
    .clk(CK),
    .d(\DFF_366.D ),
    .q(\DFF_366.Q )
  );
  al_dffl _10865_ (
    .clk(CK),
    .d(\DFF_181.Q ),
    .q(\DFF_785.Q )
  );
  al_dffl _10866_ (
    .clk(CK),
    .d(\DFF_785.Q ),
    .q(\DFF_642.Q )
  );
  al_dffl _10867_ (
    .clk(CK),
    .d(\DFF_642.Q ),
    .q(\DFF_367.Q )
  );
  al_dffl _10868_ (
    .clk(CK),
    .d(\DFF_368.D ),
    .q(\DFF_368.Q )
  );
  al_dffl _10869_ (
    .clk(CK),
    .d(\DFF_370.D ),
    .q(\DFF_370.Q )
  );
  al_dffl _10870_ (
    .clk(CK),
    .d(\DFF_146.Q ),
    .q(\DFF_1110.Q )
  );
  al_dffl _10871_ (
    .clk(CK),
    .d(\DFF_1110.Q ),
    .q(\DFF_372.Q )
  );
  al_dffl _10872_ (
    .clk(CK),
    .d(\DFF_1225.D ),
    .q(\DFF_1225.Q )
  );
  al_dffl _10873_ (
    .clk(CK),
    .d(\DFF_1225.Q ),
    .q(\DFF_373.Q )
  );
  al_dffl _10874_ (
    .clk(CK),
    .d(\DFF_374.D ),
    .q(\DFF_374.Q )
  );
  al_dffl _10875_ (
    .clk(CK),
    .d(\DFF_375.D ),
    .q(\DFF_375.Q )
  );
  al_dffl _10876_ (
    .clk(CK),
    .d(\DFF_1316.D ),
    .q(\DFF_1316.Q )
  );
  al_dffl _10877_ (
    .clk(CK),
    .d(\DFF_1316.Q ),
    .q(\DFF_377.Q )
  );
  al_dffl _10878_ (
    .clk(CK),
    .d(\DFF_378.D ),
    .q(\DFF_378.Q )
  );
  al_dffl _10879_ (
    .clk(CK),
    .d(\DFF_379.D ),
    .q(\DFF_379.Q )
  );
  al_dffl _10880_ (
    .clk(CK),
    .d(\DFF_152.Q ),
    .q(\DFF_404.Q )
  );
  al_dffl _10881_ (
    .clk(CK),
    .d(\DFF_404.Q ),
    .q(\DFF_380.Q )
  );
  al_dffl _10882_ (
    .clk(CK),
    .d(\DFF_381.D ),
    .q(\DFF_381.Q )
  );
  al_dffl _10883_ (
    .clk(CK),
    .d(\DFF_382.D ),
    .q(\DFF_382.Q )
  );
  al_dffl _10884_ (
    .clk(CK),
    .d(\DFF_383.D ),
    .q(\DFF_383.Q )
  );
  al_dffl _10885_ (
    .clk(CK),
    .d(\DFF_384.D ),
    .q(\DFF_384.Q )
  );
  al_dffl _10886_ (
    .clk(CK),
    .d(\DFF_385.D ),
    .q(\DFF_385.Q )
  );
  al_dffl _10887_ (
    .clk(CK),
    .d(\DFF_386.D ),
    .q(\DFF_386.Q )
  );
  al_dffl _10888_ (
    .clk(CK),
    .d(\DFF_387.D ),
    .q(\DFF_387.Q )
  );
  al_dffl _10889_ (
    .clk(CK),
    .d(\DFF_388.D ),
    .q(\DFF_388.Q )
  );
  al_dffl _10890_ (
    .clk(CK),
    .d(\DFF_390.D ),
    .q(\DFF_390.Q )
  );
  al_dffl _10891_ (
    .clk(CK),
    .d(\DFF_391.D ),
    .q(\DFF_391.Q )
  );
  al_dffl _10892_ (
    .clk(CK),
    .d(\DFF_392.D ),
    .q(\DFF_392.Q )
  );
  al_dffl _10893_ (
    .clk(CK),
    .d(\DFF_393.D ),
    .q(\DFF_393.Q )
  );
  al_dffl _10894_ (
    .clk(CK),
    .d(\DFF_394.D ),
    .q(\DFF_394.Q )
  );
  al_dffl _10895_ (
    .clk(CK),
    .d(\DFF_395.D ),
    .q(\DFF_395.Q )
  );
  al_dffl _10896_ (
    .clk(CK),
    .d(\DFF_396.D ),
    .q(\DFF_396.Q )
  );
  al_dffl _10897_ (
    .clk(CK),
    .d(\DFF_397.D ),
    .q(\DFF_397.Q )
  );
  al_dffl _10898_ (
    .clk(CK),
    .d(\DFF_398.D ),
    .q(\DFF_398.Q )
  );
  al_dffl _10899_ (
    .clk(CK),
    .d(\DFF_399.D ),
    .q(\DFF_399.Q )
  );
  al_dffl _10900_ (
    .clk(CK),
    .d(\DFF_400.D ),
    .q(\DFF_400.Q )
  );
  al_dffl _10901_ (
    .clk(CK),
    .d(\DFF_402.D ),
    .q(\DFF_402.Q )
  );
  al_dffl _10902_ (
    .clk(CK),
    .d(\DFF_403.D ),
    .q(\DFF_403.Q )
  );
  al_dffl _10903_ (
    .clk(CK),
    .d(\DFF_405.D ),
    .q(\DFF_405.Q )
  );
  al_dffl _10904_ (
    .clk(CK),
    .d(\DFF_406.D ),
    .q(\DFF_406.Q )
  );
  al_dffl _10905_ (
    .clk(CK),
    .d(\DFF_407.D ),
    .q(\DFF_407.Q )
  );
  al_dffl _10906_ (
    .clk(CK),
    .d(\DFF_334.Q ),
    .q(\DFF_408.Q )
  );
  al_dffl _10907_ (
    .clk(CK),
    .d(\DFF_409.D ),
    .q(\DFF_409.Q )
  );
  al_dffl _10908_ (
    .clk(CK),
    .d(\DFF_410.D ),
    .q(\DFF_410.Q )
  );
  al_dffl _10909_ (
    .clk(CK),
    .d(\DFF_411.D ),
    .q(\DFF_411.Q )
  );
  al_dffl _10910_ (
    .clk(CK),
    .d(\DFF_412.D ),
    .q(\DFF_412.Q )
  );
  al_dffl _10911_ (
    .clk(CK),
    .d(\DFF_413.D ),
    .q(\DFF_413.Q )
  );
  al_dffl _10912_ (
    .clk(CK),
    .d(\DFF_414.D ),
    .q(\DFF_414.Q )
  );
  al_dffl _10913_ (
    .clk(CK),
    .d(\DFF_415.D ),
    .q(\DFF_415.Q )
  );
  al_dffl _10914_ (
    .clk(CK),
    .d(\DFF_416.D ),
    .q(\DFF_416.Q )
  );
  al_dffl _10915_ (
    .clk(CK),
    .d(\DFF_417.D ),
    .q(\DFF_417.Q )
  );
  al_dffl _10916_ (
    .clk(CK),
    .d(\DFF_419.D ),
    .q(\DFF_419.Q )
  );
  al_dffl _10917_ (
    .clk(CK),
    .d(\DFF_420.D ),
    .q(\DFF_420.Q )
  );
  al_dffl _10918_ (
    .clk(CK),
    .d(\DFF_421.D ),
    .q(\DFF_421.Q )
  );
  al_dffl _10919_ (
    .clk(CK),
    .d(\DFF_423.D ),
    .q(\DFF_423.Q )
  );
  al_dffl _10920_ (
    .clk(CK),
    .d(\DFF_424.D ),
    .q(\DFF_424.Q )
  );
  al_dffl _10921_ (
    .clk(CK),
    .d(\DFF_425.D ),
    .q(\DFF_425.Q )
  );
  al_dffl _10922_ (
    .clk(CK),
    .d(\DFF_426.D ),
    .q(\DFF_426.Q )
  );
  al_dffl _10923_ (
    .clk(CK),
    .d(\DFF_427.D ),
    .q(\DFF_427.Q )
  );
  al_dffl _10924_ (
    .clk(CK),
    .d(\DFF_428.D ),
    .q(\DFF_428.Q )
  );
  al_dffl _10925_ (
    .clk(CK),
    .d(\DFF_429.D ),
    .q(\DFF_429.Q )
  );
  al_dffl _10926_ (
    .clk(CK),
    .d(\DFF_430.D ),
    .q(\DFF_430.Q )
  );
  al_dffl _10927_ (
    .clk(CK),
    .d(\DFF_431.D ),
    .q(\DFF_431.Q )
  );
  al_dffl _10928_ (
    .clk(CK),
    .d(\DFF_432.D ),
    .q(\DFF_432.Q )
  );
  al_dffl _10929_ (
    .clk(CK),
    .d(\DFF_433.D ),
    .q(\DFF_433.Q )
  );
  al_dffl _10930_ (
    .clk(CK),
    .d(\DFF_434.D ),
    .q(\DFF_434.Q )
  );
  al_dffl _10931_ (
    .clk(CK),
    .d(\DFF_435.D ),
    .q(\DFF_435.Q )
  );
  al_dffl _10932_ (
    .clk(CK),
    .d(\DFF_436.D ),
    .q(\DFF_436.Q )
  );
  al_dffl _10933_ (
    .clk(CK),
    .d(\DFF_437.D ),
    .q(\DFF_437.Q )
  );
  al_dffl _10934_ (
    .clk(CK),
    .d(\DFF_438.D ),
    .q(\DFF_438.Q )
  );
  al_dffl _10935_ (
    .clk(CK),
    .d(\DFF_439.D ),
    .q(\DFF_439.Q )
  );
  al_dffl _10936_ (
    .clk(CK),
    .d(\DFF_440.D ),
    .q(\DFF_440.Q )
  );
  al_dffl _10937_ (
    .clk(CK),
    .d(\DFF_441.D ),
    .q(\DFF_441.Q )
  );
  al_dffl _10938_ (
    .clk(CK),
    .d(\DFF_442.D ),
    .q(\DFF_442.Q )
  );
  al_dffl _10939_ (
    .clk(CK),
    .d(\DFF_443.D ),
    .q(\DFF_443.Q )
  );
  al_dffl _10940_ (
    .clk(CK),
    .d(\DFF_444.D ),
    .q(\DFF_444.Q )
  );
  al_dffl _10941_ (
    .clk(CK),
    .d(\DFF_445.D ),
    .q(\DFF_445.Q )
  );
  al_dffl _10942_ (
    .clk(CK),
    .d(\DFF_446.D ),
    .q(\DFF_446.Q )
  );
  al_dffl _10943_ (
    .clk(CK),
    .d(\DFF_447.D ),
    .q(\DFF_447.Q )
  );
  al_dffl _10944_ (
    .clk(CK),
    .d(\DFF_448.D ),
    .q(\DFF_448.Q )
  );
  al_dffl _10945_ (
    .clk(CK),
    .d(\DFF_449.D ),
    .q(\DFF_449.Q )
  );
  al_dffl _10946_ (
    .clk(CK),
    .d(\DFF_460.D ),
    .q(\DFF_460.Q )
  );
  al_dffl _10947_ (
    .clk(CK),
    .d(\DFF_460.Q ),
    .q(\DFF_450.Q )
  );
  al_dffl _10948_ (
    .clk(CK),
    .d(\DFF_451.D ),
    .q(\DFF_451.Q )
  );
  al_dffl _10949_ (
    .clk(CK),
    .d(\DFF_452.D ),
    .q(\DFF_452.Q )
  );
  al_dffl _10950_ (
    .clk(CK),
    .d(\DFF_453.D ),
    .q(\DFF_453.Q )
  );
  al_dffl _10951_ (
    .clk(CK),
    .d(\DFF_454.D ),
    .q(\DFF_454.Q )
  );
  al_dffl _10952_ (
    .clk(CK),
    .d(\DFF_455.D ),
    .q(\DFF_455.Q )
  );
  al_dffl _10953_ (
    .clk(CK),
    .d(\DFF_456.D ),
    .q(\DFF_456.Q )
  );
  al_dffl _10954_ (
    .clk(CK),
    .d(\DFF_457.D ),
    .q(\DFF_457.Q )
  );
  al_dffl _10955_ (
    .clk(CK),
    .d(\DFF_678.D ),
    .q(\DFF_678.Q )
  );
  al_dffl _10956_ (
    .clk(CK),
    .d(\DFF_678.Q ),
    .q(\DFF_458.Q )
  );
  al_dffl _10957_ (
    .clk(CK),
    .d(\DFF_459.D ),
    .q(\DFF_459.Q )
  );
  al_dffl _10958_ (
    .clk(CK),
    .d(\DFF_461.D ),
    .q(\DFF_461.Q )
  );
  al_dffl _10959_ (
    .clk(CK),
    .d(\DFF_462.D ),
    .q(\DFF_462.Q )
  );
  al_dffl _10960_ (
    .clk(CK),
    .d(\DFF_463.D ),
    .q(\DFF_463.Q )
  );
  al_dffl _10961_ (
    .clk(CK),
    .d(\DFF_464.D ),
    .q(\DFF_464.Q )
  );
  al_dffl _10962_ (
    .clk(CK),
    .d(\DFF_465.D ),
    .q(\DFF_465.Q )
  );
  al_dffl _10963_ (
    .clk(CK),
    .d(\DFF_466.D ),
    .q(\DFF_466.Q )
  );
  al_dffl _10964_ (
    .clk(CK),
    .d(\DFF_467.D ),
    .q(\DFF_467.Q )
  );
  al_dffl _10965_ (
    .clk(CK),
    .d(\DFF_469.D ),
    .q(\DFF_469.Q )
  );
  al_dffl _10966_ (
    .clk(CK),
    .d(\DFF_470.D ),
    .q(\DFF_470.Q )
  );
  al_dffl _10967_ (
    .clk(CK),
    .d(\DFF_471.D ),
    .q(\DFF_471.Q )
  );
  al_dffl _10968_ (
    .clk(CK),
    .d(\DFF_472.D ),
    .q(\DFF_472.Q )
  );
  al_dffl _10969_ (
    .clk(CK),
    .d(\DFF_473.D ),
    .q(\DFF_473.Q )
  );
  al_dffl _10970_ (
    .clk(CK),
    .d(\DFF_475.D ),
    .q(\DFF_475.Q )
  );
  al_dffl _10971_ (
    .clk(CK),
    .d(\DFF_476.D ),
    .q(\DFF_476.Q )
  );
  al_dffl _10972_ (
    .clk(CK),
    .d(\DFF_477.D ),
    .q(\DFF_477.Q )
  );
  al_dffl _10973_ (
    .clk(CK),
    .d(\DFF_478.D ),
    .q(\DFF_478.Q )
  );
  al_dffl _10974_ (
    .clk(CK),
    .d(\DFF_479.D ),
    .q(\DFF_479.Q )
  );
  al_dffl _10975_ (
    .clk(CK),
    .d(\DFF_1234.D ),
    .q(\DFF_1234.Q )
  );
  al_dffl _10976_ (
    .clk(CK),
    .d(\DFF_1234.Q ),
    .q(\DFF_480.Q )
  );
  al_dffl _10977_ (
    .clk(CK),
    .d(\DFF_1275.D ),
    .q(\DFF_1275.Q )
  );
  al_dffl _10978_ (
    .clk(CK),
    .d(\DFF_1275.Q ),
    .q(\DFF_481.Q )
  );
  al_dffl _10979_ (
    .clk(CK),
    .d(\DFF_482.D ),
    .q(\DFF_482.Q )
  );
  al_dffl _10980_ (
    .clk(CK),
    .d(\DFF_483.D ),
    .q(\DFF_483.Q )
  );
  al_dffl _10981_ (
    .clk(CK),
    .d(\DFF_484.D ),
    .q(\DFF_484.Q )
  );
  al_dffl _10982_ (
    .clk(CK),
    .d(\DFF_486.D ),
    .q(\DFF_486.Q )
  );
  al_dffl _10983_ (
    .clk(CK),
    .d(\DFF_487.D ),
    .q(\DFF_487.Q )
  );
  al_dffl _10984_ (
    .clk(CK),
    .d(\DFF_488.D ),
    .q(\DFF_488.Q )
  );
  al_dffl _10985_ (
    .clk(CK),
    .d(\DFF_489.D ),
    .q(\DFF_489.Q )
  );
  al_dffl _10986_ (
    .clk(CK),
    .d(\DFF_490.D ),
    .q(\DFF_490.Q )
  );
  al_dffl _10987_ (
    .clk(CK),
    .d(\DFF_491.D ),
    .q(\DFF_491.Q )
  );
  al_dffl _10988_ (
    .clk(CK),
    .d(\DFF_1414.D ),
    .q(\DFF_1414.Q )
  );
  al_dffl _10989_ (
    .clk(CK),
    .d(\DFF_1414.Q ),
    .q(\DFF_492.Q )
  );
  al_dffl _10990_ (
    .clk(CK),
    .d(\DFF_493.D ),
    .q(\DFF_493.Q )
  );
  al_dffl _10991_ (
    .clk(CK),
    .d(\DFF_494.D ),
    .q(\DFF_494.Q )
  );
  al_dffl _10992_ (
    .clk(CK),
    .d(\DFF_495.D ),
    .q(\DFF_495.Q )
  );
  al_dffl _10993_ (
    .clk(CK),
    .d(\DFF_496.D ),
    .q(\DFF_496.Q )
  );
  al_dffl _10994_ (
    .clk(CK),
    .d(\DFF_497.D ),
    .q(\DFF_497.Q )
  );
  al_dffl _10995_ (
    .clk(CK),
    .d(\DFF_498.D ),
    .q(\DFF_498.Q )
  );
  al_dffl _10996_ (
    .clk(CK),
    .d(\DFF_499.D ),
    .q(\DFF_499.Q )
  );
  al_dffl _10997_ (
    .clk(CK),
    .d(\DFF_500.D ),
    .q(\DFF_500.Q )
  );
  al_dffl _10998_ (
    .clk(CK),
    .d(\DFF_501.D ),
    .q(\DFF_501.Q )
  );
  al_dffl _10999_ (
    .clk(CK),
    .d(\DFF_502.D ),
    .q(\DFF_502.Q )
  );
  al_dffl _11000_ (
    .clk(CK),
    .d(\DFF_503.D ),
    .q(\DFF_503.Q )
  );
  al_dffl _11001_ (
    .clk(CK),
    .d(\DFF_504.D ),
    .q(\DFF_504.Q )
  );
  al_dffl _11002_ (
    .clk(CK),
    .d(\DFF_505.D ),
    .q(\DFF_505.Q )
  );
  al_dffl _11003_ (
    .clk(CK),
    .d(\DFF_506.D ),
    .q(\DFF_506.Q )
  );
  al_dffl _11004_ (
    .clk(CK),
    .d(\DFF_507.D ),
    .q(\DFF_507.Q )
  );
  al_dffl _11005_ (
    .clk(CK),
    .d(\DFF_508.D ),
    .q(\DFF_508.Q )
  );
  al_dffl _11006_ (
    .clk(CK),
    .d(\DFF_203.Q ),
    .q(\DFF_509.Q )
  );
  al_dffl _11007_ (
    .clk(CK),
    .d(\DFF_510.D ),
    .q(\DFF_510.Q )
  );
  al_dffl _11008_ (
    .clk(CK),
    .d(\DFF_675.D ),
    .q(\DFF_675.Q )
  );
  al_dffl _11009_ (
    .clk(CK),
    .d(\DFF_675.Q ),
    .q(\DFF_1308.Q )
  );
  al_dffl _11010_ (
    .clk(CK),
    .d(\DFF_1308.Q ),
    .q(\DFF_511.Q )
  );
  al_dffl _11011_ (
    .clk(CK),
    .d(\DFF_512.D ),
    .q(\DFF_512.Q )
  );
  al_dffl _11012_ (
    .clk(CK),
    .d(\DFF_513.D ),
    .q(\DFF_513.Q )
  );
  al_dffl _11013_ (
    .clk(CK),
    .d(\DFF_514.D ),
    .q(\DFF_514.Q )
  );
  al_dffl _11014_ (
    .clk(CK),
    .d(\DFF_516.D ),
    .q(\DFF_516.Q )
  );
  al_dffl _11015_ (
    .clk(CK),
    .d(\DFF_517.D ),
    .q(\DFF_517.Q )
  );
  al_dffl _11016_ (
    .clk(CK),
    .d(\DFF_518.D ),
    .q(\DFF_518.Q )
  );
  al_dffl _11017_ (
    .clk(CK),
    .d(\DFF_519.D ),
    .q(\DFF_519.Q )
  );
  al_dffl _11018_ (
    .clk(CK),
    .d(\DFF_520.D ),
    .q(\DFF_520.Q )
  );
  al_dffl _11019_ (
    .clk(CK),
    .d(\DFF_521.D ),
    .q(\DFF_521.Q )
  );
  al_dffl _11020_ (
    .clk(CK),
    .d(\DFF_522.D ),
    .q(\DFF_522.Q )
  );
  al_dffl _11021_ (
    .clk(CK),
    .d(\DFF_523.D ),
    .q(\DFF_523.Q )
  );
  al_dffl _11022_ (
    .clk(CK),
    .d(\DFF_524.D ),
    .q(\DFF_524.Q )
  );
  al_dffl _11023_ (
    .clk(CK),
    .d(\DFF_525.D ),
    .q(\DFF_525.Q )
  );
  al_dffl _11024_ (
    .clk(CK),
    .d(\DFF_526.D ),
    .q(\DFF_526.Q )
  );
  al_dffl _11025_ (
    .clk(CK),
    .d(\DFF_527.D ),
    .q(\DFF_527.Q )
  );
  al_dffl _11026_ (
    .clk(CK),
    .d(\DFF_530.D ),
    .q(\DFF_530.Q )
  );
  al_dffl _11027_ (
    .clk(CK),
    .d(\DFF_531.D ),
    .q(\DFF_531.Q )
  );
  al_dffl _11028_ (
    .clk(CK),
    .d(\DFF_532.D ),
    .q(\DFF_532.Q )
  );
  al_dffl _11029_ (
    .clk(CK),
    .d(\DFF_533.D ),
    .q(\DFF_533.Q )
  );
  al_dffl _11030_ (
    .clk(CK),
    .d(\DFF_534.D ),
    .q(\DFF_534.Q )
  );
  al_dffl _11031_ (
    .clk(CK),
    .d(\DFF_535.D ),
    .q(\DFF_535.Q )
  );
  al_dffl _11032_ (
    .clk(CK),
    .d(\DFF_536.D ),
    .q(\DFF_536.Q )
  );
  al_dffl _11033_ (
    .clk(CK),
    .d(\DFF_538.D ),
    .q(\DFF_538.Q )
  );
  al_dffl _11034_ (
    .clk(CK),
    .d(\DFF_539.D ),
    .q(\DFF_539.Q )
  );
  al_dffl _11035_ (
    .clk(CK),
    .d(\DFF_540.D ),
    .q(\DFF_540.Q )
  );
  al_dffl _11036_ (
    .clk(CK),
    .d(\DFF_541.D ),
    .q(\DFF_541.Q )
  );
  al_dffl _11037_ (
    .clk(CK),
    .d(\DFF_542.D ),
    .q(\DFF_542.Q )
  );
  al_dffl _11038_ (
    .clk(CK),
    .d(\DFF_543.D ),
    .q(\DFF_543.Q )
  );
  al_dffl _11039_ (
    .clk(CK),
    .d(\DFF_544.D ),
    .q(\DFF_544.Q )
  );
  al_dffl _11040_ (
    .clk(CK),
    .d(\DFF_545.D ),
    .q(\DFF_545.Q )
  );
  al_dffl _11041_ (
    .clk(CK),
    .d(\DFF_546.D ),
    .q(\DFF_546.Q )
  );
  al_dffl _11042_ (
    .clk(CK),
    .d(\DFF_547.D ),
    .q(\DFF_547.Q )
  );
  al_dffl _11043_ (
    .clk(CK),
    .d(\DFF_548.D ),
    .q(\DFF_548.Q )
  );
  al_dffl _11044_ (
    .clk(CK),
    .d(\DFF_549.D ),
    .q(\DFF_549.Q )
  );
  al_dffl _11045_ (
    .clk(CK),
    .d(\DFF_550.D ),
    .q(\DFF_550.Q )
  );
  al_dffl _11046_ (
    .clk(CK),
    .d(\DFF_551.D ),
    .q(\DFF_551.Q )
  );
  al_dffl _11047_ (
    .clk(CK),
    .d(\DFF_552.D ),
    .q(\DFF_552.Q )
  );
  al_dffl _11048_ (
    .clk(CK),
    .d(\DFF_86.Q ),
    .q(\DFF_553.Q )
  );
  al_dffl _11049_ (
    .clk(CK),
    .d(\DFF_555.D ),
    .q(\DFF_555.Q )
  );
  al_dffl _11050_ (
    .clk(CK),
    .d(\DFF_556.D ),
    .q(\DFF_556.Q )
  );
  al_dffl _11051_ (
    .clk(CK),
    .d(\DFF_557.D ),
    .q(\DFF_557.Q )
  );
  al_dffl _11052_ (
    .clk(CK),
    .d(\DFF_558.D ),
    .q(\DFF_558.Q )
  );
  al_dffl _11053_ (
    .clk(CK),
    .d(\DFF_559.D ),
    .q(\DFF_559.Q )
  );
  al_dffl _11054_ (
    .clk(CK),
    .d(\DFF_560.D ),
    .q(\DFF_560.Q )
  );
  al_dffl _11055_ (
    .clk(CK),
    .d(\DFF_562.D ),
    .q(\DFF_562.Q )
  );
  al_dffl _11056_ (
    .clk(CK),
    .d(\DFF_563.D ),
    .q(\DFF_563.Q )
  );
  al_dffl _11057_ (
    .clk(CK),
    .d(\DFF_564.D ),
    .q(\DFF_564.Q )
  );
  al_dffl _11058_ (
    .clk(CK),
    .d(\DFF_480.Q ),
    .q(\DFF_909.Q )
  );
  al_dffl _11059_ (
    .clk(CK),
    .d(\DFF_909.Q ),
    .q(\DFF_565.Q )
  );
  al_dffl _11060_ (
    .clk(CK),
    .d(\DFF_567.D ),
    .q(\DFF_567.Q )
  );
  al_dffl _11061_ (
    .clk(CK),
    .d(\DFF_568.D ),
    .q(\DFF_568.Q )
  );
  al_dffl _11062_ (
    .clk(CK),
    .d(\DFF_503.Q ),
    .q(\DFF_569.Q )
  );
  al_dffl _11063_ (
    .clk(CK),
    .d(\DFF_570.D ),
    .q(\DFF_570.Q )
  );
  al_dffl _11064_ (
    .clk(CK),
    .d(\DFF_571.D ),
    .q(\DFF_571.Q )
  );
  al_dffl _11065_ (
    .clk(CK),
    .d(\DFF_572.D ),
    .q(\DFF_572.Q )
  );
  al_dffl _11066_ (
    .clk(CK),
    .d(\DFF_573.D ),
    .q(\DFF_573.Q )
  );
  al_dffl _11067_ (
    .clk(CK),
    .d(\DFF_574.D ),
    .q(\DFF_574.Q )
  );
  al_dffl _11068_ (
    .clk(CK),
    .d(\DFF_575.D ),
    .q(\DFF_575.Q )
  );
  al_dffl _11069_ (
    .clk(CK),
    .d(\DFF_576.D ),
    .q(\DFF_576.Q )
  );
  al_dffl _11070_ (
    .clk(CK),
    .d(\DFF_577.D ),
    .q(\DFF_577.Q )
  );
  al_dffl _11071_ (
    .clk(CK),
    .d(\DFF_578.D ),
    .q(\DFF_578.Q )
  );
  al_dffl _11072_ (
    .clk(CK),
    .d(\DFF_579.D ),
    .q(\DFF_579.Q )
  );
  al_dffl _11073_ (
    .clk(CK),
    .d(\DFF_580.D ),
    .q(\DFF_580.Q )
  );
  al_dffl _11074_ (
    .clk(CK),
    .d(\DFF_581.D ),
    .q(\DFF_581.Q )
  );
  al_dffl _11075_ (
    .clk(CK),
    .d(\DFF_582.D ),
    .q(\DFF_582.Q )
  );
  al_dffl _11076_ (
    .clk(CK),
    .d(\DFF_583.D ),
    .q(\DFF_583.Q )
  );
  al_dffl _11077_ (
    .clk(CK),
    .d(\DFF_584.D ),
    .q(\DFF_584.Q )
  );
  al_dffl _11078_ (
    .clk(CK),
    .d(\DFF_586.D ),
    .q(\DFF_586.Q )
  );
  al_dffl _11079_ (
    .clk(CK),
    .d(\DFF_587.D ),
    .q(\DFF_587.Q )
  );
  al_dffl _11080_ (
    .clk(CK),
    .d(\DFF_588.D ),
    .q(\DFF_588.Q )
  );
  al_dffl _11081_ (
    .clk(CK),
    .d(\DFF_589.D ),
    .q(\DFF_589.Q )
  );
  al_dffl _11082_ (
    .clk(CK),
    .d(\DFF_590.D ),
    .q(\DFF_590.Q )
  );
  al_dffl _11083_ (
    .clk(CK),
    .d(\DFF_591.D ),
    .q(\DFF_591.Q )
  );
  al_dffl _11084_ (
    .clk(CK),
    .d(\DFF_592.D ),
    .q(\DFF_592.Q )
  );
  al_dffl _11085_ (
    .clk(CK),
    .d(\DFF_593.D ),
    .q(\DFF_593.Q )
  );
  al_dffl _11086_ (
    .clk(CK),
    .d(\DFF_594.D ),
    .q(\DFF_594.Q )
  );
  al_dffl _11087_ (
    .clk(CK),
    .d(\DFF_595.D ),
    .q(\DFF_595.Q )
  );
  al_dffl _11088_ (
    .clk(CK),
    .d(\DFF_596.D ),
    .q(\DFF_596.Q )
  );
  al_dffl _11089_ (
    .clk(CK),
    .d(\DFF_597.D ),
    .q(\DFF_597.Q )
  );
  al_dffl _11090_ (
    .clk(CK),
    .d(\DFF_598.D ),
    .q(\DFF_598.Q )
  );
  al_dffl _11091_ (
    .clk(CK),
    .d(\DFF_599.D ),
    .q(\DFF_599.Q )
  );
  al_dffl _11092_ (
    .clk(CK),
    .d(\DFF_1207.D ),
    .q(\DFF_1207.Q )
  );
  al_dffl _11093_ (
    .clk(CK),
    .d(\DFF_1207.Q ),
    .q(\DFF_600.Q )
  );
  al_dffl _11094_ (
    .clk(CK),
    .d(\DFF_601.D ),
    .q(\DFF_601.Q )
  );
  al_dffl _11095_ (
    .clk(CK),
    .d(\DFF_602.D ),
    .q(\DFF_602.Q )
  );
  al_dffl _11096_ (
    .clk(CK),
    .d(\DFF_861.D ),
    .q(\DFF_861.Q )
  );
  al_dffl _11097_ (
    .clk(CK),
    .d(\DFF_861.Q ),
    .q(\DFF_603.Q )
  );
  al_dffl _11098_ (
    .clk(CK),
    .d(\DFF_604.D ),
    .q(\DFF_604.Q )
  );
  al_dffl _11099_ (
    .clk(CK),
    .d(\DFF_605.D ),
    .q(\DFF_605.Q )
  );
  al_dffl _11100_ (
    .clk(CK),
    .d(\DFF_606.D ),
    .q(\DFF_606.Q )
  );
  al_dffl _11101_ (
    .clk(CK),
    .d(\DFF_607.D ),
    .q(\DFF_607.Q )
  );
  al_dffl _11102_ (
    .clk(CK),
    .d(\DFF_608.D ),
    .q(\DFF_608.Q )
  );
  al_dffl _11103_ (
    .clk(CK),
    .d(\DFF_609.D ),
    .q(\DFF_609.Q )
  );
  al_dffl _11104_ (
    .clk(CK),
    .d(\DFF_610.D ),
    .q(\DFF_610.Q )
  );
  al_dffl _11105_ (
    .clk(CK),
    .d(\DFF_611.D ),
    .q(\DFF_611.Q )
  );
  al_dffl _11106_ (
    .clk(CK),
    .d(\DFF_612.D ),
    .q(\DFF_612.Q )
  );
  al_dffl _11107_ (
    .clk(CK),
    .d(\DFF_234.Q ),
    .q(\DFF_613.Q )
  );
  al_dffl _11108_ (
    .clk(CK),
    .d(\DFF_614.D ),
    .q(\DFF_614.Q )
  );
  al_dffl _11109_ (
    .clk(CK),
    .d(\DFF_549.Q ),
    .q(\DFF_615.Q )
  );
  al_dffl _11110_ (
    .clk(CK),
    .d(\DFF_617.D ),
    .q(\DFF_617.Q )
  );
  al_dffl _11111_ (
    .clk(CK),
    .d(\DFF_618.D ),
    .q(\DFF_618.Q )
  );
  al_dffl _11112_ (
    .clk(CK),
    .d(\DFF_619.D ),
    .q(\DFF_619.Q )
  );
  al_dffl _11113_ (
    .clk(CK),
    .d(\DFF_620.D ),
    .q(\DFF_620.Q )
  );
  al_dffl _11114_ (
    .clk(CK),
    .d(\DFF_621.D ),
    .q(\DFF_621.Q )
  );
  al_dffl _11115_ (
    .clk(CK),
    .d(\DFF_622.D ),
    .q(\DFF_622.Q )
  );
  al_dffl _11116_ (
    .clk(CK),
    .d(\DFF_623.D ),
    .q(\DFF_623.Q )
  );
  al_dffl _11117_ (
    .clk(CK),
    .d(\DFF_624.D ),
    .q(\DFF_624.Q )
  );
  al_dffl _11118_ (
    .clk(CK),
    .d(\DFF_625.D ),
    .q(\DFF_625.Q )
  );
  al_dffl _11119_ (
    .clk(CK),
    .d(\DFF_626.D ),
    .q(\DFF_626.Q )
  );
  al_dffl _11120_ (
    .clk(CK),
    .d(\DFF_627.D ),
    .q(\DFF_627.Q )
  );
  al_dffl _11121_ (
    .clk(CK),
    .d(\DFF_628.D ),
    .q(\DFF_628.Q )
  );
  al_dffl _11122_ (
    .clk(CK),
    .d(\DFF_629.D ),
    .q(\DFF_629.Q )
  );
  al_dffl _11123_ (
    .clk(CK),
    .d(\DFF_630.D ),
    .q(\DFF_630.Q )
  );
  al_dffl _11124_ (
    .clk(CK),
    .d(\DFF_631.D ),
    .q(\DFF_631.Q )
  );
  al_dffl _11125_ (
    .clk(CK),
    .d(\DFF_632.D ),
    .q(\DFF_632.Q )
  );
  al_dffl _11126_ (
    .clk(CK),
    .d(\DFF_633.D ),
    .q(\DFF_633.Q )
  );
  al_dffl _11127_ (
    .clk(CK),
    .d(\DFF_634.D ),
    .q(\DFF_634.Q )
  );
  al_dffl _11128_ (
    .clk(CK),
    .d(\DFF_635.D ),
    .q(\DFF_635.Q )
  );
  al_dffl _11129_ (
    .clk(CK),
    .d(\DFF_636.D ),
    .q(\DFF_636.Q )
  );
  al_dffl _11130_ (
    .clk(CK),
    .d(\DFF_637.D ),
    .q(\DFF_637.Q )
  );
  al_dffl _11131_ (
    .clk(CK),
    .d(\DFF_638.D ),
    .q(\DFF_638.Q )
  );
  al_dffl _11132_ (
    .clk(CK),
    .d(\DFF_639.D ),
    .q(\DFF_639.Q )
  );
  al_dffl _11133_ (
    .clk(CK),
    .d(\DFF_640.D ),
    .q(\DFF_640.Q )
  );
  al_dffl _11134_ (
    .clk(CK),
    .d(\DFF_641.D ),
    .q(\DFF_641.Q )
  );
  al_dffl _11135_ (
    .clk(CK),
    .d(\DFF_644.D ),
    .q(\DFF_644.Q )
  );
  al_dffl _11136_ (
    .clk(CK),
    .d(\DFF_645.D ),
    .q(\DFF_645.Q )
  );
  al_dffl _11137_ (
    .clk(CK),
    .d(\DFF_646.D ),
    .q(\DFF_646.Q )
  );
  al_dffl _11138_ (
    .clk(CK),
    .d(\DFF_647.D ),
    .q(\DFF_647.Q )
  );
  al_dffl _11139_ (
    .clk(CK),
    .d(\DFF_648.D ),
    .q(\DFF_648.Q )
  );
  al_dffl _11140_ (
    .clk(CK),
    .d(\DFF_649.D ),
    .q(\DFF_649.Q )
  );
  al_dffl _11141_ (
    .clk(CK),
    .d(g6752),
    .q(\DFF_650.Q )
  );
  al_dffl _11142_ (
    .clk(CK),
    .d(\DFF_651.D ),
    .q(\DFF_651.Q )
  );
  al_dffl _11143_ (
    .clk(CK),
    .d(\DFF_652.D ),
    .q(\DFF_652.Q )
  );
  al_dffl _11144_ (
    .clk(CK),
    .d(\DFF_653.D ),
    .q(\DFF_653.Q )
  );
  al_dffl _11145_ (
    .clk(CK),
    .d(\DFF_654.D ),
    .q(\DFF_654.Q )
  );
  al_dffl _11146_ (
    .clk(CK),
    .d(\DFF_656.D ),
    .q(\DFF_656.Q )
  );
  al_dffl _11147_ (
    .clk(CK),
    .d(\DFF_657.D ),
    .q(\DFF_657.Q )
  );
  al_dffl _11148_ (
    .clk(CK),
    .d(\DFF_658.D ),
    .q(\DFF_658.Q )
  );
  al_dffl _11149_ (
    .clk(CK),
    .d(\DFF_659.D ),
    .q(\DFF_659.Q )
  );
  al_dffl _11150_ (
    .clk(CK),
    .d(\DFF_660.D ),
    .q(\DFF_660.Q )
  );
  al_dffl _11151_ (
    .clk(CK),
    .d(\DFF_661.D ),
    .q(\DFF_661.Q )
  );
  al_dffl _11152_ (
    .clk(CK),
    .d(\DFF_367.Q ),
    .q(\DFF_662.Q )
  );
  al_dffl _11153_ (
    .clk(CK),
    .d(\DFF_1265.D ),
    .q(\DFF_1265.Q )
  );
  al_dffl _11154_ (
    .clk(CK),
    .d(\DFF_1265.Q ),
    .q(\DFF_663.Q )
  );
  al_dffl _11155_ (
    .clk(CK),
    .d(\DFF_664.D ),
    .q(\DFF_664.Q )
  );
  al_dffl _11156_ (
    .clk(CK),
    .d(\DFF_665.D ),
    .q(\DFF_665.Q )
  );
  al_dffl _11157_ (
    .clk(CK),
    .d(\DFF_101.Q ),
    .q(\DFF_1352.Q )
  );
  al_dffl _11158_ (
    .clk(CK),
    .d(\DFF_1352.Q ),
    .q(\DFF_695.Q )
  );
  al_dffl _11159_ (
    .clk(CK),
    .d(\DFF_695.Q ),
    .q(\DFF_1262.Q )
  );
  al_dffl _11160_ (
    .clk(CK),
    .d(\DFF_1262.Q ),
    .q(\DFF_783.Q )
  );
  al_dffl _11161_ (
    .clk(CK),
    .d(\DFF_783.Q ),
    .q(\DFF_666.Q )
  );
  al_dffl _11162_ (
    .clk(CK),
    .d(\DFF_667.D ),
    .q(\DFF_667.Q )
  );
  al_dffl _11163_ (
    .clk(CK),
    .d(\DFF_668.D ),
    .q(\DFF_668.Q )
  );
  al_dffl _11164_ (
    .clk(CK),
    .d(\DFF_669.D ),
    .q(\DFF_669.Q )
  );
  al_dffl _11165_ (
    .clk(CK),
    .d(\DFF_670.D ),
    .q(\DFF_670.Q )
  );
  al_dffl _11166_ (
    .clk(CK),
    .d(\DFF_671.D ),
    .q(\DFF_671.Q )
  );
  al_dffl _11167_ (
    .clk(CK),
    .d(\DFF_672.D ),
    .q(\DFF_672.Q )
  );
  al_dffl _11168_ (
    .clk(CK),
    .d(\DFF_673.D ),
    .q(\DFF_673.Q )
  );
  al_dffl _11169_ (
    .clk(CK),
    .d(\DFF_674.D ),
    .q(\DFF_674.Q )
  );
  al_dffl _11170_ (
    .clk(CK),
    .d(\DFF_676.D ),
    .q(\DFF_676.Q )
  );
  al_dffl _11171_ (
    .clk(CK),
    .d(\DFF_677.D ),
    .q(\DFF_677.Q )
  );
  al_dffl _11172_ (
    .clk(CK),
    .d(\DFF_679.D ),
    .q(\DFF_679.Q )
  );
  al_dffl _11173_ (
    .clk(CK),
    .d(\DFF_680.D ),
    .q(\DFF_680.Q )
  );
  al_dffl _11174_ (
    .clk(CK),
    .d(\DFF_681.D ),
    .q(\DFF_681.Q )
  );
  al_dffl _11175_ (
    .clk(CK),
    .d(\DFF_682.D ),
    .q(\DFF_682.Q )
  );
  al_dffl _11176_ (
    .clk(CK),
    .d(\DFF_683.D ),
    .q(\DFF_683.Q )
  );
  al_dffl _11177_ (
    .clk(CK),
    .d(\DFF_684.D ),
    .q(\DFF_684.Q )
  );
  al_dffl _11178_ (
    .clk(CK),
    .d(\DFF_685.D ),
    .q(\DFF_685.Q )
  );
  al_dffl _11179_ (
    .clk(CK),
    .d(\DFF_686.D ),
    .q(\DFF_686.Q )
  );
  al_dffl _11180_ (
    .clk(CK),
    .d(\DFF_348.Q ),
    .q(\DFF_687.Q )
  );
  al_dffl _11181_ (
    .clk(CK),
    .d(\DFF_688.D ),
    .q(\DFF_688.Q )
  );
  al_dffl _11182_ (
    .clk(CK),
    .d(\DFF_689.D ),
    .q(\DFF_689.Q )
  );
  al_dffl _11183_ (
    .clk(CK),
    .d(\DFF_690.D ),
    .q(\DFF_690.Q )
  );
  al_dffl _11184_ (
    .clk(CK),
    .d(\DFF_691.D ),
    .q(\DFF_691.Q )
  );
  al_dffl _11185_ (
    .clk(CK),
    .d(\DFF_692.D ),
    .q(\DFF_692.Q )
  );
  al_dffl _11186_ (
    .clk(CK),
    .d(\DFF_693.D ),
    .q(\DFF_693.Q )
  );
  al_dffl _11187_ (
    .clk(CK),
    .d(\DFF_694.D ),
    .q(\DFF_694.Q )
  );
  al_dffl _11188_ (
    .clk(CK),
    .d(\DFF_696.D ),
    .q(\DFF_696.Q )
  );
  al_dffl _11189_ (
    .clk(CK),
    .d(\DFF_697.D ),
    .q(\DFF_697.Q )
  );
  al_dffl _11190_ (
    .clk(CK),
    .d(\DFF_600.Q ),
    .q(\DFF_698.Q )
  );
  al_dffl _11191_ (
    .clk(CK),
    .d(\DFF_699.D ),
    .q(\DFF_699.Q )
  );
  al_dffl _11192_ (
    .clk(CK),
    .d(\DFF_700.D ),
    .q(\DFF_700.Q )
  );
  al_dffl _11193_ (
    .clk(CK),
    .d(\DFF_701.D ),
    .q(\DFF_701.Q )
  );
  al_dffl _11194_ (
    .clk(CK),
    .d(\DFF_702.D ),
    .q(\DFF_702.Q )
  );
  al_dffl _11195_ (
    .clk(CK),
    .d(\DFF_703.D ),
    .q(\DFF_703.Q )
  );
  al_dffl _11196_ (
    .clk(CK),
    .d(\DFF_565.Q ),
    .q(\DFF_1224.Q )
  );
  al_dffl _11197_ (
    .clk(CK),
    .d(\DFF_1224.Q ),
    .q(\DFF_1416.Q )
  );
  al_dffl _11198_ (
    .clk(CK),
    .d(\DFF_1416.Q ),
    .q(\DFF_1049.Q )
  );
  al_dffl _11199_ (
    .clk(CK),
    .d(\DFF_1049.Q ),
    .q(\DFF_704.Q )
  );
  al_dffl _11200_ (
    .clk(CK),
    .d(\DFF_705.D ),
    .q(\DFF_705.Q )
  );
  al_dffl _11201_ (
    .clk(CK),
    .d(\DFF_706.D ),
    .q(\DFF_706.Q )
  );
  al_dffl _11202_ (
    .clk(CK),
    .d(\DFF_707.D ),
    .q(\DFF_707.Q )
  );
  al_dffl _11203_ (
    .clk(CK),
    .d(\DFF_708.D ),
    .q(\DFF_708.Q )
  );
  al_dffl _11204_ (
    .clk(CK),
    .d(\DFF_709.D ),
    .q(\DFF_709.Q )
  );
  al_dffl _11205_ (
    .clk(CK),
    .d(\DFF_710.D ),
    .q(\DFF_710.Q )
  );
  al_dffl _11206_ (
    .clk(CK),
    .d(\DFF_712.D ),
    .q(\DFF_712.Q )
  );
  al_dffl _11207_ (
    .clk(CK),
    .d(\DFF_713.D ),
    .q(\DFF_713.Q )
  );
  al_dffl _11208_ (
    .clk(CK),
    .d(\DFF_714.D ),
    .q(\DFF_714.Q )
  );
  al_dffl _11209_ (
    .clk(CK),
    .d(\DFF_715.D ),
    .q(\DFF_715.Q )
  );
  al_dffl _11210_ (
    .clk(CK),
    .d(\DFF_716.D ),
    .q(\DFF_716.Q )
  );
  al_dffl _11211_ (
    .clk(CK),
    .d(\DFF_717.D ),
    .q(\DFF_717.Q )
  );
  al_dffl _11212_ (
    .clk(CK),
    .d(\DFF_718.D ),
    .q(\DFF_718.Q )
  );
  al_dffl _11213_ (
    .clk(CK),
    .d(\DFF_719.D ),
    .q(\DFF_719.Q )
  );
  al_dffl _11214_ (
    .clk(CK),
    .d(\DFF_720.D ),
    .q(\DFF_720.Q )
  );
  al_dffl _11215_ (
    .clk(CK),
    .d(\DFF_721.D ),
    .q(\DFF_721.Q )
  );
  al_dffl _11216_ (
    .clk(CK),
    .d(\DFF_722.D ),
    .q(\DFF_722.Q )
  );
  al_dffl _11217_ (
    .clk(CK),
    .d(\DFF_723.D ),
    .q(\DFF_723.Q )
  );
  al_dffl _11218_ (
    .clk(CK),
    .d(\DFF_724.D ),
    .q(\DFF_724.Q )
  );
  al_dffl _11219_ (
    .clk(CK),
    .d(\DFF_725.D ),
    .q(\DFF_725.Q )
  );
  al_dffl _11220_ (
    .clk(CK),
    .d(\DFF_726.D ),
    .q(\DFF_726.Q )
  );
  al_dffl _11221_ (
    .clk(CK),
    .d(\DFF_727.D ),
    .q(\DFF_727.Q )
  );
  al_dffl _11222_ (
    .clk(CK),
    .d(\DFF_728.D ),
    .q(\DFF_728.Q )
  );
  al_dffl _11223_ (
    .clk(CK),
    .d(\DFF_729.D ),
    .q(\DFF_729.Q )
  );
  al_dffl _11224_ (
    .clk(CK),
    .d(\DFF_730.D ),
    .q(\DFF_730.Q )
  );
  al_dffl _11225_ (
    .clk(CK),
    .d(\DFF_731.D ),
    .q(\DFF_731.Q )
  );
  al_dffl _11226_ (
    .clk(CK),
    .d(\DFF_732.D ),
    .q(\DFF_732.Q )
  );
  al_dffl _11227_ (
    .clk(CK),
    .d(\DFF_733.D ),
    .q(\DFF_733.Q )
  );
  al_dffl _11228_ (
    .clk(CK),
    .d(\DFF_734.D ),
    .q(\DFF_734.Q )
  );
  al_dffl _11229_ (
    .clk(CK),
    .d(\DFF_735.D ),
    .q(\DFF_735.Q )
  );
  al_dffl _11230_ (
    .clk(CK),
    .d(\DFF_736.D ),
    .q(\DFF_736.Q )
  );
  al_dffl _11231_ (
    .clk(CK),
    .d(\DFF_738.D ),
    .q(\DFF_738.Q )
  );
  al_dffl _11232_ (
    .clk(CK),
    .d(\DFF_740.D ),
    .q(\DFF_740.Q )
  );
  al_dffl _11233_ (
    .clk(CK),
    .d(\DFF_741.D ),
    .q(\DFF_741.Q )
  );
  al_dffl _11234_ (
    .clk(CK),
    .d(\DFF_742.D ),
    .q(\DFF_742.Q )
  );
  al_dffl _11235_ (
    .clk(CK),
    .d(\DFF_743.D ),
    .q(\DFF_743.Q )
  );
  al_dffl _11236_ (
    .clk(CK),
    .d(\DFF_744.D ),
    .q(\DFF_744.Q )
  );
  al_dffl _11237_ (
    .clk(CK),
    .d(\DFF_745.D ),
    .q(\DFF_745.Q )
  );
  al_dffl _11238_ (
    .clk(CK),
    .d(\DFF_746.D ),
    .q(\DFF_746.Q )
  );
  al_dffl _11239_ (
    .clk(CK),
    .d(\DFF_747.D ),
    .q(\DFF_747.Q )
  );
  al_dffl _11240_ (
    .clk(CK),
    .d(\DFF_748.D ),
    .q(\DFF_748.Q )
  );
  al_dffl _11241_ (
    .clk(CK),
    .d(\DFF_749.D ),
    .q(\DFF_749.Q )
  );
  al_dffl _11242_ (
    .clk(CK),
    .d(\DFF_750.D ),
    .q(\DFF_750.Q )
  );
  al_dffl _11243_ (
    .clk(CK),
    .d(\DFF_751.D ),
    .q(\DFF_751.Q )
  );
  al_dffl _11244_ (
    .clk(CK),
    .d(\DFF_753.D ),
    .q(\DFF_753.Q )
  );
  al_dffl _11245_ (
    .clk(CK),
    .d(\DFF_754.D ),
    .q(\DFF_754.Q )
  );
  al_dffl _11246_ (
    .clk(CK),
    .d(\DFF_755.D ),
    .q(\DFF_755.Q )
  );
  al_dffl _11247_ (
    .clk(CK),
    .d(\DFF_756.D ),
    .q(\DFF_756.Q )
  );
  al_dffl _11248_ (
    .clk(CK),
    .d(\DFF_757.D ),
    .q(\DFF_757.Q )
  );
  al_dffl _11249_ (
    .clk(CK),
    .d(\DFF_758.D ),
    .q(\DFF_758.Q )
  );
  al_dffl _11250_ (
    .clk(CK),
    .d(\DFF_759.D ),
    .q(\DFF_759.Q )
  );
  al_dffl _11251_ (
    .clk(CK),
    .d(\DFF_760.D ),
    .q(\DFF_760.Q )
  );
  al_dffl _11252_ (
    .clk(CK),
    .d(\DFF_761.D ),
    .q(\DFF_761.Q )
  );
  al_dffl _11253_ (
    .clk(CK),
    .d(\DFF_762.D ),
    .q(\DFF_762.Q )
  );
  al_dffl _11254_ (
    .clk(CK),
    .d(\DFF_763.D ),
    .q(\DFF_763.Q )
  );
  al_dffl _11255_ (
    .clk(CK),
    .d(\DFF_380.Q ),
    .q(\DFF_764.Q )
  );
  al_dffl _11256_ (
    .clk(CK),
    .d(\DFF_766.D ),
    .q(\DFF_766.Q )
  );
  al_dffl _11257_ (
    .clk(CK),
    .d(\DFF_767.D ),
    .q(\DFF_767.Q )
  );
  al_dffl _11258_ (
    .clk(CK),
    .d(\DFF_768.D ),
    .q(\DFF_768.Q )
  );
  al_dffl _11259_ (
    .clk(CK),
    .d(\DFF_769.D ),
    .q(\DFF_769.Q )
  );
  al_dffl _11260_ (
    .clk(CK),
    .d(\DFF_770.D ),
    .q(\DFF_770.Q )
  );
  al_dffl _11261_ (
    .clk(CK),
    .d(\DFF_771.D ),
    .q(\DFF_771.Q )
  );
  al_dffl _11262_ (
    .clk(CK),
    .d(\DFF_772.D ),
    .q(\DFF_772.Q )
  );
  al_dffl _11263_ (
    .clk(CK),
    .d(\DFF_773.D ),
    .q(\DFF_773.Q )
  );
  al_dffl _11264_ (
    .clk(CK),
    .d(\DFF_774.D ),
    .q(\DFF_774.Q )
  );
  al_dffl _11265_ (
    .clk(CK),
    .d(\DFF_775.D ),
    .q(\DFF_775.Q )
  );
  al_dffl _11266_ (
    .clk(CK),
    .d(\DFF_776.D ),
    .q(\DFF_776.Q )
  );
  al_dffl _11267_ (
    .clk(CK),
    .d(\DFF_777.D ),
    .q(\DFF_777.Q )
  );
  al_dffl _11268_ (
    .clk(CK),
    .d(\DFF_778.D ),
    .q(\DFF_778.Q )
  );
  al_dffl _11269_ (
    .clk(CK),
    .d(\DFF_779.D ),
    .q(\DFF_779.Q )
  );
  al_dffl _11270_ (
    .clk(CK),
    .d(\DFF_163.Q ),
    .q(\DFF_971.Q )
  );
  al_dffl _11271_ (
    .clk(CK),
    .d(\DFF_971.Q ),
    .q(\DFF_836.Q )
  );
  al_dffl _11272_ (
    .clk(CK),
    .d(\DFF_836.Q ),
    .q(\DFF_780.Q )
  );
  al_dffl _11273_ (
    .clk(CK),
    .d(\DFF_781.D ),
    .q(\DFF_781.Q )
  );
  al_dffl _11274_ (
    .clk(CK),
    .d(\DFF_782.D ),
    .q(\DFF_782.Q )
  );
  al_dffl _11275_ (
    .clk(CK),
    .d(\DFF_784.D ),
    .q(\DFF_784.Q )
  );
  al_dffl _11276_ (
    .clk(CK),
    .d(\DFF_786.D ),
    .q(\DFF_786.Q )
  );
  al_dffl _11277_ (
    .clk(CK),
    .d(\DFF_787.D ),
    .q(\DFF_787.Q )
  );
  al_dffl _11278_ (
    .clk(CK),
    .d(\DFF_788.D ),
    .q(\DFF_788.Q )
  );
  al_dffl _11279_ (
    .clk(CK),
    .d(\DFF_789.D ),
    .q(\DFF_789.Q )
  );
  al_dffl _11280_ (
    .clk(CK),
    .d(\DFF_790.D ),
    .q(\DFF_790.Q )
  );
  al_dffl _11281_ (
    .clk(CK),
    .d(\DFF_185.Q ),
    .q(\DFF_791.Q )
  );
  al_dffl _11282_ (
    .clk(CK),
    .d(\DFF_792.D ),
    .q(\DFF_792.Q )
  );
  al_dffl _11283_ (
    .clk(CK),
    .d(\DFF_793.D ),
    .q(\DFF_793.Q )
  );
  al_dffl _11284_ (
    .clk(CK),
    .d(\DFF_794.D ),
    .q(\DFF_794.Q )
  );
  al_dffl _11285_ (
    .clk(CK),
    .d(\DFF_795.D ),
    .q(\DFF_795.Q )
  );
  al_dffl _11286_ (
    .clk(CK),
    .d(\DFF_796.D ),
    .q(\DFF_796.Q )
  );
  al_dffl _11287_ (
    .clk(CK),
    .d(\DFF_269.Q ),
    .q(\DFF_798.Q )
  );
  al_dffl _11288_ (
    .clk(CK),
    .d(\DFF_799.D ),
    .q(\DFF_799.Q )
  );
  al_dffl _11289_ (
    .clk(CK),
    .d(\DFF_800.D ),
    .q(\DFF_800.Q )
  );
  al_dffl _11290_ (
    .clk(CK),
    .d(\DFF_801.D ),
    .q(\DFF_801.Q )
  );
  al_dffl _11291_ (
    .clk(CK),
    .d(\DFF_802.D ),
    .q(\DFF_802.Q )
  );
  al_dffl _11292_ (
    .clk(CK),
    .d(\DFF_803.D ),
    .q(\DFF_803.Q )
  );
  al_dffl _11293_ (
    .clk(CK),
    .d(\DFF_804.D ),
    .q(\DFF_804.Q )
  );
  al_dffl _11294_ (
    .clk(CK),
    .d(\DFF_805.D ),
    .q(\DFF_805.Q )
  );
  al_dffl _11295_ (
    .clk(CK),
    .d(\DFF_807.D ),
    .q(\DFF_807.Q )
  );
  al_dffl _11296_ (
    .clk(CK),
    .d(\DFF_808.D ),
    .q(\DFF_808.Q )
  );
  al_dffl _11297_ (
    .clk(CK),
    .d(\DFF_809.D ),
    .q(\DFF_809.Q )
  );
  al_dffl _11298_ (
    .clk(CK),
    .d(\DFF_830.D ),
    .q(\DFF_830.Q )
  );
  al_dffl _11299_ (
    .clk(CK),
    .d(\DFF_830.Q ),
    .q(\DFF_810.Q )
  );
  al_dffl _11300_ (
    .clk(CK),
    .d(\DFF_811.D ),
    .q(\DFF_811.Q )
  );
  al_dffl _11301_ (
    .clk(CK),
    .d(\DFF_812.D ),
    .q(\DFF_812.Q )
  );
  al_dffl _11302_ (
    .clk(CK),
    .d(\DFF_813.D ),
    .q(\DFF_813.Q )
  );
  al_dffl _11303_ (
    .clk(CK),
    .d(\DFF_814.D ),
    .q(\DFF_814.Q )
  );
  al_dffl _11304_ (
    .clk(CK),
    .d(\DFF_815.D ),
    .q(\DFF_815.Q )
  );
  al_dffl _11305_ (
    .clk(CK),
    .d(\DFF_816.D ),
    .q(\DFF_816.Q )
  );
  al_dffl _11306_ (
    .clk(CK),
    .d(\DFF_1256.D ),
    .q(\DFF_1256.Q )
  );
  al_dffl _11307_ (
    .clk(CK),
    .d(\DFF_1256.Q ),
    .q(\DFF_817.Q )
  );
  al_dffl _11308_ (
    .clk(CK),
    .d(\DFF_818.D ),
    .q(\DFF_818.Q )
  );
  al_dffl _11309_ (
    .clk(CK),
    .d(\DFF_820.D ),
    .q(\DFF_820.Q )
  );
  al_dffl _11310_ (
    .clk(CK),
    .d(\DFF_821.D ),
    .q(\DFF_821.Q )
  );
  al_dffl _11311_ (
    .clk(CK),
    .d(\DFF_822.D ),
    .q(\DFF_822.Q )
  );
  al_dffl _11312_ (
    .clk(CK),
    .d(\DFF_823.D ),
    .q(\DFF_823.Q )
  );
  al_dffl _11313_ (
    .clk(CK),
    .d(\DFF_824.D ),
    .q(\DFF_824.Q )
  );
  al_dffl _11314_ (
    .clk(CK),
    .d(\DFF_825.D ),
    .q(\DFF_825.Q )
  );
  al_dffl _11315_ (
    .clk(CK),
    .d(\DFF_826.D ),
    .q(\DFF_826.Q )
  );
  al_dffl _11316_ (
    .clk(CK),
    .d(\DFF_827.D ),
    .q(\DFF_827.Q )
  );
  al_dffl _11317_ (
    .clk(CK),
    .d(\DFF_339.Q ),
    .q(\DFF_828.Q )
  );
  al_dffl _11318_ (
    .clk(CK),
    .d(\DFF_829.D ),
    .q(\DFF_829.Q )
  );
  al_dffl _11319_ (
    .clk(CK),
    .d(\DFF_832.D ),
    .q(\DFF_832.Q )
  );
  al_dffl _11320_ (
    .clk(CK),
    .d(\DFF_833.D ),
    .q(\DFF_833.Q )
  );
  al_dffl _11321_ (
    .clk(CK),
    .d(\DFF_834.D ),
    .q(\DFF_834.Q )
  );
  al_dffl _11322_ (
    .clk(CK),
    .d(\DFF_835.D ),
    .q(\DFF_835.Q )
  );
  al_dffl _11323_ (
    .clk(CK),
    .d(\DFF_837.D ),
    .q(\DFF_837.Q )
  );
  al_dffl _11324_ (
    .clk(CK),
    .d(\DFF_838.D ),
    .q(\DFF_838.Q )
  );
  al_dffl _11325_ (
    .clk(CK),
    .d(\DFF_839.D ),
    .q(\DFF_839.Q )
  );
  al_dffl _11326_ (
    .clk(CK),
    .d(\DFF_840.D ),
    .q(\DFF_840.Q )
  );
  al_dffl _11327_ (
    .clk(CK),
    .d(\DFF_841.D ),
    .q(\DFF_841.Q )
  );
  al_dffl _11328_ (
    .clk(CK),
    .d(\DFF_824.Q ),
    .q(\DFF_842.Q )
  );
  al_dffl _11329_ (
    .clk(CK),
    .d(\DFF_843.D ),
    .q(\DFF_843.Q )
  );
  al_dffl _11330_ (
    .clk(CK),
    .d(\DFF_844.D ),
    .q(\DFF_844.Q )
  );
  al_dffl _11331_ (
    .clk(CK),
    .d(\DFF_845.D ),
    .q(\DFF_845.Q )
  );
  al_dffl _11332_ (
    .clk(CK),
    .d(\DFF_846.D ),
    .q(\DFF_846.Q )
  );
  al_dffl _11333_ (
    .clk(CK),
    .d(\DFF_847.D ),
    .q(\DFF_847.Q )
  );
  al_dffl _11334_ (
    .clk(CK),
    .d(\DFF_849.D ),
    .q(\DFF_849.Q )
  );
  al_dffl _11335_ (
    .clk(CK),
    .d(\DFF_850.D ),
    .q(\DFF_850.Q )
  );
  al_dffl _11336_ (
    .clk(CK),
    .d(\DFF_851.D ),
    .q(\DFF_851.Q )
  );
  al_dffl _11337_ (
    .clk(CK),
    .d(\DFF_852.D ),
    .q(\DFF_852.Q )
  );
  al_dffl _11338_ (
    .clk(CK),
    .d(\DFF_853.D ),
    .q(\DFF_853.Q )
  );
  al_dffl _11339_ (
    .clk(CK),
    .d(\DFF_854.D ),
    .q(\DFF_854.Q )
  );
  al_dffl _11340_ (
    .clk(CK),
    .d(\DFF_855.D ),
    .q(\DFF_855.Q )
  );
  al_dffl _11341_ (
    .clk(CK),
    .d(\DFF_857.D ),
    .q(\DFF_857.Q )
  );
  al_dffl _11342_ (
    .clk(CK),
    .d(\DFF_858.D ),
    .q(\DFF_858.Q )
  );
  al_dffl _11343_ (
    .clk(CK),
    .d(\DFF_859.D ),
    .q(\DFF_859.Q )
  );
  al_dffl _11344_ (
    .clk(CK),
    .d(\DFF_860.D ),
    .q(\DFF_860.Q )
  );
  al_dffl _11345_ (
    .clk(CK),
    .d(\DFF_862.D ),
    .q(\DFF_862.Q )
  );
  al_dffl _11346_ (
    .clk(CK),
    .d(\DFF_863.D ),
    .q(\DFF_863.Q )
  );
  al_dffl _11347_ (
    .clk(CK),
    .d(\DFF_864.D ),
    .q(\DFF_864.Q )
  );
  al_dffl _11348_ (
    .clk(CK),
    .d(\DFF_865.D ),
    .q(\DFF_865.Q )
  );
  al_dffl _11349_ (
    .clk(CK),
    .d(\DFF_866.D ),
    .q(\DFF_866.Q )
  );
  al_dffl _11350_ (
    .clk(CK),
    .d(\DFF_867.D ),
    .q(\DFF_867.Q )
  );
  al_dffl _11351_ (
    .clk(CK),
    .d(\DFF_868.D ),
    .q(\DFF_868.Q )
  );
  al_dffl _11352_ (
    .clk(CK),
    .d(\DFF_869.D ),
    .q(\DFF_869.Q )
  );
  al_dffl _11353_ (
    .clk(CK),
    .d(\DFF_870.D ),
    .q(\DFF_870.Q )
  );
  al_dffl _11354_ (
    .clk(CK),
    .d(\DFF_871.D ),
    .q(\DFF_871.Q )
  );
  al_dffl _11355_ (
    .clk(CK),
    .d(\DFF_872.D ),
    .q(\DFF_872.Q )
  );
  al_dffl _11356_ (
    .clk(CK),
    .d(\DFF_874.D ),
    .q(\DFF_874.Q )
  );
  al_dffl _11357_ (
    .clk(CK),
    .d(\DFF_875.D ),
    .q(\DFF_875.Q )
  );
  al_dffl _11358_ (
    .clk(CK),
    .d(\DFF_876.D ),
    .q(\DFF_876.Q )
  );
  al_dffl _11359_ (
    .clk(CK),
    .d(\DFF_877.D ),
    .q(\DFF_877.Q )
  );
  al_dffl _11360_ (
    .clk(CK),
    .d(\DFF_878.D ),
    .q(\DFF_878.Q )
  );
  al_dffl _11361_ (
    .clk(CK),
    .d(\DFF_879.D ),
    .q(\DFF_879.Q )
  );
  al_dffl _11362_ (
    .clk(CK),
    .d(\DFF_880.D ),
    .q(\DFF_880.Q )
  );
  al_dffl _11363_ (
    .clk(CK),
    .d(\DFF_881.D ),
    .q(\DFF_881.Q )
  );
  al_dffl _11364_ (
    .clk(CK),
    .d(\DFF_882.D ),
    .q(\DFF_882.Q )
  );
  al_dffl _11365_ (
    .clk(CK),
    .d(\DFF_883.D ),
    .q(\DFF_883.Q )
  );
  al_dffl _11366_ (
    .clk(CK),
    .d(\DFF_884.D ),
    .q(\DFF_884.Q )
  );
  al_dffl _11367_ (
    .clk(CK),
    .d(\DFF_886.D ),
    .q(\DFF_886.Q )
  );
  al_dffl _11368_ (
    .clk(CK),
    .d(\DFF_887.D ),
    .q(\DFF_887.Q )
  );
  al_dffl _11369_ (
    .clk(CK),
    .d(\DFF_888.D ),
    .q(\DFF_888.Q )
  );
  al_dffl _11370_ (
    .clk(CK),
    .d(\DFF_889.D ),
    .q(\DFF_889.Q )
  );
  al_dffl _11371_ (
    .clk(CK),
    .d(\DFF_890.D ),
    .q(\DFF_890.Q )
  );
  al_dffl _11372_ (
    .clk(CK),
    .d(\DFF_891.D ),
    .q(\DFF_891.Q )
  );
  al_dffl _11373_ (
    .clk(CK),
    .d(\DFF_892.D ),
    .q(\DFF_892.Q )
  );
  al_dffl _11374_ (
    .clk(CK),
    .d(\DFF_893.D ),
    .q(\DFF_893.Q )
  );
  al_dffl _11375_ (
    .clk(CK),
    .d(\DFF_894.D ),
    .q(\DFF_894.Q )
  );
  al_dffl _11376_ (
    .clk(CK),
    .d(\DFF_895.D ),
    .q(\DFF_895.Q )
  );
  al_dffl _11377_ (
    .clk(CK),
    .d(\DFF_896.D ),
    .q(\DFF_896.Q )
  );
  al_dffl _11378_ (
    .clk(CK),
    .d(\DFF_897.D ),
    .q(\DFF_897.Q )
  );
  al_dffl _11379_ (
    .clk(CK),
    .d(\DFF_899.D ),
    .q(\DFF_899.Q )
  );
  al_dffl _11380_ (
    .clk(CK),
    .d(\DFF_900.D ),
    .q(\DFF_900.Q )
  );
  al_dffl _11381_ (
    .clk(CK),
    .d(\DFF_901.D ),
    .q(\DFF_901.Q )
  );
  al_dffl _11382_ (
    .clk(CK),
    .d(\DFF_902.D ),
    .q(\DFF_902.Q )
  );
  al_dffl _11383_ (
    .clk(CK),
    .d(\DFF_903.D ),
    .q(\DFF_903.Q )
  );
  al_dffl _11384_ (
    .clk(CK),
    .d(\DFF_904.D ),
    .q(\DFF_904.Q )
  );
  al_dffl _11385_ (
    .clk(CK),
    .d(\DFF_907.D ),
    .q(\DFF_907.Q )
  );
  al_dffl _11386_ (
    .clk(CK),
    .d(\DFF_908.D ),
    .q(\DFF_908.Q )
  );
  al_dffl _11387_ (
    .clk(CK),
    .d(\DFF_910.D ),
    .q(\DFF_910.Q )
  );
  al_dffl _11388_ (
    .clk(CK),
    .d(\DFF_911.D ),
    .q(\DFF_911.Q )
  );
  al_dffl _11389_ (
    .clk(CK),
    .d(\DFF_912.D ),
    .q(\DFF_912.Q )
  );
  al_dffl _11390_ (
    .clk(CK),
    .d(\DFF_913.D ),
    .q(\DFF_913.Q )
  );
  al_dffl _11391_ (
    .clk(CK),
    .d(\DFF_914.D ),
    .q(\DFF_914.Q )
  );
  al_dffl _11392_ (
    .clk(CK),
    .d(\DFF_915.D ),
    .q(\DFF_915.Q )
  );
  al_dffl _11393_ (
    .clk(CK),
    .d(\DFF_916.D ),
    .q(\DFF_916.Q )
  );
  al_dffl _11394_ (
    .clk(CK),
    .d(\DFF_917.D ),
    .q(\DFF_917.Q )
  );
  al_dffl _11395_ (
    .clk(CK),
    .d(\DFF_918.D ),
    .q(\DFF_918.Q )
  );
  al_dffl _11396_ (
    .clk(CK),
    .d(\DFF_919.D ),
    .q(\DFF_919.Q )
  );
  al_dffl _11397_ (
    .clk(CK),
    .d(\DFF_920.D ),
    .q(\DFF_920.Q )
  );
  al_dffl _11398_ (
    .clk(CK),
    .d(\DFF_921.D ),
    .q(\DFF_921.Q )
  );
  al_dffl _11399_ (
    .clk(CK),
    .d(\DFF_922.D ),
    .q(\DFF_922.Q )
  );
  al_dffl _11400_ (
    .clk(CK),
    .d(\DFF_923.D ),
    .q(\DFF_923.Q )
  );
  al_dffl _11401_ (
    .clk(CK),
    .d(\DFF_924.D ),
    .q(\DFF_924.Q )
  );
  al_dffl _11402_ (
    .clk(CK),
    .d(\DFF_925.D ),
    .q(\DFF_925.Q )
  );
  al_dffl _11403_ (
    .clk(CK),
    .d(\DFF_926.D ),
    .q(\DFF_926.Q )
  );
  al_dffl _11404_ (
    .clk(CK),
    .d(\DFF_928.D ),
    .q(\DFF_928.Q )
  );
  al_dffl _11405_ (
    .clk(CK),
    .d(\DFF_929.D ),
    .q(\DFF_929.Q )
  );
  al_dffl _11406_ (
    .clk(CK),
    .d(\DFF_930.D ),
    .q(\DFF_930.Q )
  );
  al_dffl _11407_ (
    .clk(CK),
    .d(\DFF_931.D ),
    .q(\DFF_931.Q )
  );
  al_dffl _11408_ (
    .clk(CK),
    .d(\DFF_932.D ),
    .q(\DFF_932.Q )
  );
  al_dffl _11409_ (
    .clk(CK),
    .d(\DFF_933.D ),
    .q(\DFF_933.Q )
  );
  al_dffl _11410_ (
    .clk(CK),
    .d(\DFF_934.D ),
    .q(\DFF_934.Q )
  );
  al_dffl _11411_ (
    .clk(CK),
    .d(\DFF_935.D ),
    .q(\DFF_935.Q )
  );
  al_dffl _11412_ (
    .clk(CK),
    .d(\DFF_936.D ),
    .q(\DFF_936.Q )
  );
  al_dffl _11413_ (
    .clk(CK),
    .d(\DFF_938.D ),
    .q(\DFF_938.Q )
  );
  al_dffl _11414_ (
    .clk(CK),
    .d(\DFF_939.D ),
    .q(\DFF_939.Q )
  );
  al_dffl _11415_ (
    .clk(CK),
    .d(\DFF_940.D ),
    .q(\DFF_940.Q )
  );
  al_dffl _11416_ (
    .clk(CK),
    .d(\DFF_941.D ),
    .q(\DFF_941.Q )
  );
  al_dffl _11417_ (
    .clk(CK),
    .d(\DFF_943.D ),
    .q(\DFF_943.Q )
  );
  al_dffl _11418_ (
    .clk(CK),
    .d(\DFF_945.D ),
    .q(\DFF_945.Q )
  );
  al_dffl _11419_ (
    .clk(CK),
    .d(\DFF_946.D ),
    .q(\DFF_946.Q )
  );
  al_dffl _11420_ (
    .clk(CK),
    .d(\DFF_947.D ),
    .q(\DFF_947.Q )
  );
  al_dffl _11421_ (
    .clk(CK),
    .d(\DFF_948.D ),
    .q(\DFF_948.Q )
  );
  al_dffl _11422_ (
    .clk(CK),
    .d(\DFF_949.D ),
    .q(\DFF_949.Q )
  );
  al_dffl _11423_ (
    .clk(CK),
    .d(\DFF_950.D ),
    .q(\DFF_950.Q )
  );
  al_dffl _11424_ (
    .clk(CK),
    .d(\DFF_951.D ),
    .q(\DFF_951.Q )
  );
  al_dffl _11425_ (
    .clk(CK),
    .d(\DFF_952.D ),
    .q(\DFF_952.Q )
  );
  al_dffl _11426_ (
    .clk(CK),
    .d(\DFF_953.D ),
    .q(\DFF_953.Q )
  );
  al_dffl _11427_ (
    .clk(CK),
    .d(\DFF_954.D ),
    .q(\DFF_954.Q )
  );
  al_dffl _11428_ (
    .clk(CK),
    .d(\DFF_955.D ),
    .q(\DFF_955.Q )
  );
  al_dffl _11429_ (
    .clk(CK),
    .d(\DFF_956.D ),
    .q(\DFF_956.Q )
  );
  al_dffl _11430_ (
    .clk(CK),
    .d(\DFF_957.D ),
    .q(\DFF_957.Q )
  );
  al_dffl _11431_ (
    .clk(CK),
    .d(\DFF_958.D ),
    .q(\DFF_958.Q )
  );
  al_dffl _11432_ (
    .clk(CK),
    .d(\DFF_959.D ),
    .q(\DFF_959.Q )
  );
  al_dffl _11433_ (
    .clk(CK),
    .d(\DFF_960.D ),
    .q(\DFF_960.Q )
  );
  al_dffl _11434_ (
    .clk(CK),
    .d(\DFF_961.D ),
    .q(\DFF_961.Q )
  );
  al_dffl _11435_ (
    .clk(CK),
    .d(\DFF_962.D ),
    .q(\DFF_962.Q )
  );
  al_dffl _11436_ (
    .clk(CK),
    .d(\DFF_963.D ),
    .q(\DFF_963.Q )
  );
  al_dffl _11437_ (
    .clk(CK),
    .d(\DFF_964.D ),
    .q(\DFF_964.Q )
  );
  al_dffl _11438_ (
    .clk(CK),
    .d(\DFF_965.D ),
    .q(\DFF_965.Q )
  );
  al_dffl _11439_ (
    .clk(CK),
    .d(\DFF_966.D ),
    .q(\DFF_966.Q )
  );
  al_dffl _11440_ (
    .clk(CK),
    .d(\DFF_967.D ),
    .q(\DFF_967.Q )
  );
  al_dffl _11441_ (
    .clk(CK),
    .d(\DFF_968.D ),
    .q(\DFF_968.Q )
  );
  al_dffl _11442_ (
    .clk(CK),
    .d(\DFF_969.D ),
    .q(\DFF_969.Q )
  );
  al_dffl _11443_ (
    .clk(CK),
    .d(\DFF_972.D ),
    .q(\DFF_972.Q )
  );
  al_dffl _11444_ (
    .clk(CK),
    .d(\DFF_973.D ),
    .q(\DFF_973.Q )
  );
  al_dffl _11445_ (
    .clk(CK),
    .d(\DFF_974.D ),
    .q(\DFF_974.Q )
  );
  al_dffl _11446_ (
    .clk(CK),
    .d(\DFF_975.D ),
    .q(\DFF_975.Q )
  );
  al_dffl _11447_ (
    .clk(CK),
    .d(\DFF_976.D ),
    .q(\DFF_976.Q )
  );
  al_dffl _11448_ (
    .clk(CK),
    .d(\DFF_977.D ),
    .q(\DFF_977.Q )
  );
  al_dffl _11449_ (
    .clk(CK),
    .d(\DFF_978.D ),
    .q(\DFF_978.Q )
  );
  al_dffl _11450_ (
    .clk(CK),
    .d(\DFF_979.D ),
    .q(\DFF_979.Q )
  );
  al_dffl _11451_ (
    .clk(CK),
    .d(\DFF_980.D ),
    .q(\DFF_980.Q )
  );
  al_dffl _11452_ (
    .clk(CK),
    .d(\DFF_672.Q ),
    .q(\DFF_981.Q )
  );
  al_dffl _11453_ (
    .clk(CK),
    .d(\DFF_982.D ),
    .q(\DFF_982.Q )
  );
  al_dffl _11454_ (
    .clk(CK),
    .d(\DFF_983.D ),
    .q(\DFF_983.Q )
  );
  al_dffl _11455_ (
    .clk(CK),
    .d(\DFF_984.D ),
    .q(\DFF_984.Q )
  );
  al_dffl _11456_ (
    .clk(CK),
    .d(\DFF_985.D ),
    .q(\DFF_985.Q )
  );
  al_dffl _11457_ (
    .clk(CK),
    .d(\DFF_986.D ),
    .q(\DFF_986.Q )
  );
  al_dffl _11458_ (
    .clk(CK),
    .d(\DFF_987.D ),
    .q(\DFF_987.Q )
  );
  al_dffl _11459_ (
    .clk(CK),
    .d(\DFF_988.D ),
    .q(\DFF_988.Q )
  );
  al_dffl _11460_ (
    .clk(CK),
    .d(\DFF_989.D ),
    .q(\DFF_989.Q )
  );
  al_dffl _11461_ (
    .clk(CK),
    .d(\DFF_327.Q ),
    .q(\DFF_990.Q )
  );
  al_dffl _11462_ (
    .clk(CK),
    .d(\DFF_1345.Q ),
    .q(\DFF_991.Q )
  );
  al_dffl _11463_ (
    .clk(CK),
    .d(\DFF_993.D ),
    .q(\DFF_993.Q )
  );
  al_dffl _11464_ (
    .clk(CK),
    .d(\DFF_994.D ),
    .q(\DFF_994.Q )
  );
  al_dffl _11465_ (
    .clk(CK),
    .d(\DFF_662.Q ),
    .q(\DFF_1219.Q )
  );
  al_dffl _11466_ (
    .clk(CK),
    .d(\DFF_1219.Q ),
    .q(\DFF_995.Q )
  );
  al_dffl _11467_ (
    .clk(CK),
    .d(\DFF_996.D ),
    .q(\DFF_996.Q )
  );
  al_dffl _11468_ (
    .clk(CK),
    .d(\DFF_178.Q ),
    .q(\DFF_997.Q )
  );
  al_dffl _11469_ (
    .clk(CK),
    .d(\DFF_998.D ),
    .q(\DFF_998.Q )
  );
  al_dffl _11470_ (
    .clk(CK),
    .d(\DFF_999.D ),
    .q(\DFF_999.Q )
  );
  al_dffl _11471_ (
    .clk(CK),
    .d(\DFF_1000.D ),
    .q(\DFF_1000.Q )
  );
  al_dffl _11472_ (
    .clk(CK),
    .d(\DFF_1073.D ),
    .q(\DFF_1073.Q )
  );
  al_dffl _11473_ (
    .clk(CK),
    .d(\DFF_1073.Q ),
    .q(\DFF_1002.Q )
  );
  al_dffl _11474_ (
    .clk(CK),
    .d(\DFF_764.Q ),
    .q(\DFF_1003.Q )
  );
  al_dffl _11475_ (
    .clk(CK),
    .d(\DFF_1004.D ),
    .q(\DFF_1004.Q )
  );
  al_dffl _11476_ (
    .clk(CK),
    .d(\DFF_1005.D ),
    .q(\DFF_1005.Q )
  );
  al_dffl _11477_ (
    .clk(CK),
    .d(\DFF_1006.D ),
    .q(\DFF_1006.Q )
  );
  al_dffl _11478_ (
    .clk(CK),
    .d(\DFF_1007.D ),
    .q(\DFF_1007.Q )
  );
  al_dffl _11479_ (
    .clk(CK),
    .d(\DFF_1008.D ),
    .q(\DFF_1008.Q )
  );
  al_dffl _11480_ (
    .clk(CK),
    .d(\DFF_1009.D ),
    .q(\DFF_1009.Q )
  );
  al_dffl _11481_ (
    .clk(CK),
    .d(\DFF_1010.D ),
    .q(\DFF_1010.Q )
  );
  al_dffl _11482_ (
    .clk(CK),
    .d(\DFF_1011.D ),
    .q(\DFF_1011.Q )
  );
  al_dffl _11483_ (
    .clk(CK),
    .d(\DFF_1012.D ),
    .q(\DFF_1012.Q )
  );
  al_dffl _11484_ (
    .clk(CK),
    .d(\DFF_1013.D ),
    .q(\DFF_1013.Q )
  );
  al_dffl _11485_ (
    .clk(CK),
    .d(\DFF_686.Q ),
    .q(\DFF_1014.Q )
  );
  al_dffl _11486_ (
    .clk(CK),
    .d(\DFF_1015.D ),
    .q(\DFF_1015.Q )
  );
  al_dffl _11487_ (
    .clk(CK),
    .d(\DFF_1016.D ),
    .q(\DFF_1016.Q )
  );
  al_dffl _11488_ (
    .clk(CK),
    .d(\DFF_1017.D ),
    .q(\DFF_1017.Q )
  );
  al_dffl _11489_ (
    .clk(CK),
    .d(\DFF_1018.D ),
    .q(\DFF_1018.Q )
  );
  al_dffl _11490_ (
    .clk(CK),
    .d(\DFF_1019.D ),
    .q(\DFF_1019.Q )
  );
  al_dffl _11491_ (
    .clk(CK),
    .d(\DFF_1020.D ),
    .q(\DFF_1020.Q )
  );
  al_dffl _11492_ (
    .clk(CK),
    .d(\DFF_1021.D ),
    .q(\DFF_1021.Q )
  );
  al_dffl _11493_ (
    .clk(CK),
    .d(\DFF_1022.D ),
    .q(\DFF_1022.Q )
  );
  al_dffl _11494_ (
    .clk(CK),
    .d(\DFF_780.Q ),
    .q(\DFF_1023.Q )
  );
  al_dffl _11495_ (
    .clk(CK),
    .d(\DFF_1024.D ),
    .q(\DFF_1024.Q )
  );
  al_dffl _11496_ (
    .clk(CK),
    .d(\DFF_1025.D ),
    .q(\DFF_1025.Q )
  );
  al_dffl _11497_ (
    .clk(CK),
    .d(\DFF_1026.D ),
    .q(\DFF_1026.Q )
  );
  al_dffl _11498_ (
    .clk(CK),
    .d(\DFF_1027.D ),
    .q(\DFF_1027.Q )
  );
  al_dffl _11499_ (
    .clk(CK),
    .d(\DFF_1028.D ),
    .q(\DFF_1028.Q )
  );
  al_dffl _11500_ (
    .clk(CK),
    .d(\DFF_1029.D ),
    .q(\DFF_1029.Q )
  );
  al_dffl _11501_ (
    .clk(CK),
    .d(\DFF_1030.D ),
    .q(\DFF_1030.Q )
  );
  al_dffl _11502_ (
    .clk(CK),
    .d(\DFF_1031.D ),
    .q(\DFF_1031.Q )
  );
  al_dffl _11503_ (
    .clk(CK),
    .d(\DFF_1032.D ),
    .q(\DFF_1032.Q )
  );
  al_dffl _11504_ (
    .clk(CK),
    .d(\DFF_1033.D ),
    .q(\DFF_1033.Q )
  );
  al_dffl _11505_ (
    .clk(CK),
    .d(\DFF_1034.D ),
    .q(\DFF_1034.Q )
  );
  al_dffl _11506_ (
    .clk(CK),
    .d(\DFF_1035.D ),
    .q(\DFF_1035.Q )
  );
  al_dffl _11507_ (
    .clk(CK),
    .d(\DFF_1036.D ),
    .q(\DFF_1036.Q )
  );
  al_dffl _11508_ (
    .clk(CK),
    .d(\DFF_1037.D ),
    .q(\DFF_1037.Q )
  );
  al_dffl _11509_ (
    .clk(CK),
    .d(\DFF_1039.D ),
    .q(\DFF_1039.Q )
  );
  al_dffl _11510_ (
    .clk(CK),
    .d(\DFF_1040.D ),
    .q(\DFF_1040.Q )
  );
  al_dffl _11511_ (
    .clk(CK),
    .d(\DFF_1041.D ),
    .q(\DFF_1041.Q )
  );
  al_dffl _11512_ (
    .clk(CK),
    .d(\DFF_1042.D ),
    .q(\DFF_1042.Q )
  );
  al_dffl _11513_ (
    .clk(CK),
    .d(\DFF_1027.Q ),
    .q(\DFF_1043.Q )
  );
  al_dffl _11514_ (
    .clk(CK),
    .d(\DFF_1044.D ),
    .q(\DFF_1044.Q )
  );
  al_dffl _11515_ (
    .clk(CK),
    .d(\DFF_1045.D ),
    .q(\DFF_1045.Q )
  );
  al_dffl _11516_ (
    .clk(CK),
    .d(\DFF_1046.D ),
    .q(\DFF_1046.Q )
  );
  al_dffl _11517_ (
    .clk(CK),
    .d(\DFF_1047.D ),
    .q(\DFF_1047.Q )
  );
  al_dffl _11518_ (
    .clk(CK),
    .d(\DFF_1048.D ),
    .q(\DFF_1048.Q )
  );
  al_dffl _11519_ (
    .clk(CK),
    .d(\DFF_1050.D ),
    .q(\DFF_1050.Q )
  );
  al_dffl _11520_ (
    .clk(CK),
    .d(\DFF_1051.D ),
    .q(\DFF_1051.Q )
  );
  al_dffl _11521_ (
    .clk(CK),
    .d(\DFF_1052.D ),
    .q(\DFF_1052.Q )
  );
  al_dffl _11522_ (
    .clk(CK),
    .d(\DFF_1053.D ),
    .q(\DFF_1053.Q )
  );
  al_dffl _11523_ (
    .clk(CK),
    .d(\DFF_1054.D ),
    .q(\DFF_1054.Q )
  );
  al_dffl _11524_ (
    .clk(CK),
    .d(\DFF_1055.D ),
    .q(\DFF_1055.Q )
  );
  al_dffl _11525_ (
    .clk(CK),
    .d(\DFF_1056.D ),
    .q(\DFF_1056.Q )
  );
  al_dffl _11526_ (
    .clk(CK),
    .d(\DFF_1057.D ),
    .q(\DFF_1057.Q )
  );
  al_dffl _11527_ (
    .clk(CK),
    .d(\DFF_1058.D ),
    .q(\DFF_1058.Q )
  );
  al_dffl _11528_ (
    .clk(CK),
    .d(\DFF_1059.D ),
    .q(\DFF_1059.Q )
  );
  al_dffl _11529_ (
    .clk(CK),
    .d(\DFF_1060.D ),
    .q(\DFF_1060.Q )
  );
  al_dffl _11530_ (
    .clk(CK),
    .d(\DFF_612.Q ),
    .q(\DFF_1061.Q )
  );
  al_dffl _11531_ (
    .clk(CK),
    .d(\DFF_1062.D ),
    .q(\DFF_1062.Q )
  );
  al_dffl _11532_ (
    .clk(CK),
    .d(\DFF_1063.D ),
    .q(\DFF_1063.Q )
  );
  al_dffl _11533_ (
    .clk(CK),
    .d(\DFF_1064.D ),
    .q(\DFF_1064.Q )
  );
  al_dffl _11534_ (
    .clk(CK),
    .d(\DFF_1065.D ),
    .q(\DFF_1065.Q )
  );
  al_dffl _11535_ (
    .clk(CK),
    .d(\DFF_1066.D ),
    .q(\DFF_1066.Q )
  );
  al_dffl _11536_ (
    .clk(CK),
    .d(\DFF_1067.D ),
    .q(\DFF_1067.Q )
  );
  al_dffl _11537_ (
    .clk(CK),
    .d(\DFF_1068.D ),
    .q(\DFF_1068.Q )
  );
  al_dffl _11538_ (
    .clk(CK),
    .d(\DFF_1069.D ),
    .q(\DFF_1069.Q )
  );
  al_dffl _11539_ (
    .clk(CK),
    .d(\DFF_1070.D ),
    .q(\DFF_1070.Q )
  );
  al_dffl _11540_ (
    .clk(CK),
    .d(\DFF_1071.D ),
    .q(\DFF_1071.Q )
  );
  al_dffl _11541_ (
    .clk(CK),
    .d(\DFF_1074.D ),
    .q(\DFF_1074.Q )
  );
  al_dffl _11542_ (
    .clk(CK),
    .d(\DFF_1075.D ),
    .q(\DFF_1075.Q )
  );
  al_dffl _11543_ (
    .clk(CK),
    .d(\DFF_1076.D ),
    .q(\DFF_1076.Q )
  );
  al_dffl _11544_ (
    .clk(CK),
    .d(\DFF_1077.D ),
    .q(\DFF_1077.Q )
  );
  al_dffl _11545_ (
    .clk(CK),
    .d(\DFF_1078.D ),
    .q(\DFF_1078.Q )
  );
  al_dffl _11546_ (
    .clk(CK),
    .d(\DFF_1079.D ),
    .q(\DFF_1079.Q )
  );
  al_dffl _11547_ (
    .clk(CK),
    .d(\DFF_1080.D ),
    .q(\DFF_1080.Q )
  );
  al_dffl _11548_ (
    .clk(CK),
    .d(\DFF_1082.D ),
    .q(\DFF_1082.Q )
  );
  al_dffl _11549_ (
    .clk(CK),
    .d(\DFF_1083.D ),
    .q(\DFF_1083.Q )
  );
  al_dffl _11550_ (
    .clk(CK),
    .d(\DFF_1084.D ),
    .q(\DFF_1084.Q )
  );
  al_dffl _11551_ (
    .clk(CK),
    .d(\DFF_1085.D ),
    .q(\DFF_1085.Q )
  );
  al_dffl _11552_ (
    .clk(CK),
    .d(\DFF_1086.D ),
    .q(\DFF_1086.Q )
  );
  al_dffl _11553_ (
    .clk(CK),
    .d(\DFF_1089.D ),
    .q(\DFF_1089.Q )
  );
  al_dffl _11554_ (
    .clk(CK),
    .d(\DFF_1090.D ),
    .q(\DFF_1090.Q )
  );
  al_dffl _11555_ (
    .clk(CK),
    .d(\DFF_1091.D ),
    .q(\DFF_1091.Q )
  );
  al_dffl _11556_ (
    .clk(CK),
    .d(\DFF_1092.D ),
    .q(\DFF_1092.Q )
  );
  al_dffl _11557_ (
    .clk(CK),
    .d(\DFF_1093.D ),
    .q(\DFF_1093.Q )
  );
  al_dffl _11558_ (
    .clk(CK),
    .d(\DFF_1094.D ),
    .q(\DFF_1094.Q )
  );
  al_dffl _11559_ (
    .clk(CK),
    .d(\DFF_1095.D ),
    .q(\DFF_1095.Q )
  );
  al_dffl _11560_ (
    .clk(CK),
    .d(\DFF_1096.D ),
    .q(\DFF_1096.Q )
  );
  al_dffl _11561_ (
    .clk(CK),
    .d(\DFF_1097.D ),
    .q(\DFF_1097.Q )
  );
  al_dffl _11562_ (
    .clk(CK),
    .d(\DFF_1098.D ),
    .q(\DFF_1098.Q )
  );
  al_dffl _11563_ (
    .clk(CK),
    .d(\DFF_1099.D ),
    .q(\DFF_1099.Q )
  );
  al_dffl _11564_ (
    .clk(CK),
    .d(\DFF_981.Q ),
    .q(\DFF_1100.Q )
  );
  al_dffl _11565_ (
    .clk(CK),
    .d(\DFF_1101.D ),
    .q(\DFF_1101.Q )
  );
  al_dffl _11566_ (
    .clk(CK),
    .d(\DFF_1103.D ),
    .q(\DFF_1103.Q )
  );
  al_dffl _11567_ (
    .clk(CK),
    .d(\DFF_1104.D ),
    .q(\DFF_1104.Q )
  );
  al_dffl _11568_ (
    .clk(CK),
    .d(\DFF_1105.D ),
    .q(\DFF_1105.Q )
  );
  al_dffl _11569_ (
    .clk(CK),
    .d(\DFF_1107.D ),
    .q(\DFF_1107.Q )
  );
  al_dffl _11570_ (
    .clk(CK),
    .d(\DFF_1108.D ),
    .q(\DFF_1108.Q )
  );
  al_dffl _11571_ (
    .clk(CK),
    .d(\DFF_1109.D ),
    .q(\DFF_1109.Q )
  );
  al_dffl _11572_ (
    .clk(CK),
    .d(\DFF_1111.D ),
    .q(\DFF_1111.Q )
  );
  al_dffl _11573_ (
    .clk(CK),
    .d(\DFF_1112.D ),
    .q(\DFF_1112.Q )
  );
  al_dffl _11574_ (
    .clk(CK),
    .d(\DFF_1113.D ),
    .q(\DFF_1113.Q )
  );
  al_dffl _11575_ (
    .clk(CK),
    .d(\DFF_1114.D ),
    .q(\DFF_1114.Q )
  );
  al_dffl _11576_ (
    .clk(CK),
    .d(\DFF_1115.D ),
    .q(\DFF_1115.Q )
  );
  al_dffl _11577_ (
    .clk(CK),
    .d(\DFF_1116.D ),
    .q(\DFF_1116.Q )
  );
  al_dffl _11578_ (
    .clk(CK),
    .d(\DFF_1117.D ),
    .q(\DFF_1117.Q )
  );
  al_dffl _11579_ (
    .clk(CK),
    .d(\DFF_997.Q ),
    .q(\DFF_1118.Q )
  );
  al_dffl _11580_ (
    .clk(CK),
    .d(\DFF_1120.D ),
    .q(\DFF_1120.Q )
  );
  al_dffl _11581_ (
    .clk(CK),
    .d(\DFF_1121.D ),
    .q(\DFF_1121.Q )
  );
  al_dffl _11582_ (
    .clk(CK),
    .d(\DFF_1123.D ),
    .q(\DFF_1123.Q )
  );
  al_dffl _11583_ (
    .clk(CK),
    .d(\DFF_1124.D ),
    .q(\DFF_1124.Q )
  );
  al_dffl _11584_ (
    .clk(CK),
    .d(\DFF_1125.D ),
    .q(\DFF_1125.Q )
  );
  al_dffl _11585_ (
    .clk(CK),
    .d(\DFF_1126.D ),
    .q(\DFF_1126.Q )
  );
  al_dffl _11586_ (
    .clk(CK),
    .d(\DFF_1127.D ),
    .q(\DFF_1127.Q )
  );
  al_dffl _11587_ (
    .clk(CK),
    .d(\DFF_1128.D ),
    .q(\DFF_1128.Q )
  );
  al_dffl _11588_ (
    .clk(CK),
    .d(\DFF_1129.D ),
    .q(\DFF_1129.Q )
  );
  al_dffl _11589_ (
    .clk(CK),
    .d(\DFF_1130.D ),
    .q(\DFF_1130.Q )
  );
  al_dffl _11590_ (
    .clk(CK),
    .d(\DFF_1131.D ),
    .q(\DFF_1131.Q )
  );
  al_dffl _11591_ (
    .clk(CK),
    .d(\DFF_1132.D ),
    .q(\DFF_1132.Q )
  );
  al_dffl _11592_ (
    .clk(CK),
    .d(\DFF_1133.D ),
    .q(\DFF_1133.Q )
  );
  al_dffl _11593_ (
    .clk(CK),
    .d(\DFF_1134.D ),
    .q(\DFF_1134.Q )
  );
  al_dffl _11594_ (
    .clk(CK),
    .d(\DFF_1135.D ),
    .q(\DFF_1135.Q )
  );
  al_dffl _11595_ (
    .clk(CK),
    .d(\DFF_1136.D ),
    .q(\DFF_1136.Q )
  );
  al_dffl _11596_ (
    .clk(CK),
    .d(\DFF_1137.D ),
    .q(\DFF_1137.Q )
  );
  al_dffl _11597_ (
    .clk(CK),
    .d(\DFF_1138.D ),
    .q(\DFF_1138.Q )
  );
  al_dffl _11598_ (
    .clk(CK),
    .d(\DFF_1139.D ),
    .q(\DFF_1139.Q )
  );
  al_dffl _11599_ (
    .clk(CK),
    .d(\DFF_1140.D ),
    .q(\DFF_1140.Q )
  );
  al_dffl _11600_ (
    .clk(CK),
    .d(\DFF_1141.D ),
    .q(\DFF_1141.Q )
  );
  al_dffl _11601_ (
    .clk(CK),
    .d(\DFF_1142.D ),
    .q(\DFF_1142.Q )
  );
  al_dffl _11602_ (
    .clk(CK),
    .d(\DFF_1143.D ),
    .q(\DFF_1143.Q )
  );
  al_dffl _11603_ (
    .clk(CK),
    .d(\DFF_1144.D ),
    .q(\DFF_1144.Q )
  );
  al_dffl _11604_ (
    .clk(CK),
    .d(\DFF_1145.D ),
    .q(\DFF_1145.Q )
  );
  al_dffl _11605_ (
    .clk(CK),
    .d(\DFF_1146.D ),
    .q(\DFF_1146.Q )
  );
  al_dffl _11606_ (
    .clk(CK),
    .d(\DFF_1147.D ),
    .q(\DFF_1147.Q )
  );
  al_dffl _11607_ (
    .clk(CK),
    .d(\DFF_1148.D ),
    .q(\DFF_1148.Q )
  );
  al_dffl _11608_ (
    .clk(CK),
    .d(\DFF_1149.D ),
    .q(\DFF_1149.Q )
  );
  al_dffl _11609_ (
    .clk(CK),
    .d(\DFF_1150.D ),
    .q(\DFF_1150.Q )
  );
  al_dffl _11610_ (
    .clk(CK),
    .d(\DFF_1151.D ),
    .q(\DFF_1151.Q )
  );
  al_dffl _11611_ (
    .clk(CK),
    .d(\DFF_1152.D ),
    .q(\DFF_1152.Q )
  );
  al_dffl _11612_ (
    .clk(CK),
    .d(\DFF_1153.D ),
    .q(\DFF_1153.Q )
  );
  al_dffl _11613_ (
    .clk(CK),
    .d(\DFF_1154.D ),
    .q(\DFF_1154.Q )
  );
  al_dffl _11614_ (
    .clk(CK),
    .d(\DFF_1156.D ),
    .q(\DFF_1156.Q )
  );
  al_dffl _11615_ (
    .clk(CK),
    .d(\DFF_1157.D ),
    .q(\DFF_1157.Q )
  );
  al_dffl _11616_ (
    .clk(CK),
    .d(\DFF_1159.D ),
    .q(\DFF_1159.Q )
  );
  al_dffl _11617_ (
    .clk(CK),
    .d(\DFF_1160.D ),
    .q(\DFF_1160.Q )
  );
  al_dffl _11618_ (
    .clk(CK),
    .d(\DFF_1161.D ),
    .q(\DFF_1161.Q )
  );
  al_dffl _11619_ (
    .clk(CK),
    .d(\DFF_1162.D ),
    .q(\DFF_1162.Q )
  );
  al_dffl _11620_ (
    .clk(CK),
    .d(\DFF_1163.D ),
    .q(\DFF_1163.Q )
  );
  al_dffl _11621_ (
    .clk(CK),
    .d(\DFF_1164.D ),
    .q(\DFF_1164.Q )
  );
  al_dffl _11622_ (
    .clk(CK),
    .d(\DFF_1165.D ),
    .q(\DFF_1165.Q )
  );
  al_dffl _11623_ (
    .clk(CK),
    .d(\DFF_1166.D ),
    .q(\DFF_1166.Q )
  );
  al_dffl _11624_ (
    .clk(CK),
    .d(\DFF_1167.D ),
    .q(\DFF_1167.Q )
  );
  al_dffl _11625_ (
    .clk(CK),
    .d(\DFF_1168.D ),
    .q(\DFF_1168.Q )
  );
  al_dffl _11626_ (
    .clk(CK),
    .d(\DFF_1169.D ),
    .q(\DFF_1169.Q )
  );
  al_dffl _11627_ (
    .clk(CK),
    .d(\DFF_1170.D ),
    .q(\DFF_1170.Q )
  );
  al_dffl _11628_ (
    .clk(CK),
    .d(\DFF_1171.D ),
    .q(\DFF_1171.Q )
  );
  al_dffl _11629_ (
    .clk(CK),
    .d(\DFF_1172.D ),
    .q(\DFF_1172.Q )
  );
  al_dffl _11630_ (
    .clk(CK),
    .d(\DFF_1173.D ),
    .q(\DFF_1173.Q )
  );
  al_dffl _11631_ (
    .clk(CK),
    .d(\DFF_1174.D ),
    .q(\DFF_1174.Q )
  );
  al_dffl _11632_ (
    .clk(CK),
    .d(\DFF_1175.D ),
    .q(\DFF_1175.Q )
  );
  al_dffl _11633_ (
    .clk(CK),
    .d(\DFF_1100.Q ),
    .q(\DFF_1176.Q )
  );
  al_dffl _11634_ (
    .clk(CK),
    .d(\DFF_1177.D ),
    .q(\DFF_1177.Q )
  );
  al_dffl _11635_ (
    .clk(CK),
    .d(\DFF_1178.D ),
    .q(\DFF_1178.Q )
  );
  al_dffl _11636_ (
    .clk(CK),
    .d(\DFF_1179.D ),
    .q(\DFF_1179.Q )
  );
  al_dffl _11637_ (
    .clk(CK),
    .d(\DFF_1180.D ),
    .q(\DFF_1180.Q )
  );
  al_dffl _11638_ (
    .clk(CK),
    .d(\DFF_1181.D ),
    .q(\DFF_1181.Q )
  );
  al_dffl _11639_ (
    .clk(CK),
    .d(\DFF_1182.D ),
    .q(\DFF_1182.Q )
  );
  al_dffl _11640_ (
    .clk(CK),
    .d(\DFF_1183.D ),
    .q(\DFF_1183.Q )
  );
  al_dffl _11641_ (
    .clk(CK),
    .d(\DFF_1184.D ),
    .q(\DFF_1184.Q )
  );
  al_dffl _11642_ (
    .clk(CK),
    .d(\DFF_1186.D ),
    .q(\DFF_1186.Q )
  );
  al_dffl _11643_ (
    .clk(CK),
    .d(\DFF_1187.D ),
    .q(\DFF_1187.Q )
  );
  al_dffl _11644_ (
    .clk(CK),
    .d(\DFF_1188.D ),
    .q(\DFF_1188.Q )
  );
  al_dffl _11645_ (
    .clk(CK),
    .d(\DFF_1189.D ),
    .q(\DFF_1189.Q )
  );
  al_dffl _11646_ (
    .clk(CK),
    .d(\DFF_1190.D ),
    .q(\DFF_1190.Q )
  );
  al_dffl _11647_ (
    .clk(CK),
    .d(\DFF_1118.Q ),
    .q(\DFF_1191.Q )
  );
  al_dffl _11648_ (
    .clk(CK),
    .d(\DFF_1192.D ),
    .q(\DFF_1192.Q )
  );
  al_dffl _11649_ (
    .clk(CK),
    .d(\DFF_1193.D ),
    .q(\DFF_1193.Q )
  );
  al_dffl _11650_ (
    .clk(CK),
    .d(\DFF_1194.D ),
    .q(\DFF_1194.Q )
  );
  al_dffl _11651_ (
    .clk(CK),
    .d(\DFF_1195.D ),
    .q(\DFF_1195.Q )
  );
  al_dffl _11652_ (
    .clk(CK),
    .d(\DFF_1197.D ),
    .q(\DFF_1197.Q )
  );
  al_dffl _11653_ (
    .clk(CK),
    .d(\DFF_1198.D ),
    .q(\DFF_1198.Q )
  );
  al_dffl _11654_ (
    .clk(CK),
    .d(\DFF_1199.D ),
    .q(\DFF_1199.Q )
  );
  al_dffl _11655_ (
    .clk(CK),
    .d(\DFF_1200.D ),
    .q(\DFF_1200.Q )
  );
  al_dffl _11656_ (
    .clk(CK),
    .d(\DFF_1201.D ),
    .q(\DFF_1201.Q )
  );
  al_dffl _11657_ (
    .clk(CK),
    .d(\DFF_1202.D ),
    .q(\DFF_1202.Q )
  );
  al_dffl _11658_ (
    .clk(CK),
    .d(\DFF_1203.D ),
    .q(\DFF_1203.Q )
  );
  al_dffl _11659_ (
    .clk(CK),
    .d(\DFF_1204.D ),
    .q(\DFF_1204.Q )
  );
  al_dffl _11660_ (
    .clk(CK),
    .d(\DFF_1205.D ),
    .q(\DFF_1205.Q )
  );
  al_dffl _11661_ (
    .clk(CK),
    .d(\DFF_1206.D ),
    .q(\DFF_1206.Q )
  );
  al_dffl _11662_ (
    .clk(CK),
    .d(\DFF_1208.D ),
    .q(\DFF_1208.Q )
  );
  al_dffl _11663_ (
    .clk(CK),
    .d(\DFF_991.Q ),
    .q(\DFF_1209.Q )
  );
  al_dffl _11664_ (
    .clk(CK),
    .d(\DFF_1210.D ),
    .q(\DFF_1210.Q )
  );
  al_dffl _11665_ (
    .clk(CK),
    .d(\DFF_1211.D ),
    .q(\DFF_1211.Q )
  );
  al_dffl _11666_ (
    .clk(CK),
    .d(\DFF_1212.D ),
    .q(\DFF_1212.Q )
  );
  al_dffl _11667_ (
    .clk(CK),
    .d(\DFF_1213.D ),
    .q(\DFF_1213.Q )
  );
  al_dffl _11668_ (
    .clk(CK),
    .d(\DFF_1214.D ),
    .q(\DFF_1214.Q )
  );
  al_dffl _11669_ (
    .clk(CK),
    .d(\DFF_1215.D ),
    .q(\DFF_1215.Q )
  );
  al_dffl _11670_ (
    .clk(CK),
    .d(\DFF_1216.D ),
    .q(\DFF_1216.Q )
  );
  al_dffl _11671_ (
    .clk(CK),
    .d(\DFF_1217.D ),
    .q(\DFF_1217.Q )
  );
  al_dffl _11672_ (
    .clk(CK),
    .d(\DFF_1218.D ),
    .q(\DFF_1218.Q )
  );
  al_dffl _11673_ (
    .clk(CK),
    .d(\DFF_1220.D ),
    .q(\DFF_1220.Q )
  );
  al_dffl _11674_ (
    .clk(CK),
    .d(\DFF_1221.D ),
    .q(\DFF_1221.Q )
  );
  al_dffl _11675_ (
    .clk(CK),
    .d(\DFF_1222.D ),
    .q(\DFF_1222.Q )
  );
  al_dffl _11676_ (
    .clk(CK),
    .d(\DFF_1223.D ),
    .q(\DFF_1223.Q )
  );
  al_dffl _11677_ (
    .clk(CK),
    .d(\DFF_1226.D ),
    .q(\DFF_1226.Q )
  );
  al_dffl _11678_ (
    .clk(CK),
    .d(\DFF_1227.D ),
    .q(\DFF_1227.Q )
  );
  al_dffl _11679_ (
    .clk(CK),
    .d(\DFF_545.Q ),
    .q(\DFF_1228.Q )
  );
  al_dffl _11680_ (
    .clk(CK),
    .d(\DFF_1229.D ),
    .q(\DFF_1229.Q )
  );
  al_dffl _11681_ (
    .clk(CK),
    .d(\DFF_1230.D ),
    .q(\DFF_1230.Q )
  );
  al_dffl _11682_ (
    .clk(CK),
    .d(\DFF_1231.D ),
    .q(\DFF_1231.Q )
  );
  al_dffl _11683_ (
    .clk(CK),
    .d(\DFF_1232.D ),
    .q(\DFF_1232.Q )
  );
  al_dffl _11684_ (
    .clk(CK),
    .d(\DFF_1233.D ),
    .q(\DFF_1233.Q )
  );
  al_dffl _11685_ (
    .clk(CK),
    .d(\DFF_1235.D ),
    .q(\DFF_1235.Q )
  );
  al_dffl _11686_ (
    .clk(CK),
    .d(\DFF_1236.D ),
    .q(\DFF_1236.Q )
  );
  al_dffl _11687_ (
    .clk(CK),
    .d(\DFF_1237.D ),
    .q(\DFF_1237.Q )
  );
  al_dffl _11688_ (
    .clk(CK),
    .d(\DFF_1238.D ),
    .q(\DFF_1238.Q )
  );
  al_dffl _11689_ (
    .clk(CK),
    .d(\DFF_1239.D ),
    .q(\DFF_1239.Q )
  );
  al_dffl _11690_ (
    .clk(CK),
    .d(\DFF_1240.D ),
    .q(\DFF_1240.Q )
  );
  al_dffl _11691_ (
    .clk(CK),
    .d(\DFF_1241.D ),
    .q(\DFF_1241.Q )
  );
  al_dffl _11692_ (
    .clk(CK),
    .d(\DFF_1242.D ),
    .q(\DFF_1242.Q )
  );
  al_dffl _11693_ (
    .clk(CK),
    .d(\DFF_1243.D ),
    .q(\DFF_1243.Q )
  );
  al_dffl _11694_ (
    .clk(CK),
    .d(\DFF_1244.D ),
    .q(\DFF_1244.Q )
  );
  al_dffl _11695_ (
    .clk(CK),
    .d(\DFF_1245.D ),
    .q(\DFF_1245.Q )
  );
  al_dffl _11696_ (
    .clk(CK),
    .d(\DFF_1246.D ),
    .q(\DFF_1246.Q )
  );
  al_dffl _11697_ (
    .clk(CK),
    .d(\DFF_1247.D ),
    .q(\DFF_1247.Q )
  );
  al_dffl _11698_ (
    .clk(CK),
    .d(\DFF_1249.D ),
    .q(\DFF_1249.Q )
  );
  al_dffl _11699_ (
    .clk(CK),
    .d(\DFF_1250.D ),
    .q(\DFF_1250.Q )
  );
  al_dffl _11700_ (
    .clk(CK),
    .d(\DFF_1251.D ),
    .q(\DFF_1251.Q )
  );
  al_dffl _11701_ (
    .clk(CK),
    .d(\DFF_1252.D ),
    .q(\DFF_1252.Q )
  );
  al_dffl _11702_ (
    .clk(CK),
    .d(\DFF_1253.D ),
    .q(\DFF_1253.Q )
  );
  al_dffl _11703_ (
    .clk(CK),
    .d(\DFF_1254.D ),
    .q(\DFF_1254.Q )
  );
  al_dffl _11704_ (
    .clk(CK),
    .d(\DFF_1255.D ),
    .q(\DFF_1255.Q )
  );
  al_dffl _11705_ (
    .clk(CK),
    .d(\DFF_1257.D ),
    .q(\DFF_1257.Q )
  );
  al_dffl _11706_ (
    .clk(CK),
    .d(\DFF_1258.D ),
    .q(\DFF_1258.Q )
  );
  al_dffl _11707_ (
    .clk(CK),
    .d(\DFF_1259.D ),
    .q(\DFF_1259.Q )
  );
  al_dffl _11708_ (
    .clk(CK),
    .d(\DFF_1260.D ),
    .q(\DFF_1260.Q )
  );
  al_dffl _11709_ (
    .clk(CK),
    .d(\DFF_1261.D ),
    .q(\DFF_1261.Q )
  );
  al_dffl _11710_ (
    .clk(CK),
    .d(\DFF_1263.D ),
    .q(\DFF_1263.Q )
  );
  al_dffl _11711_ (
    .clk(CK),
    .d(\DFF_1264.D ),
    .q(\DFF_1264.Q )
  );
  al_dffl _11712_ (
    .clk(CK),
    .d(\DFF_1266.D ),
    .q(\DFF_1266.Q )
  );
  al_dffl _11713_ (
    .clk(CK),
    .d(\DFF_1267.D ),
    .q(\DFF_1267.Q )
  );
  al_dffl _11714_ (
    .clk(CK),
    .d(\DFF_1268.D ),
    .q(\DFF_1268.Q )
  );
  al_dffl _11715_ (
    .clk(CK),
    .d(\DFF_1269.D ),
    .q(\DFF_1269.Q )
  );
  al_dffl _11716_ (
    .clk(CK),
    .d(\DFF_1270.D ),
    .q(\DFF_1270.Q )
  );
  al_dffl _11717_ (
    .clk(CK),
    .d(\DFF_1271.D ),
    .q(\DFF_1271.Q )
  );
  al_dffl _11718_ (
    .clk(CK),
    .d(\DFF_1272.D ),
    .q(\DFF_1272.Q )
  );
  al_dffl _11719_ (
    .clk(CK),
    .d(\DFF_1273.D ),
    .q(\DFF_1273.Q )
  );
  al_dffl _11720_ (
    .clk(CK),
    .d(\DFF_1274.D ),
    .q(\DFF_1274.Q )
  );
  al_dffl _11721_ (
    .clk(CK),
    .d(\DFF_1276.D ),
    .q(\DFF_1276.Q )
  );
  al_dffl _11722_ (
    .clk(CK),
    .d(\DFF_1277.D ),
    .q(\DFF_1277.Q )
  );
  al_dffl _11723_ (
    .clk(CK),
    .d(\DFF_1278.D ),
    .q(\DFF_1278.Q )
  );
  al_dffl _11724_ (
    .clk(CK),
    .d(\DFF_1279.D ),
    .q(\DFF_1279.Q )
  );
  al_dffl _11725_ (
    .clk(CK),
    .d(\DFF_1280.D ),
    .q(\DFF_1280.Q )
  );
  al_dffl _11726_ (
    .clk(CK),
    .d(\DFF_1281.D ),
    .q(\DFF_1281.Q )
  );
  al_dffl _11727_ (
    .clk(CK),
    .d(\DFF_1282.D ),
    .q(\DFF_1282.Q )
  );
  al_dffl _11728_ (
    .clk(CK),
    .d(\DFF_1283.D ),
    .q(\DFF_1283.Q )
  );
  al_dffl _11729_ (
    .clk(CK),
    .d(\DFF_1284.D ),
    .q(\DFF_1284.Q )
  );
  al_dffl _11730_ (
    .clk(CK),
    .d(\DFF_1285.D ),
    .q(\DFF_1285.Q )
  );
  al_dffl _11731_ (
    .clk(CK),
    .d(\DFF_1287.D ),
    .q(\DFF_1287.Q )
  );
  al_dffl _11732_ (
    .clk(CK),
    .d(\DFF_1288.D ),
    .q(\DFF_1288.Q )
  );
  al_dffl _11733_ (
    .clk(CK),
    .d(\DFF_1289.D ),
    .q(\DFF_1289.Q )
  );
  al_dffl _11734_ (
    .clk(CK),
    .d(\DFF_1290.D ),
    .q(\DFF_1290.Q )
  );
  al_dffl _11735_ (
    .clk(CK),
    .d(\DFF_1291.D ),
    .q(\DFF_1291.Q )
  );
  al_dffl _11736_ (
    .clk(CK),
    .d(\DFF_1292.D ),
    .q(\DFF_1292.Q )
  );
  al_dffl _11737_ (
    .clk(CK),
    .d(\DFF_1294.D ),
    .q(\DFF_1294.Q )
  );
  al_dffl _11738_ (
    .clk(CK),
    .d(\DFF_1295.D ),
    .q(\DFF_1295.Q )
  );
  al_dffl _11739_ (
    .clk(CK),
    .d(\DFF_1296.D ),
    .q(\DFF_1296.Q )
  );
  al_dffl _11740_ (
    .clk(CK),
    .d(\DFF_1297.D ),
    .q(\DFF_1297.Q )
  );
  al_dffl _11741_ (
    .clk(CK),
    .d(\DFF_1298.D ),
    .q(\DFF_1298.Q )
  );
  al_dffl _11742_ (
    .clk(CK),
    .d(\DFF_1299.D ),
    .q(\DFF_1299.Q )
  );
  al_dffl _11743_ (
    .clk(CK),
    .d(\DFF_1301.D ),
    .q(\DFF_1301.Q )
  );
  al_dffl _11744_ (
    .clk(CK),
    .d(\DFF_1302.D ),
    .q(\DFF_1302.Q )
  );
  al_dffl _11745_ (
    .clk(CK),
    .d(\DFF_76.Q ),
    .q(\DFF_1359.Q )
  );
  al_dffl _11746_ (
    .clk(CK),
    .d(\DFF_1359.Q ),
    .q(\DFF_1303.Q )
  );
  al_dffl _11747_ (
    .clk(CK),
    .d(\DFF_1304.D ),
    .q(\DFF_1304.Q )
  );
  al_dffl _11748_ (
    .clk(CK),
    .d(\DFF_1305.D ),
    .q(\DFF_1305.Q )
  );
  al_dffl _11749_ (
    .clk(CK),
    .d(\DFF_1306.D ),
    .q(\DFF_1306.Q )
  );
  al_dffl _11750_ (
    .clk(CK),
    .d(\DFF_1307.D ),
    .q(\DFF_1307.Q )
  );
  al_dffl _11751_ (
    .clk(CK),
    .d(\DFF_1309.D ),
    .q(\DFF_1309.Q )
  );
  al_dffl _11752_ (
    .clk(CK),
    .d(\DFF_1310.D ),
    .q(\DFF_1310.Q )
  );
  al_dffl _11753_ (
    .clk(CK),
    .d(\DFF_1311.D ),
    .q(\DFF_1311.Q )
  );
  al_dffl _11754_ (
    .clk(CK),
    .d(\DFF_1312.D ),
    .q(\DFF_1312.Q )
  );
  al_dffl _11755_ (
    .clk(CK),
    .d(\DFF_1313.D ),
    .q(\DFF_1313.Q )
  );
  al_dffl _11756_ (
    .clk(CK),
    .d(\DFF_1314.D ),
    .q(\DFF_1314.Q )
  );
  al_dffl _11757_ (
    .clk(CK),
    .d(\DFF_1315.D ),
    .q(\DFF_1315.Q )
  );
  al_dffl _11758_ (
    .clk(CK),
    .d(\DFF_1317.D ),
    .q(\DFF_1317.Q )
  );
  al_dffl _11759_ (
    .clk(CK),
    .d(\DFF_1318.D ),
    .q(\DFF_1318.Q )
  );
  al_dffl _11760_ (
    .clk(CK),
    .d(\DFF_1319.D ),
    .q(\DFF_1319.Q )
  );
  al_dffl _11761_ (
    .clk(CK),
    .d(\DFF_1320.D ),
    .q(\DFF_1320.Q )
  );
  al_dffl _11762_ (
    .clk(CK),
    .d(\DFF_1321.D ),
    .q(\DFF_1321.Q )
  );
  al_dffl _11763_ (
    .clk(CK),
    .d(\DFF_1322.D ),
    .q(\DFF_1322.Q )
  );
  al_dffl _11764_ (
    .clk(CK),
    .d(\DFF_1323.D ),
    .q(\DFF_1323.Q )
  );
  al_dffl _11765_ (
    .clk(CK),
    .d(\DFF_1324.D ),
    .q(\DFF_1324.Q )
  );
  al_dffl _11766_ (
    .clk(CK),
    .d(\DFF_1325.D ),
    .q(\DFF_1325.Q )
  );
  al_dffl _11767_ (
    .clk(CK),
    .d(\DFF_1326.D ),
    .q(\DFF_1326.Q )
  );
  al_dffl _11768_ (
    .clk(CK),
    .d(\DFF_1327.D ),
    .q(\DFF_1327.Q )
  );
  al_dffl _11769_ (
    .clk(CK),
    .d(\DFF_1328.D ),
    .q(\DFF_1328.Q )
  );
  al_dffl _11770_ (
    .clk(CK),
    .d(\DFF_1329.D ),
    .q(\DFF_1329.Q )
  );
  al_dffl _11771_ (
    .clk(CK),
    .d(\DFF_1330.D ),
    .q(\DFF_1330.Q )
  );
  al_dffl _11772_ (
    .clk(CK),
    .d(\DFF_1331.D ),
    .q(\DFF_1331.Q )
  );
  al_dffl _11773_ (
    .clk(CK),
    .d(\DFF_1332.D ),
    .q(\DFF_1332.Q )
  );
  al_dffl _11774_ (
    .clk(CK),
    .d(\DFF_1333.D ),
    .q(\DFF_1333.Q )
  );
  al_dffl _11775_ (
    .clk(CK),
    .d(\DFF_1334.D ),
    .q(\DFF_1334.Q )
  );
  al_dffl _11776_ (
    .clk(CK),
    .d(\DFF_1336.D ),
    .q(\DFF_1336.Q )
  );
  al_dffl _11777_ (
    .clk(CK),
    .d(\DFF_1337.D ),
    .q(\DFF_1337.Q )
  );
  al_dffl _11778_ (
    .clk(CK),
    .d(\DFF_1339.D ),
    .q(\DFF_1339.Q )
  );
  al_dffl _11779_ (
    .clk(CK),
    .d(\DFF_1340.D ),
    .q(\DFF_1340.Q )
  );
  al_dffl _11780_ (
    .clk(CK),
    .d(\DFF_1341.D ),
    .q(\DFF_1341.Q )
  );
  al_dffl _11781_ (
    .clk(CK),
    .d(\DFF_1342.D ),
    .q(\DFF_1342.Q )
  );
  al_dffl _11782_ (
    .clk(CK),
    .d(\DFF_1343.D ),
    .q(\DFF_1343.Q )
  );
  al_dffl _11783_ (
    .clk(CK),
    .d(\DFF_1344.D ),
    .q(\DFF_1344.Q )
  );
  al_dffl _11784_ (
    .clk(CK),
    .d(\DFF_1345.D ),
    .q(\DFF_1345.Q )
  );
  al_dffl _11785_ (
    .clk(CK),
    .d(\DFF_1346.D ),
    .q(\DFF_1346.Q )
  );
  al_dffl _11786_ (
    .clk(CK),
    .d(\DFF_1347.D ),
    .q(\DFF_1347.Q )
  );
  al_dffl _11787_ (
    .clk(CK),
    .d(\DFF_1348.D ),
    .q(\DFF_1348.Q )
  );
  al_dffl _11788_ (
    .clk(CK),
    .d(\DFF_1349.D ),
    .q(\DFF_1349.Q )
  );
  al_dffl _11789_ (
    .clk(CK),
    .d(\DFF_1350.D ),
    .q(\DFF_1350.Q )
  );
  al_dffl _11790_ (
    .clk(CK),
    .d(\DFF_1351.D ),
    .q(\DFF_1351.Q )
  );
  al_dffl _11791_ (
    .clk(CK),
    .d(\DFF_1353.D ),
    .q(\DFF_1353.Q )
  );
  al_dffl _11792_ (
    .clk(CK),
    .d(\DFF_1355.D ),
    .q(\DFF_1355.Q )
  );
  al_dffl _11793_ (
    .clk(CK),
    .d(\DFF_1356.D ),
    .q(\DFF_1356.Q )
  );
  al_dffl _11794_ (
    .clk(CK),
    .d(\DFF_1357.D ),
    .q(\DFF_1357.Q )
  );
  al_dffl _11795_ (
    .clk(CK),
    .d(\DFF_1358.D ),
    .q(\DFF_1358.Q )
  );
  al_dffl _11796_ (
    .clk(CK),
    .d(\DFF_1360.D ),
    .q(\DFF_1360.Q )
  );
  al_dffl _11797_ (
    .clk(CK),
    .d(\DFF_1361.D ),
    .q(\DFF_1361.Q )
  );
  al_dffl _11798_ (
    .clk(CK),
    .d(\DFF_1362.D ),
    .q(\DFF_1362.Q )
  );
  al_dffl _11799_ (
    .clk(CK),
    .d(\DFF_1363.D ),
    .q(\DFF_1363.Q )
  );
  al_dffl _11800_ (
    .clk(CK),
    .d(\DFF_1364.D ),
    .q(\DFF_1364.Q )
  );
  al_dffl _11801_ (
    .clk(CK),
    .d(\DFF_1365.D ),
    .q(\DFF_1365.Q )
  );
  al_dffl _11802_ (
    .clk(CK),
    .d(\DFF_1366.D ),
    .q(\DFF_1366.Q )
  );
  al_dffl _11803_ (
    .clk(CK),
    .d(\DFF_1367.D ),
    .q(\DFF_1367.Q )
  );
  al_dffl _11804_ (
    .clk(CK),
    .d(\DFF_1368.D ),
    .q(\DFF_1368.Q )
  );
  al_dffl _11805_ (
    .clk(CK),
    .d(\DFF_1369.D ),
    .q(\DFF_1369.Q )
  );
  al_dffl _11806_ (
    .clk(CK),
    .d(\DFF_1370.D ),
    .q(\DFF_1370.Q )
  );
  al_dffl _11807_ (
    .clk(CK),
    .d(\DFF_1371.D ),
    .q(\DFF_1371.Q )
  );
  al_dffl _11808_ (
    .clk(CK),
    .d(\DFF_1372.D ),
    .q(\DFF_1372.Q )
  );
  al_dffl _11809_ (
    .clk(CK),
    .d(\DFF_1373.D ),
    .q(\DFF_1373.Q )
  );
  al_dffl _11810_ (
    .clk(CK),
    .d(\DFF_1374.D ),
    .q(\DFF_1374.Q )
  );
  al_dffl _11811_ (
    .clk(CK),
    .d(\DFF_1375.D ),
    .q(\DFF_1375.Q )
  );
  al_dffl _11812_ (
    .clk(CK),
    .d(\DFF_1376.D ),
    .q(\DFF_1376.Q )
  );
  al_dffl _11813_ (
    .clk(CK),
    .d(\DFF_1377.D ),
    .q(\DFF_1377.Q )
  );
  al_dffl _11814_ (
    .clk(CK),
    .d(\DFF_1378.D ),
    .q(\DFF_1378.Q )
  );
  al_dffl _11815_ (
    .clk(CK),
    .d(\DFF_1379.D ),
    .q(\DFF_1379.Q )
  );
  al_dffl _11816_ (
    .clk(CK),
    .d(\DFF_1380.D ),
    .q(\DFF_1380.Q )
  );
  al_dffl _11817_ (
    .clk(CK),
    .d(\DFF_1381.D ),
    .q(\DFF_1381.Q )
  );
  al_dffl _11818_ (
    .clk(CK),
    .d(\DFF_1382.D ),
    .q(\DFF_1382.Q )
  );
  al_dffl _11819_ (
    .clk(CK),
    .d(\DFF_1383.D ),
    .q(\DFF_1383.Q )
  );
  al_dffl _11820_ (
    .clk(CK),
    .d(\DFF_1384.D ),
    .q(\DFF_1384.Q )
  );
  al_dffl _11821_ (
    .clk(CK),
    .d(\DFF_1385.D ),
    .q(\DFF_1385.Q )
  );
  al_dffl _11822_ (
    .clk(CK),
    .d(\DFF_1386.D ),
    .q(\DFF_1386.Q )
  );
  al_dffl _11823_ (
    .clk(CK),
    .d(\DFF_1387.D ),
    .q(\DFF_1387.Q )
  );
  al_dffl _11824_ (
    .clk(CK),
    .d(\DFF_1388.D ),
    .q(\DFF_1388.Q )
  );
  al_dffl _11825_ (
    .clk(CK),
    .d(\DFF_704.Q ),
    .q(\DFF_1389.Q )
  );
  al_dffl _11826_ (
    .clk(CK),
    .d(\DFF_1390.D ),
    .q(\DFF_1390.Q )
  );
  al_dffl _11827_ (
    .clk(CK),
    .d(\DFF_1391.D ),
    .q(\DFF_1391.Q )
  );
  al_dffl _11828_ (
    .clk(CK),
    .d(\DFF_1392.D ),
    .q(\DFF_1392.Q )
  );
  al_dffl _11829_ (
    .clk(CK),
    .d(\DFF_1393.D ),
    .q(\DFF_1393.Q )
  );
  al_dffl _11830_ (
    .clk(CK),
    .d(\DFF_1394.D ),
    .q(\DFF_1394.Q )
  );
  al_dffl _11831_ (
    .clk(CK),
    .d(\DFF_1395.D ),
    .q(\DFF_1395.Q )
  );
  al_dffl _11832_ (
    .clk(CK),
    .d(\DFF_630.Q ),
    .q(\DFF_1396.Q )
  );
  al_dffl _11833_ (
    .clk(CK),
    .d(\DFF_1397.D ),
    .q(\DFF_1397.Q )
  );
  al_dffl _11834_ (
    .clk(CK),
    .d(\DFF_1398.D ),
    .q(\DFF_1398.Q )
  );
  al_dffl _11835_ (
    .clk(CK),
    .d(\DFF_1399.D ),
    .q(\DFF_1399.Q )
  );
  al_dffl _11836_ (
    .clk(CK),
    .d(\DFF_1400.D ),
    .q(\DFF_1400.Q )
  );
  al_dffl _11837_ (
    .clk(CK),
    .d(\DFF_1401.D ),
    .q(\DFF_1401.Q )
  );
  al_dffl _11838_ (
    .clk(CK),
    .d(\DFF_1402.D ),
    .q(\DFF_1402.Q )
  );
  al_dffl _11839_ (
    .clk(CK),
    .d(\DFF_1403.D ),
    .q(\DFF_1403.Q )
  );
  al_dffl _11840_ (
    .clk(CK),
    .d(\DFF_1404.D ),
    .q(\DFF_1404.Q )
  );
  al_dffl _11841_ (
    .clk(CK),
    .d(\DFF_1405.D ),
    .q(\DFF_1405.Q )
  );
  al_dffl _11842_ (
    .clk(CK),
    .d(\DFF_1406.D ),
    .q(\DFF_1406.Q )
  );
  al_dffl _11843_ (
    .clk(CK),
    .d(\DFF_1407.D ),
    .q(\DFF_1407.Q )
  );
  al_dffl _11844_ (
    .clk(CK),
    .d(\DFF_1408.D ),
    .q(\DFF_1408.Q )
  );
  al_dffl _11845_ (
    .clk(CK),
    .d(\DFF_1409.D ),
    .q(\DFF_1409.Q )
  );
  al_dffl _11846_ (
    .clk(CK),
    .d(\DFF_1410.D ),
    .q(\DFF_1410.Q )
  );
  al_dffl _11847_ (
    .clk(CK),
    .d(\DFF_1411.D ),
    .q(\DFF_1411.Q )
  );
  al_dffl _11848_ (
    .clk(CK),
    .d(\DFF_1412.D ),
    .q(\DFF_1412.Q )
  );
  al_dffl _11849_ (
    .clk(CK),
    .d(\DFF_1413.D ),
    .q(\DFF_1413.Q )
  );
  al_dffl _11850_ (
    .clk(CK),
    .d(\DFF_1415.D ),
    .q(\DFF_1415.Q )
  );
  al_dffl _11851_ (
    .clk(CK),
    .d(\DFF_1417.D ),
    .q(\DFF_1417.Q )
  );
  al_dffl _11852_ (
    .clk(CK),
    .d(\DFF_1418.D ),
    .q(\DFF_1418.Q )
  );
  al_dffl _11853_ (
    .clk(CK),
    .d(\DFF_1419.D ),
    .q(\DFF_1419.Q )
  );
  al_dffl _11854_ (
    .clk(CK),
    .d(\DFF_1422.D ),
    .q(\DFF_1422.Q )
  );
  al_dffl _11855_ (
    .clk(CK),
    .d(\DFF_1423.D ),
    .q(\DFF_1423.Q )
  );
  al_dffl _11856_ (
    .clk(CK),
    .d(\DFF_1424.D ),
    .q(\DFF_1424.Q )
  );
  al_dffl _11857_ (
    .clk(CK),
    .d(\DFF_1425.D ),
    .q(\DFF_1425.Q )
  );
  assign \DFF_0.CK  = CK;
  assign \DFF_1.CK  = CK;
  assign \DFF_10.CK  = CK;
  assign \DFF_100.CK  = CK;
  assign \DFF_1000.CK  = CK;
  assign \DFF_1001.CK  = CK;
  assign \DFF_1002.CK  = CK;
  assign \DFF_1002.D  = \DFF_1073.Q ;
  assign \DFF_1003.CK  = CK;
  assign \DFF_1003.D  = \DFF_764.Q ;
  assign \DFF_1004.CK  = CK;
  assign \DFF_1005.CK  = CK;
  assign \DFF_1006.CK  = CK;
  assign \DFF_1007.CK  = CK;
  assign \DFF_1008.CK  = CK;
  assign \DFF_1009.CK  = CK;
  assign \DFF_101.CK  = CK;
  assign \DFF_101.D  = \DFF_263.Q ;
  assign \DFF_1010.CK  = CK;
  assign \DFF_1011.CK  = CK;
  assign \DFF_1012.CK  = CK;
  assign \DFF_1013.CK  = CK;
  assign \DFF_1014.CK  = CK;
  assign \DFF_1014.D  = \DFF_686.Q ;
  assign \DFF_1015.CK  = CK;
  assign \DFF_1016.CK  = CK;
  assign \DFF_1017.CK  = CK;
  assign \DFF_1018.CK  = CK;
  assign \DFF_1019.CK  = CK;
  assign \DFF_102.CK  = CK;
  assign \DFF_1020.CK  = CK;
  assign \DFF_1021.CK  = CK;
  assign \DFF_1022.CK  = CK;
  assign \DFF_1023.CK  = CK;
  assign \DFF_1023.D  = \DFF_780.Q ;
  assign \DFF_1024.CK  = CK;
  assign \DFF_1025.CK  = CK;
  assign \DFF_1026.CK  = CK;
  assign \DFF_1027.CK  = CK;
  assign \DFF_1028.CK  = CK;
  assign \DFF_1029.CK  = CK;
  assign \DFF_103.CK  = CK;
  assign \DFF_1030.CK  = CK;
  assign \DFF_1031.CK  = CK;
  assign \DFF_1032.CK  = CK;
  assign \DFF_1033.CK  = CK;
  assign \DFF_1034.CK  = CK;
  assign \DFF_1035.CK  = CK;
  assign \DFF_1036.CK  = CK;
  assign \DFF_1037.CK  = CK;
  assign \DFF_1038.CK  = CK;
  assign \DFF_1038.D  = \DFF_529.Q ;
  assign \DFF_1039.CK  = CK;
  assign \DFF_104.CK  = CK;
  assign \DFF_1040.CK  = CK;
  assign \DFF_1041.CK  = CK;
  assign \DFF_1042.CK  = CK;
  assign \DFF_1043.CK  = CK;
  assign \DFF_1043.D  = \DFF_1027.Q ;
  assign \DFF_1044.CK  = CK;
  assign \DFF_1045.CK  = CK;
  assign \DFF_1046.CK  = CK;
  assign \DFF_1047.CK  = CK;
  assign \DFF_1048.CK  = CK;
  assign \DFF_1049.CK  = CK;
  assign \DFF_1049.D  = \DFF_1416.Q ;
  assign \DFF_105.CK  = CK;
  assign \DFF_1050.CK  = CK;
  assign \DFF_1051.CK  = CK;
  assign \DFF_1052.CK  = CK;
  assign \DFF_1053.CK  = CK;
  assign \DFF_1054.CK  = CK;
  assign \DFF_1055.CK  = CK;
  assign \DFF_1056.CK  = CK;
  assign \DFF_1057.CK  = CK;
  assign \DFF_1058.CK  = CK;
  assign \DFF_1059.CK  = CK;
  assign \DFF_106.CK  = CK;
  assign \DFF_1060.CK  = CK;
  assign \DFF_1061.CK  = CK;
  assign \DFF_1061.D  = \DFF_612.Q ;
  assign \DFF_1062.CK  = CK;
  assign \DFF_1063.CK  = CK;
  assign \DFF_1064.CK  = CK;
  assign \DFF_1065.CK  = CK;
  assign \DFF_1066.CK  = CK;
  assign \DFF_1067.CK  = CK;
  assign \DFF_1068.CK  = CK;
  assign \DFF_1069.CK  = CK;
  assign \DFF_107.CK  = CK;
  assign \DFF_1070.CK  = CK;
  assign \DFF_1071.CK  = CK;
  assign \DFF_1072.CK  = CK;
  assign \DFF_1073.CK  = CK;
  assign \DFF_1074.CK  = CK;
  assign \DFF_1075.CK  = CK;
  assign \DFF_1076.CK  = CK;
  assign \DFF_1077.CK  = CK;
  assign \DFF_1078.CK  = CK;
  assign \DFF_1079.CK  = CK;
  assign \DFF_108.CK  = CK;
  assign \DFF_1080.CK  = CK;
  assign \DFF_1081.CK  = CK;
  assign \DFF_1081.D  = \DFF_515.Q ;
  assign \DFF_1082.CK  = CK;
  assign \DFF_1083.CK  = CK;
  assign \DFF_1084.CK  = CK;
  assign \DFF_1085.CK  = CK;
  assign \DFF_1086.CK  = CK;
  assign \DFF_1087.CK  = CK;
  assign \DFF_1087.D  = \DFF_737.Q ;
  assign \DFF_1088.CK  = CK;
  assign \DFF_1089.CK  = CK;
  assign \DFF_109.CK  = CK;
  assign \DFF_109.D  = \DFF_752.Q ;
  assign \DFF_1090.CK  = CK;
  assign \DFF_1091.CK  = CK;
  assign \DFF_1092.CK  = CK;
  assign \DFF_1093.CK  = CK;
  assign \DFF_1094.CK  = CK;
  assign \DFF_1095.CK  = CK;
  assign \DFF_1096.CK  = CK;
  assign \DFF_1097.CK  = CK;
  assign \DFF_1098.CK  = CK;
  assign \DFF_1099.CK  = CK;
  assign \DFF_11.CK  = CK;
  assign \DFF_110.CK  = CK;
  assign \DFF_110.D  = \DFF_797.Q ;
  assign \DFF_1100.CK  = CK;
  assign \DFF_1100.D  = \DFF_981.Q ;
  assign \DFF_1101.CK  = CK;
  assign \DFF_1102.CK  = CK;
  assign \DFF_1102.D  = \DFF_848.Q ;
  assign \DFF_1103.CK  = CK;
  assign \DFF_1104.CK  = CK;
  assign \DFF_1105.CK  = CK;
  assign \DFF_1106.CK  = CK;
  assign \DFF_1106.D  = \DFF_561.Q ;
  assign \DFF_1107.CK  = CK;
  assign \DFF_1108.CK  = CK;
  assign \DFF_1109.CK  = CK;
  assign \DFF_111.CK  = CK;
  assign \DFF_1110.CK  = CK;
  assign \DFF_1110.D  = \DFF_146.Q ;
  assign \DFF_1111.CK  = CK;
  assign \DFF_1112.CK  = CK;
  assign \DFF_1113.CK  = CK;
  assign \DFF_1114.CK  = CK;
  assign \DFF_1115.CK  = CK;
  assign \DFF_1116.CK  = CK;
  assign \DFF_1117.CK  = CK;
  assign \DFF_1118.CK  = CK;
  assign \DFF_1118.D  = \DFF_997.Q ;
  assign \DFF_1119.CK  = CK;
  assign \DFF_1119.D  = \DFF_123.Q ;
  assign \DFF_112.CK  = CK;
  assign \DFF_1120.CK  = CK;
  assign \DFF_1121.CK  = CK;
  assign \DFF_1122.CK  = CK;
  assign \DFF_1122.D  = \DFF_643.Q ;
  assign \DFF_1123.CK  = CK;
  assign \DFF_1124.CK  = CK;
  assign \DFF_1125.CK  = CK;
  assign \DFF_1126.CK  = CK;
  assign \DFF_1127.CK  = CK;
  assign \DFF_1128.CK  = CK;
  assign \DFF_1129.CK  = CK;
  assign \DFF_113.CK  = CK;
  assign \DFF_1130.CK  = CK;
  assign \DFF_1131.CK  = CK;
  assign \DFF_1132.CK  = CK;
  assign \DFF_1133.CK  = CK;
  assign \DFF_1134.CK  = CK;
  assign \DFF_1135.CK  = CK;
  assign \DFF_1136.CK  = CK;
  assign \DFF_1137.CK  = CK;
  assign \DFF_1138.CK  = CK;
  assign \DFF_1139.CK  = CK;
  assign \DFF_114.CK  = CK;
  assign \DFF_1140.CK  = CK;
  assign \DFF_1141.CK  = CK;
  assign \DFF_1142.CK  = CK;
  assign \DFF_1143.CK  = CK;
  assign \DFF_1144.CK  = CK;
  assign \DFF_1145.CK  = CK;
  assign \DFF_1146.CK  = CK;
  assign \DFF_1147.CK  = CK;
  assign \DFF_1148.CK  = CK;
  assign \DFF_1149.CK  = CK;
  assign \DFF_115.CK  = CK;
  assign \DFF_1150.CK  = CK;
  assign \DFF_1151.CK  = CK;
  assign \DFF_1152.CK  = CK;
  assign \DFF_1153.CK  = CK;
  assign \DFF_1154.CK  = CK;
  assign \DFF_1155.CK  = CK;
  assign \DFF_1155.D  = \DFF_1354.Q ;
  assign \DFF_1156.CK  = CK;
  assign \DFF_1157.CK  = CK;
  assign \DFF_1158.CK  = CK;
  assign \DFF_1159.CK  = CK;
  assign \DFF_116.CK  = CK;
  assign \DFF_1160.CK  = CK;
  assign \DFF_1161.CK  = CK;
  assign \DFF_1162.CK  = CK;
  assign \DFF_1163.CK  = CK;
  assign \DFF_1164.CK  = CK;
  assign \DFF_1165.CK  = CK;
  assign \DFF_1166.CK  = CK;
  assign \DFF_1167.CK  = CK;
  assign \DFF_1168.CK  = CK;
  assign \DFF_1169.CK  = CK;
  assign \DFF_117.CK  = CK;
  assign \DFF_117.D  = \DFF_1335.Q ;
  assign \DFF_1170.CK  = CK;
  assign \DFF_1171.CK  = CK;
  assign \DFF_1172.CK  = CK;
  assign \DFF_1173.CK  = CK;
  assign \DFF_1174.CK  = CK;
  assign \DFF_1175.CK  = CK;
  assign \DFF_1176.CK  = CK;
  assign \DFF_1176.D  = \DFF_1100.Q ;
  assign \DFF_1177.CK  = CK;
  assign \DFF_1178.CK  = CK;
  assign \DFF_1179.CK  = CK;
  assign \DFF_118.CK  = CK;
  assign \DFF_1180.CK  = CK;
  assign \DFF_1181.CK  = CK;
  assign \DFF_1182.CK  = CK;
  assign \DFF_1183.CK  = CK;
  assign \DFF_1184.CK  = CK;
  assign \DFF_1185.CK  = CK;
  assign \DFF_1185.D  = \DFF_1248.Q ;
  assign \DFF_1186.CK  = CK;
  assign \DFF_1187.CK  = CK;
  assign \DFF_1188.CK  = CK;
  assign \DFF_1189.CK  = CK;
  assign \DFF_119.CK  = CK;
  assign \DFF_1190.CK  = CK;
  assign \DFF_1191.CK  = CK;
  assign \DFF_1191.D  = \DFF_1118.Q ;
  assign \DFF_1192.CK  = CK;
  assign \DFF_1193.CK  = CK;
  assign \DFF_1194.CK  = CK;
  assign \DFF_1195.CK  = CK;
  assign \DFF_1196.CK  = CK;
  assign \DFF_1196.D  = \DFF_806.Q ;
  assign \DFF_1197.CK  = CK;
  assign \DFF_1198.CK  = CK;
  assign \DFF_1199.CK  = CK;
  assign \DFF_12.CK  = CK;
  assign \DFF_120.CK  = CK;
  assign \DFF_1200.CK  = CK;
  assign \DFF_1201.CK  = CK;
  assign \DFF_1202.CK  = CK;
  assign \DFF_1203.CK  = CK;
  assign \DFF_1204.CK  = CK;
  assign \DFF_1205.CK  = CK;
  assign \DFF_1206.CK  = CK;
  assign \DFF_1207.CK  = CK;
  assign \DFF_1208.CK  = CK;
  assign \DFF_1209.CK  = CK;
  assign \DFF_1209.D  = \DFF_991.Q ;
  assign \DFF_121.CK  = CK;
  assign \DFF_1210.CK  = CK;
  assign \DFF_1211.CK  = CK;
  assign \DFF_1212.CK  = CK;
  assign \DFF_1213.CK  = CK;
  assign \DFF_1214.CK  = CK;
  assign \DFF_1215.CK  = CK;
  assign \DFF_1216.CK  = CK;
  assign \DFF_1217.CK  = CK;
  assign \DFF_1218.CK  = CK;
  assign \DFF_1219.CK  = CK;
  assign \DFF_1219.D  = \DFF_662.Q ;
  assign \DFF_122.CK  = CK;
  assign \DFF_1220.CK  = CK;
  assign \DFF_1221.CK  = CK;
  assign \DFF_1222.CK  = CK;
  assign \DFF_1223.CK  = CK;
  assign \DFF_1224.CK  = CK;
  assign \DFF_1224.D  = \DFF_565.Q ;
  assign \DFF_1225.CK  = CK;
  assign \DFF_1226.CK  = CK;
  assign \DFF_1227.CK  = CK;
  assign \DFF_1228.CK  = CK;
  assign \DFF_1228.D  = \DFF_545.Q ;
  assign \DFF_1229.CK  = CK;
  assign \DFF_123.CK  = CK;
  assign \DFF_123.D  = \DFF_315.Q ;
  assign \DFF_1230.CK  = CK;
  assign \DFF_1231.CK  = CK;
  assign \DFF_1232.CK  = CK;
  assign \DFF_1233.CK  = CK;
  assign \DFF_1234.CK  = CK;
  assign \DFF_1235.CK  = CK;
  assign \DFF_1236.CK  = CK;
  assign \DFF_1237.CK  = CK;
  assign \DFF_1238.CK  = CK;
  assign \DFF_1239.CK  = CK;
  assign \DFF_124.CK  = CK;
  assign \DFF_1240.CK  = CK;
  assign \DFF_1241.CK  = CK;
  assign \DFF_1242.CK  = CK;
  assign \DFF_1243.CK  = CK;
  assign \DFF_1244.CK  = CK;
  assign \DFF_1245.CK  = CK;
  assign \DFF_1246.CK  = CK;
  assign \DFF_1247.CK  = CK;
  assign \DFF_1248.CK  = CK;
  assign \DFF_1248.D  = \DFF_1196.Q ;
  assign \DFF_1249.CK  = CK;
  assign \DFF_125.CK  = CK;
  assign \DFF_1250.CK  = CK;
  assign \DFF_1251.CK  = CK;
  assign \DFF_1252.CK  = CK;
  assign \DFF_1253.CK  = CK;
  assign \DFF_1254.CK  = CK;
  assign \DFF_1255.CK  = CK;
  assign \DFF_1256.CK  = CK;
  assign \DFF_1257.CK  = CK;
  assign \DFF_1258.CK  = CK;
  assign \DFF_1259.CK  = CK;
  assign \DFF_126.CK  = CK;
  assign \DFF_1260.CK  = CK;
  assign \DFF_1261.CK  = CK;
  assign \DFF_1262.CK  = CK;
  assign \DFF_1262.D  = \DFF_695.Q ;
  assign \DFF_1263.CK  = CK;
  assign \DFF_1264.CK  = CK;
  assign \DFF_1265.CK  = CK;
  assign \DFF_1266.CK  = CK;
  assign \DFF_1267.CK  = CK;
  assign \DFF_1268.CK  = CK;
  assign \DFF_1269.CK  = CK;
  assign \DFF_127.CK  = CK;
  assign \DFF_1270.CK  = CK;
  assign \DFF_1271.CK  = CK;
  assign \DFF_1272.CK  = CK;
  assign \DFF_1273.CK  = CK;
  assign \DFF_1274.CK  = CK;
  assign \DFF_1275.CK  = CK;
  assign \DFF_1276.CK  = CK;
  assign \DFF_1277.CK  = CK;
  assign \DFF_1278.CK  = CK;
  assign \DFF_1279.CK  = CK;
  assign \DFF_128.CK  = CK;
  assign \DFF_1280.CK  = CK;
  assign \DFF_1281.CK  = CK;
  assign \DFF_1282.CK  = CK;
  assign \DFF_1283.CK  = CK;
  assign \DFF_1284.CK  = CK;
  assign \DFF_1285.CK  = CK;
  assign \DFF_1286.CK  = CK;
  assign \DFF_1286.D  = \DFF_389.Q ;
  assign \DFF_1287.CK  = CK;
  assign \DFF_1288.CK  = CK;
  assign \DFF_1289.CK  = CK;
  assign \DFF_129.CK  = CK;
  assign \DFF_1290.CK  = CK;
  assign \DFF_1291.CK  = CK;
  assign \DFF_1292.CK  = CK;
  assign \DFF_1293.CK  = CK;
  assign \DFF_1293.D  = \DFF_1038.Q ;
  assign \DFF_1294.CK  = CK;
  assign \DFF_1295.CK  = CK;
  assign \DFF_1296.CK  = CK;
  assign \DFF_1297.CK  = CK;
  assign \DFF_1298.CK  = CK;
  assign \DFF_1299.CK  = CK;
  assign \DFF_13.CK  = CK;
  assign \DFF_130.CK  = CK;
  assign \DFF_1300.CK  = CK;
  assign \DFF_1300.D  = \DFF_369.Q ;
  assign \DFF_1301.CK  = CK;
  assign \DFF_1302.CK  = CK;
  assign \DFF_1303.CK  = CK;
  assign \DFF_1303.D  = \DFF_1359.Q ;
  assign \DFF_1304.CK  = CK;
  assign \DFF_1305.CK  = CK;
  assign \DFF_1306.CK  = CK;
  assign \DFF_1307.CK  = CK;
  assign \DFF_1308.CK  = CK;
  assign \DFF_1308.D  = \DFF_675.Q ;
  assign \DFF_1309.CK  = CK;
  assign \DFF_131.CK  = CK;
  assign \DFF_1310.CK  = CK;
  assign \DFF_1311.CK  = CK;
  assign \DFF_1312.CK  = CK;
  assign \DFF_1313.CK  = CK;
  assign \DFF_1314.CK  = CK;
  assign \DFF_1315.CK  = CK;
  assign \DFF_1316.CK  = CK;
  assign \DFF_1317.CK  = CK;
  assign \DFF_1318.CK  = CK;
  assign \DFF_1319.CK  = CK;
  assign \DFF_132.CK  = CK;
  assign \DFF_1320.CK  = CK;
  assign \DFF_1321.CK  = CK;
  assign \DFF_1322.CK  = CK;
  assign \DFF_1323.CK  = CK;
  assign \DFF_1324.CK  = CK;
  assign \DFF_1325.CK  = CK;
  assign \DFF_1326.CK  = CK;
  assign \DFF_1327.CK  = CK;
  assign \DFF_1328.CK  = CK;
  assign \DFF_1329.CK  = CK;
  assign \DFF_133.CK  = CK;
  assign \DFF_1330.CK  = CK;
  assign \DFF_1331.CK  = CK;
  assign \DFF_1332.CK  = CK;
  assign \DFF_1333.CK  = CK;
  assign \DFF_1334.CK  = CK;
  assign \DFF_1335.CK  = CK;
  assign \DFF_1335.D  = \DFF_46.Q ;
  assign \DFF_1336.CK  = CK;
  assign \DFF_1337.CK  = CK;
  assign \DFF_1338.CK  = CK;
  assign \DFF_1338.D  = \DFF_944.Q ;
  assign \DFF_1339.CK  = CK;
  assign \DFF_134.CK  = CK;
  assign \DFF_1340.CK  = CK;
  assign \DFF_1341.CK  = CK;
  assign \DFF_1342.CK  = CK;
  assign \DFF_1343.CK  = CK;
  assign \DFF_1344.CK  = CK;
  assign \DFF_1345.CK  = CK;
  assign \DFF_1346.CK  = CK;
  assign \DFF_1347.CK  = CK;
  assign \DFF_1348.CK  = CK;
  assign \DFF_1349.CK  = CK;
  assign \DFF_135.CK  = CK;
  assign \DFF_1350.CK  = CK;
  assign \DFF_1351.CK  = CK;
  assign \DFF_1352.CK  = CK;
  assign \DFF_1352.D  = \DFF_101.Q ;
  assign \DFF_1353.CK  = CK;
  assign \DFF_1354.CK  = CK;
  assign \DFF_1354.D  = \DFF_1293.Q ;
  assign \DFF_1355.CK  = CK;
  assign \DFF_1356.CK  = CK;
  assign \DFF_1357.CK  = CK;
  assign \DFF_1358.CK  = CK;
  assign \DFF_1359.CK  = CK;
  assign \DFF_1359.D  = \DFF_76.Q ;
  assign \DFF_136.CK  = CK;
  assign \DFF_1360.CK  = CK;
  assign \DFF_1361.CK  = CK;
  assign \DFF_1362.CK  = CK;
  assign \DFF_1363.CK  = CK;
  assign \DFF_1364.CK  = CK;
  assign \DFF_1365.CK  = CK;
  assign \DFF_1366.CK  = CK;
  assign \DFF_1367.CK  = CK;
  assign \DFF_1368.CK  = CK;
  assign \DFF_1369.CK  = CK;
  assign \DFF_137.CK  = CK;
  assign \DFF_1370.CK  = CK;
  assign \DFF_1371.CK  = CK;
  assign \DFF_1372.CK  = CK;
  assign \DFF_1373.CK  = CK;
  assign \DFF_1374.CK  = CK;
  assign \DFF_1375.CK  = CK;
  assign \DFF_1376.CK  = CK;
  assign \DFF_1377.CK  = CK;
  assign \DFF_1378.CK  = CK;
  assign \DFF_1379.CK  = CK;
  assign \DFF_138.CK  = CK;
  assign \DFF_1380.CK  = CK;
  assign \DFF_1381.CK  = CK;
  assign \DFF_1382.CK  = CK;
  assign \DFF_1383.CK  = CK;
  assign \DFF_1384.CK  = CK;
  assign \DFF_1385.CK  = CK;
  assign \DFF_1386.CK  = CK;
  assign \DFF_1387.CK  = CK;
  assign \DFF_1388.CK  = CK;
  assign \DFF_1389.CK  = CK;
  assign \DFF_1389.D  = \DFF_704.Q ;
  assign \DFF_139.CK  = CK;
  assign \DFF_1390.CK  = CK;
  assign \DFF_1391.CK  = CK;
  assign \DFF_1392.CK  = CK;
  assign \DFF_1393.CK  = CK;
  assign \DFF_1394.CK  = CK;
  assign \DFF_1395.CK  = CK;
  assign \DFF_1396.CK  = CK;
  assign \DFF_1396.D  = \DFF_630.Q ;
  assign \DFF_1397.CK  = CK;
  assign \DFF_1398.CK  = CK;
  assign \DFF_1399.CK  = CK;
  assign \DFF_14.CK  = CK;
  assign \DFF_140.CK  = CK;
  assign \DFF_1400.CK  = CK;
  assign \DFF_1401.CK  = CK;
  assign \DFF_1402.CK  = CK;
  assign \DFF_1403.CK  = CK;
  assign \DFF_1404.CK  = CK;
  assign \DFF_1405.CK  = CK;
  assign \DFF_1406.CK  = CK;
  assign \DFF_1407.CK  = CK;
  assign \DFF_1408.CK  = CK;
  assign \DFF_1409.CK  = CK;
  assign \DFF_141.CK  = CK;
  assign \DFF_1410.CK  = CK;
  assign \DFF_1411.CK  = CK;
  assign \DFF_1412.CK  = CK;
  assign \DFF_1413.CK  = CK;
  assign \DFF_1414.CK  = CK;
  assign \DFF_1415.CK  = CK;
  assign \DFF_1416.CK  = CK;
  assign \DFF_1416.D  = \DFF_1224.Q ;
  assign \DFF_1417.CK  = CK;
  assign \DFF_1418.CK  = CK;
  assign \DFF_1419.CK  = CK;
  assign \DFF_142.CK  = CK;
  assign \DFF_1420.CK  = CK;
  assign \DFF_1421.CK  = CK;
  assign \DFF_1422.CK  = CK;
  assign \DFF_1423.CK  = CK;
  assign \DFF_1424.CK  = CK;
  assign \DFF_1425.CK  = CK;
  assign \DFF_143.CK  = CK;
  assign \DFF_144.CK  = CK;
  assign \DFF_145.CK  = CK;
  assign \DFF_146.CK  = CK;
  assign \DFF_146.D  = \DFF_422.Q ;
  assign \DFF_147.CK  = CK;
  assign \DFF_148.CK  = CK;
  assign \DFF_149.CK  = CK;
  assign \DFF_15.CK  = CK;
  assign \DFF_150.CK  = CK;
  assign \DFF_151.CK  = CK;
  assign \DFF_152.CK  = CK;
  assign \DFF_152.D  = \DFF_1106.Q ;
  assign \DFF_153.CK  = CK;
  assign \DFF_154.CK  = CK;
  assign \DFF_155.CK  = CK;
  assign \DFF_156.CK  = CK;
  assign \DFF_157.CK  = CK;
  assign \DFF_158.CK  = CK;
  assign \DFF_159.CK  = CK;
  assign \DFF_16.CK  = CK;
  assign \DFF_160.CK  = CK;
  assign \DFF_161.CK  = CK;
  assign \DFF_162.CK  = CK;
  assign \DFF_163.CK  = CK;
  assign \DFF_163.D  = \DFF_1185.Q ;
  assign \DFF_164.CK  = CK;
  assign \DFF_165.CK  = CK;
  assign \DFF_166.CK  = CK;
  assign \DFF_166.D  = \DFF_317.Q ;
  assign \DFF_167.CK  = CK;
  assign \DFF_168.CK  = CK;
  assign \DFF_168.D  = \DFF_371.Q ;
  assign \DFF_169.CK  = CK;
  assign \DFF_17.CK  = CK;
  assign \DFF_170.CK  = CK;
  assign \DFF_171.CK  = CK;
  assign \DFF_171.D  = \DFF_1072.Q ;
  assign \DFF_172.CK  = CK;
  assign \DFF_173.CK  = CK;
  assign \DFF_174.CK  = CK;
  assign \DFF_175.CK  = CK;
  assign \DFF_176.CK  = CK;
  assign \DFF_177.CK  = CK;
  assign \DFF_178.CK  = CK;
  assign \DFF_179.CK  = CK;
  assign \DFF_18.CK  = CK;
  assign \DFF_180.CK  = CK;
  assign \DFF_181.CK  = CK;
  assign \DFF_181.D  = \DFF_305.Q ;
  assign \DFF_182.CK  = CK;
  assign \DFF_183.CK  = CK;
  assign \DFF_184.CK  = CK;
  assign \DFF_185.CK  = CK;
  assign \DFF_186.CK  = CK;
  assign \DFF_187.CK  = CK;
  assign \DFF_188.CK  = CK;
  assign \DFF_188.D  = \DFF_554.Q ;
  assign \DFF_189.CK  = CK;
  assign \DFF_19.CK  = CK;
  assign \DFF_190.CK  = CK;
  assign \DFF_191.CK  = CK;
  assign \DFF_192.CK  = CK;
  assign \DFF_193.CK  = CK;
  assign \DFF_194.CK  = CK;
  assign \DFF_195.CK  = CK;
  assign \DFF_196.CK  = CK;
  assign \DFF_197.CK  = CK;
  assign \DFF_198.CK  = CK;
  assign \DFF_199.CK  = CK;
  assign \DFF_2.CK  = CK;
  assign \DFF_20.CK  = CK;
  assign \DFF_200.CK  = CK;
  assign \DFF_201.CK  = CK;
  assign \DFF_202.CK  = CK;
  assign \DFF_203.CK  = CK;
  assign \DFF_204.CK  = CK;
  assign \DFF_205.CK  = CK;
  assign \DFF_206.CK  = CK;
  assign \DFF_207.CK  = CK;
  assign \DFF_208.CK  = CK;
  assign \DFF_209.CK  = CK;
  assign \DFF_21.CK  = CK;
  assign \DFF_210.CK  = CK;
  assign \DFF_211.CK  = CK;
  assign \DFF_212.CK  = CK;
  assign \DFF_213.CK  = CK;
  assign \DFF_214.CK  = CK;
  assign \DFF_215.CK  = CK;
  assign \DFF_216.CK  = CK;
  assign \DFF_217.CK  = CK;
  assign \DFF_218.CK  = CK;
  assign \DFF_219.CK  = CK;
  assign \DFF_22.CK  = CK;
  assign \DFF_22.D  = \DFF_279.Q ;
  assign \DFF_220.CK  = CK;
  assign \DFF_220.D  = \DFF_942.Q ;
  assign \DFF_221.CK  = CK;
  assign \DFF_222.CK  = CK;
  assign \DFF_223.CK  = CK;
  assign \DFF_224.CK  = CK;
  assign \DFF_225.CK  = CK;
  assign \DFF_226.CK  = CK;
  assign \DFF_227.CK  = CK;
  assign \DFF_228.CK  = CK;
  assign \DFF_229.CK  = CK;
  assign \DFF_23.CK  = CK;
  assign \DFF_230.CK  = CK;
  assign \DFF_231.CK  = CK;
  assign \DFF_232.CK  = CK;
  assign \DFF_233.CK  = CK;
  assign \DFF_234.CK  = CK;
  assign \DFF_235.CK  = CK;
  assign \DFF_235.D  = \DFF_85.Q ;
  assign \DFF_236.CK  = CK;
  assign \DFF_237.CK  = CK;
  assign \DFF_238.CK  = CK;
  assign \DFF_239.CK  = CK;
  assign \DFF_24.CK  = CK;
  assign \DFF_240.CK  = CK;
  assign \DFF_241.CK  = CK;
  assign \DFF_242.CK  = CK;
  assign \DFF_243.CK  = CK;
  assign \DFF_244.CK  = CK;
  assign \DFF_245.CK  = CK;
  assign \DFF_246.CK  = CK;
  assign \DFF_247.CK  = CK;
  assign \DFF_248.CK  = CK;
  assign \DFF_249.CK  = CK;
  assign \DFF_25.CK  = CK;
  assign \DFF_250.CK  = CK;
  assign \DFF_251.CK  = CK;
  assign \DFF_252.CK  = CK;
  assign \DFF_253.CK  = CK;
  assign \DFF_254.CK  = CK;
  assign \DFF_255.CK  = CK;
  assign \DFF_256.CK  = CK;
  assign \DFF_256.D  = \DFF_1081.Q ;
  assign \DFF_257.CK  = CK;
  assign \DFF_258.CK  = CK;
  assign \DFF_259.CK  = CK;
  assign \DFF_26.CK  = CK;
  assign \DFF_260.CK  = CK;
  assign \DFF_261.CK  = CK;
  assign \DFF_262.CK  = CK;
  assign \DFF_263.CK  = CK;
  assign \DFF_263.D  = \DFF_117.Q ;
  assign \DFF_264.CK  = CK;
  assign \DFF_265.CK  = CK;
  assign \DFF_266.CK  = CK;
  assign \DFF_267.CK  = CK;
  assign \DFF_268.CK  = CK;
  assign \DFF_269.CK  = CK;
  assign \DFF_27.CK  = CK;
  assign \DFF_270.CK  = CK;
  assign \DFF_271.CK  = CK;
  assign \DFF_272.CK  = CK;
  assign \DFF_273.CK  = CK;
  assign \DFF_274.CK  = CK;
  assign \DFF_275.CK  = CK;
  assign \DFF_276.CK  = CK;
  assign \DFF_277.CK  = CK;
  assign \DFF_278.CK  = CK;
  assign \DFF_279.CK  = CK;
  assign \DFF_279.D  = \DFF_1102.Q ;
  assign \DFF_28.CK  = CK;
  assign \DFF_280.CK  = CK;
  assign \DFF_281.CK  = CK;
  assign \DFF_281.D  = \DFF_360.Q ;
  assign \DFF_282.CK  = CK;
  assign \DFF_283.CK  = CK;
  assign \DFF_284.CK  = CK;
  assign \DFF_285.CK  = CK;
  assign \DFF_286.CK  = CK;
  assign \DFF_287.CK  = CK;
  assign \DFF_288.CK  = CK;
  assign \DFF_289.CK  = CK;
  assign \DFF_29.CK  = CK;
  assign \DFF_290.CK  = CK;
  assign \DFF_290.D  = \DFF_1300.Q ;
  assign \DFF_291.CK  = CK;
  assign \DFF_292.CK  = CK;
  assign \DFF_293.CK  = CK;
  assign \DFF_294.CK  = CK;
  assign \DFF_295.CK  = CK;
  assign \DFF_295.D  = \DFF_1122.Q ;
  assign \DFF_296.CK  = CK;
  assign \DFF_297.CK  = CK;
  assign \DFF_298.CK  = CK;
  assign \DFF_299.CK  = CK;
  assign \DFF_299.D  = \DFF_147.Q ;
  assign \DFF_3.CK  = CK;
  assign \DFF_30.CK  = CK;
  assign \DFF_300.CK  = CK;
  assign \DFF_301.CK  = CK;
  assign \DFF_302.CK  = CK;
  assign \DFF_303.CK  = CK;
  assign \DFF_304.CK  = CK;
  assign \DFF_305.CK  = CK;
  assign \DFF_305.D  = \DFF_401.Q ;
  assign \DFF_306.CK  = CK;
  assign \DFF_307.CK  = CK;
  assign \DFF_308.CK  = CK;
  assign \DFF_309.CK  = CK;
  assign \DFF_31.CK  = CK;
  assign \DFF_31.D  = \DFF_1338.Q ;
  assign \DFF_310.CK  = CK;
  assign \DFF_311.CK  = CK;
  assign \DFF_312.CK  = CK;
  assign \DFF_313.CK  = CK;
  assign \DFF_314.CK  = CK;
  assign \DFF_315.CK  = CK;
  assign \DFF_315.D  = \DFF_474.Q ;
  assign \DFF_316.CK  = CK;
  assign \DFF_317.CK  = CK;
  assign \DFF_318.CK  = CK;
  assign \DFF_319.CK  = CK;
  assign \DFF_32.CK  = CK;
  assign \DFF_320.CK  = CK;
  assign \DFF_320.D  = \DFF_831.Q ;
  assign \DFF_321.CK  = CK;
  assign \DFF_322.CK  = CK;
  assign \DFF_323.CK  = CK;
  assign \DFF_324.CK  = CK;
  assign \DFF_325.CK  = CK;
  assign \DFF_325.D  = \DFF_739.Q ;
  assign \DFF_326.CK  = CK;
  assign \DFF_326.D  = \DFF_30.Q ;
  assign \DFF_327.CK  = CK;
  assign \DFF_327.D  = \DFF_937.Q ;
  assign \DFF_328.CK  = CK;
  assign \DFF_329.CK  = CK;
  assign \DFF_33.CK  = CK;
  assign \DFF_330.CK  = CK;
  assign \DFF_331.CK  = CK;
  assign \DFF_332.CK  = CK;
  assign \DFF_333.CK  = CK;
  assign \DFF_334.CK  = CK;
  assign \DFF_334.D  = \DFF_60.Q ;
  assign \DFF_335.CK  = CK;
  assign \DFF_336.CK  = CK;
  assign \DFF_337.CK  = CK;
  assign \DFF_338.CK  = CK;
  assign \DFF_339.CK  = CK;
  assign \DFF_34.CK  = CK;
  assign \DFF_34.D  = \DFF_81.Q ;
  assign \DFF_340.CK  = CK;
  assign \DFF_341.CK  = CK;
  assign \DFF_342.CK  = CK;
  assign \DFF_343.CK  = CK;
  assign \DFF_344.CK  = CK;
  assign \DFF_345.CK  = CK;
  assign \DFF_346.CK  = CK;
  assign \DFF_347.CK  = CK;
  assign \DFF_348.CK  = CK;
  assign \DFF_349.CK  = CK;
  assign \DFF_35.CK  = CK;
  assign \DFF_350.CK  = CK;
  assign \DFF_351.CK  = CK;
  assign \DFF_352.CK  = CK;
  assign \DFF_353.CK  = CK;
  assign \DFF_354.CK  = CK;
  assign \DFF_355.CK  = CK;
  assign \DFF_356.CK  = CK;
  assign \DFF_357.CK  = CK;
  assign \DFF_358.CK  = CK;
  assign \DFF_359.CK  = CK;
  assign \DFF_36.CK  = CK;
  assign \DFF_360.CK  = CK;
  assign \DFF_360.D  = \DFF_537.Q ;
  assign \DFF_361.CK  = CK;
  assign \DFF_362.CK  = CK;
  assign \DFF_363.CK  = CK;
  assign \DFF_364.CK  = CK;
  assign \DFF_365.CK  = CK;
  assign \DFF_365.D  = \DFF_376.Q ;
  assign \DFF_366.CK  = CK;
  assign \DFF_367.CK  = CK;
  assign \DFF_367.D  = \DFF_642.Q ;
  assign \DFF_368.CK  = CK;
  assign \DFF_369.CK  = CK;
  assign \DFF_369.D  = \DFF_873.Q ;
  assign \DFF_37.CK  = CK;
  assign \DFF_370.CK  = CK;
  assign \DFF_371.CK  = CK;
  assign \DFF_372.CK  = CK;
  assign \DFF_372.D  = \DFF_1110.Q ;
  assign \DFF_373.CK  = CK;
  assign \DFF_373.D  = \DFF_1225.Q ;
  assign \DFF_374.CK  = CK;
  assign \DFF_375.CK  = CK;
  assign \DFF_376.CK  = CK;
  assign \DFF_377.CK  = CK;
  assign \DFF_377.D  = \DFF_1316.Q ;
  assign \DFF_378.CK  = CK;
  assign \DFF_379.CK  = CK;
  assign \DFF_38.CK  = CK;
  assign \DFF_38.D  = \DFF_528.Q ;
  assign \DFF_380.CK  = CK;
  assign \DFF_380.D  = \DFF_404.Q ;
  assign \DFF_381.CK  = CK;
  assign \DFF_382.CK  = CK;
  assign \DFF_383.CK  = CK;
  assign \DFF_384.CK  = CK;
  assign \DFF_385.CK  = CK;
  assign \DFF_386.CK  = CK;
  assign \DFF_387.CK  = CK;
  assign \DFF_388.CK  = CK;
  assign \DFF_389.CK  = CK;
  assign \DFF_39.CK  = CK;
  assign \DFF_390.CK  = CK;
  assign \DFF_391.CK  = CK;
  assign \DFF_392.CK  = CK;
  assign \DFF_393.CK  = CK;
  assign \DFF_394.CK  = CK;
  assign \DFF_395.CK  = CK;
  assign \DFF_396.CK  = CK;
  assign \DFF_397.CK  = CK;
  assign \DFF_398.CK  = CK;
  assign \DFF_399.CK  = CK;
  assign \DFF_4.CK  = CK;
  assign \DFF_40.CK  = CK;
  assign \DFF_400.CK  = CK;
  assign \DFF_401.CK  = CK;
  assign \DFF_401.D  = \DFF_1001.Q ;
  assign \DFF_402.CK  = CK;
  assign \DFF_403.CK  = CK;
  assign \DFF_404.CK  = CK;
  assign \DFF_404.D  = \DFF_152.Q ;
  assign \DFF_405.CK  = CK;
  assign \DFF_406.CK  = CK;
  assign \DFF_407.CK  = CK;
  assign \DFF_408.CK  = CK;
  assign \DFF_408.D  = \DFF_334.Q ;
  assign \DFF_409.CK  = CK;
  assign \DFF_41.CK  = CK;
  assign \DFF_410.CK  = CK;
  assign \DFF_411.CK  = CK;
  assign \DFF_412.CK  = CK;
  assign \DFF_413.CK  = CK;
  assign \DFF_414.CK  = CK;
  assign \DFF_415.CK  = CK;
  assign \DFF_416.CK  = CK;
  assign \DFF_417.CK  = CK;
  assign \DFF_418.CK  = CK;
  assign \DFF_418.D  = \DFF_885.Q ;
  assign \DFF_419.CK  = CK;
  assign \DFF_42.CK  = CK;
  assign \DFF_420.CK  = CK;
  assign \DFF_421.CK  = CK;
  assign \DFF_422.CK  = CK;
  assign \DFF_423.CK  = CK;
  assign \DFF_424.CK  = CK;
  assign \DFF_425.CK  = CK;
  assign \DFF_426.CK  = CK;
  assign \DFF_427.CK  = CK;
  assign \DFF_428.CK  = CK;
  assign \DFF_429.CK  = CK;
  assign \DFF_43.CK  = CK;
  assign \DFF_430.CK  = CK;
  assign \DFF_431.CK  = CK;
  assign \DFF_432.CK  = CK;
  assign \DFF_433.CK  = CK;
  assign \DFF_434.CK  = CK;
  assign \DFF_435.CK  = CK;
  assign \DFF_436.CK  = CK;
  assign \DFF_437.CK  = CK;
  assign \DFF_438.CK  = CK;
  assign \DFF_439.CK  = CK;
  assign \DFF_44.CK  = CK;
  assign \DFF_440.CK  = CK;
  assign \DFF_441.CK  = CK;
  assign \DFF_442.CK  = CK;
  assign \DFF_443.CK  = CK;
  assign \DFF_444.CK  = CK;
  assign \DFF_445.CK  = CK;
  assign \DFF_446.CK  = CK;
  assign \DFF_447.CK  = CK;
  assign \DFF_448.CK  = CK;
  assign \DFF_449.CK  = CK;
  assign \DFF_45.CK  = CK;
  assign \DFF_450.CK  = CK;
  assign \DFF_450.D  = \DFF_460.Q ;
  assign \DFF_451.CK  = CK;
  assign \DFF_452.CK  = CK;
  assign \DFF_453.CK  = CK;
  assign \DFF_454.CK  = CK;
  assign \DFF_455.CK  = CK;
  assign \DFF_456.CK  = CK;
  assign \DFF_457.CK  = CK;
  assign \DFF_458.CK  = CK;
  assign \DFF_458.D  = \DFF_678.Q ;
  assign \DFF_459.CK  = CK;
  assign \DFF_46.CK  = CK;
  assign \DFF_460.CK  = CK;
  assign \DFF_461.CK  = CK;
  assign \DFF_462.CK  = CK;
  assign \DFF_463.CK  = CK;
  assign \DFF_464.CK  = CK;
  assign \DFF_465.CK  = CK;
  assign \DFF_466.CK  = CK;
  assign \DFF_467.CK  = CK;
  assign \DFF_468.CK  = CK;
  assign \DFF_468.D  = \DFF_1420.Q ;
  assign \DFF_469.CK  = CK;
  assign \DFF_47.CK  = CK;
  assign \DFF_470.CK  = CK;
  assign \DFF_471.CK  = CK;
  assign \DFF_472.CK  = CK;
  assign \DFF_473.CK  = CK;
  assign \DFF_474.CK  = CK;
  assign \DFF_474.D  = \DFF_188.Q ;
  assign \DFF_475.CK  = CK;
  assign \DFF_476.CK  = CK;
  assign \DFF_477.CK  = CK;
  assign \DFF_478.CK  = CK;
  assign \DFF_479.CK  = CK;
  assign \DFF_48.CK  = CK;
  assign \DFF_480.CK  = CK;
  assign \DFF_480.D  = \DFF_1234.Q ;
  assign \DFF_481.CK  = CK;
  assign \DFF_481.D  = \DFF_1275.Q ;
  assign \DFF_482.CK  = CK;
  assign \DFF_483.CK  = CK;
  assign \DFF_484.CK  = CK;
  assign \DFF_485.CK  = CK;
  assign \DFF_485.D  = \DFF_1286.Q ;
  assign \DFF_486.CK  = CK;
  assign \DFF_487.CK  = CK;
  assign \DFF_488.CK  = CK;
  assign \DFF_489.CK  = CK;
  assign \DFF_49.CK  = CK;
  assign \DFF_490.CK  = CK;
  assign \DFF_491.CK  = CK;
  assign \DFF_492.CK  = CK;
  assign \DFF_492.D  = \DFF_1414.Q ;
  assign \DFF_493.CK  = CK;
  assign \DFF_494.CK  = CK;
  assign \DFF_495.CK  = CK;
  assign \DFF_496.CK  = CK;
  assign \DFF_497.CK  = CK;
  assign \DFF_498.CK  = CK;
  assign \DFF_499.CK  = CK;
  assign \DFF_5.CK  = CK;
  assign \DFF_50.CK  = CK;
  assign \DFF_500.CK  = CK;
  assign \DFF_501.CK  = CK;
  assign \DFF_502.CK  = CK;
  assign \DFF_503.CK  = CK;
  assign \DFF_504.CK  = CK;
  assign \DFF_505.CK  = CK;
  assign \DFF_506.CK  = CK;
  assign \DFF_507.CK  = CK;
  assign \DFF_508.CK  = CK;
  assign \DFF_509.CK  = CK;
  assign \DFF_509.D  = \DFF_203.Q ;
  assign \DFF_51.CK  = CK;
  assign \DFF_510.CK  = CK;
  assign \DFF_511.CK  = CK;
  assign \DFF_511.D  = \DFF_1308.Q ;
  assign \DFF_512.CK  = CK;
  assign \DFF_513.CK  = CK;
  assign \DFF_514.CK  = CK;
  assign \DFF_515.CK  = CK;
  assign \DFF_516.CK  = CK;
  assign \DFF_517.CK  = CK;
  assign \DFF_518.CK  = CK;
  assign \DFF_519.CK  = CK;
  assign \DFF_52.CK  = CK;
  assign \DFF_520.CK  = CK;
  assign \DFF_521.CK  = CK;
  assign \DFF_522.CK  = CK;
  assign \DFF_523.CK  = CK;
  assign \DFF_524.CK  = CK;
  assign \DFF_525.CK  = CK;
  assign \DFF_526.CK  = CK;
  assign \DFF_527.CK  = CK;
  assign \DFF_528.CK  = CK;
  assign \DFF_528.D  = \DFF_1362.Q ;
  assign \DFF_529.CK  = CK;
  assign \DFF_529.D  = \DFF_819.Q ;
  assign \DFF_53.CK  = CK;
  assign \DFF_53.D  = \DFF_898.Q ;
  assign \DFF_530.CK  = CK;
  assign \DFF_531.CK  = CK;
  assign \DFF_532.CK  = CK;
  assign \DFF_533.CK  = CK;
  assign \DFF_534.CK  = CK;
  assign \DFF_535.CK  = CK;
  assign \DFF_536.CK  = CK;
  assign \DFF_537.CK  = CK;
  assign \DFF_537.D  = \DFF_765.Q ;
  assign \DFF_538.CK  = CK;
  assign \DFF_539.CK  = CK;
  assign \DFF_54.CK  = CK;
  assign \DFF_540.CK  = CK;
  assign \DFF_541.CK  = CK;
  assign \DFF_542.CK  = CK;
  assign \DFF_543.CK  = CK;
  assign \DFF_544.CK  = CK;
  assign \DFF_545.CK  = CK;
  assign \DFF_546.CK  = CK;
  assign \DFF_547.CK  = CK;
  assign \DFF_548.CK  = CK;
  assign \DFF_549.CK  = CK;
  assign \DFF_55.CK  = CK;
  assign \DFF_550.CK  = CK;
  assign \DFF_551.CK  = CK;
  assign \DFF_552.CK  = CK;
  assign \DFF_553.CK  = CK;
  assign \DFF_553.D  = \DFF_86.Q ;
  assign \DFF_554.CK  = CK;
  assign \DFF_555.CK  = CK;
  assign \DFF_556.CK  = CK;
  assign \DFF_557.CK  = CK;
  assign \DFF_558.CK  = CK;
  assign \DFF_559.CK  = CK;
  assign \DFF_56.CK  = CK;
  assign \DFF_560.CK  = CK;
  assign \DFF_561.CK  = CK;
  assign \DFF_561.D  = \DFF_585.Q ;
  assign \DFF_562.CK  = CK;
  assign \DFF_563.CK  = CK;
  assign \DFF_564.CK  = CK;
  assign \DFF_565.CK  = CK;
  assign \DFF_565.D  = \DFF_909.Q ;
  assign \DFF_566.CK  = CK;
  assign \DFF_566.D  = \DFF_906.Q ;
  assign \DFF_567.CK  = CK;
  assign \DFF_568.CK  = CK;
  assign \DFF_569.CK  = CK;
  assign \DFF_569.D  = \DFF_503.Q ;
  assign \DFF_57.CK  = CK;
  assign \DFF_570.CK  = CK;
  assign \DFF_571.CK  = CK;
  assign \DFF_572.CK  = CK;
  assign \DFF_573.CK  = CK;
  assign \DFF_574.CK  = CK;
  assign \DFF_575.CK  = CK;
  assign \DFF_576.CK  = CK;
  assign \DFF_577.CK  = CK;
  assign \DFF_578.CK  = CK;
  assign \DFF_579.CK  = CK;
  assign \DFF_58.CK  = CK;
  assign \DFF_580.CK  = CK;
  assign \DFF_581.CK  = CK;
  assign \DFF_582.CK  = CK;
  assign \DFF_583.CK  = CK;
  assign \DFF_584.CK  = CK;
  assign \DFF_585.CK  = CK;
  assign \DFF_586.CK  = CK;
  assign \DFF_587.CK  = CK;
  assign \DFF_588.CK  = CK;
  assign \DFF_589.CK  = CK;
  assign \DFF_59.CK  = CK;
  assign \DFF_590.CK  = CK;
  assign \DFF_591.CK  = CK;
  assign \DFF_592.CK  = CK;
  assign \DFF_593.CK  = CK;
  assign \DFF_594.CK  = CK;
  assign \DFF_595.CK  = CK;
  assign \DFF_596.CK  = CK;
  assign \DFF_597.CK  = CK;
  assign \DFF_598.CK  = CK;
  assign \DFF_599.CK  = CK;
  assign \DFF_6.CK  = CK;
  assign \DFF_60.CK  = CK;
  assign \DFF_600.CK  = CK;
  assign \DFF_600.D  = \DFF_1207.Q ;
  assign \DFF_601.CK  = CK;
  assign \DFF_602.CK  = CK;
  assign \DFF_603.CK  = CK;
  assign \DFF_603.D  = \DFF_861.Q ;
  assign \DFF_604.CK  = CK;
  assign \DFF_605.CK  = CK;
  assign \DFF_606.CK  = CK;
  assign \DFF_607.CK  = CK;
  assign \DFF_608.CK  = CK;
  assign \DFF_609.CK  = CK;
  assign \DFF_61.CK  = CK;
  assign \DFF_610.CK  = CK;
  assign \DFF_611.CK  = CK;
  assign \DFF_612.CK  = CK;
  assign \DFF_613.CK  = CK;
  assign \DFF_613.D  = \DFF_234.Q ;
  assign \DFF_614.CK  = CK;
  assign \DFF_615.CK  = CK;
  assign \DFF_615.D  = \DFF_549.Q ;
  assign \DFF_616.CK  = CK;
  assign \DFF_616.D  = \DFF_566.Q ;
  assign \DFF_617.CK  = CK;
  assign \DFF_618.CK  = CK;
  assign \DFF_619.CK  = CK;
  assign \DFF_62.CK  = CK;
  assign \DFF_620.CK  = CK;
  assign \DFF_621.CK  = CK;
  assign \DFF_622.CK  = CK;
  assign \DFF_623.CK  = CK;
  assign \DFF_624.CK  = CK;
  assign \DFF_625.CK  = CK;
  assign \DFF_626.CK  = CK;
  assign \DFF_627.CK  = CK;
  assign \DFF_628.CK  = CK;
  assign \DFF_629.CK  = CK;
  assign \DFF_63.CK  = CK;
  assign \DFF_630.CK  = CK;
  assign \DFF_631.CK  = CK;
  assign \DFF_632.CK  = CK;
  assign \DFF_633.CK  = CK;
  assign \DFF_634.CK  = CK;
  assign \DFF_635.CK  = CK;
  assign \DFF_636.CK  = CK;
  assign \DFF_637.CK  = CK;
  assign \DFF_638.CK  = CK;
  assign \DFF_639.CK  = CK;
  assign \DFF_64.CK  = CK;
  assign \DFF_640.CK  = CK;
  assign \DFF_641.CK  = CK;
  assign \DFF_642.CK  = CK;
  assign \DFF_642.D  = \DFF_785.Q ;
  assign \DFF_643.CK  = CK;
  assign \DFF_643.D  = \DFF_711.Q ;
  assign \DFF_644.CK  = CK;
  assign \DFF_645.CK  = CK;
  assign \DFF_646.CK  = CK;
  assign \DFF_647.CK  = CK;
  assign \DFF_648.CK  = CK;
  assign \DFF_649.CK  = CK;
  assign \DFF_65.CK  = CK;
  assign \DFF_650.CK  = CK;
  assign \DFF_650.D  = g6752;
  assign \DFF_651.CK  = CK;
  assign \DFF_652.CK  = CK;
  assign \DFF_653.CK  = CK;
  assign \DFF_654.CK  = CK;
  assign \DFF_655.CK  = CK;
  assign \DFF_655.D  = \DFF_165.Q ;
  assign \DFF_656.CK  = CK;
  assign \DFF_657.CK  = CK;
  assign \DFF_658.CK  = CK;
  assign \DFF_659.CK  = CK;
  assign \DFF_66.CK  = CK;
  assign \DFF_660.CK  = CK;
  assign \DFF_661.CK  = CK;
  assign \DFF_662.CK  = CK;
  assign \DFF_662.D  = \DFF_367.Q ;
  assign \DFF_663.CK  = CK;
  assign \DFF_663.D  = \DFF_1265.Q ;
  assign \DFF_664.CK  = CK;
  assign \DFF_665.CK  = CK;
  assign \DFF_666.CK  = CK;
  assign \DFF_666.D  = \DFF_783.Q ;
  assign \DFF_667.CK  = CK;
  assign \DFF_668.CK  = CK;
  assign \DFF_669.CK  = CK;
  assign \DFF_67.CK  = CK;
  assign \DFF_670.CK  = CK;
  assign \DFF_671.CK  = CK;
  assign \DFF_672.CK  = CK;
  assign \DFF_673.CK  = CK;
  assign \DFF_674.CK  = CK;
  assign \DFF_675.CK  = CK;
  assign \DFF_676.CK  = CK;
  assign \DFF_677.CK  = CK;
  assign \DFF_678.CK  = CK;
  assign \DFF_679.CK  = CK;
  assign \DFF_68.CK  = CK;
  assign \DFF_680.CK  = CK;
  assign \DFF_681.CK  = CK;
  assign \DFF_682.CK  = CK;
  assign \DFF_683.CK  = CK;
  assign \DFF_684.CK  = CK;
  assign \DFF_685.CK  = CK;
  assign \DFF_686.CK  = CK;
  assign \DFF_687.CK  = CK;
  assign \DFF_687.D  = \DFF_348.Q ;
  assign \DFF_688.CK  = CK;
  assign \DFF_689.CK  = CK;
  assign \DFF_69.CK  = CK;
  assign \DFF_690.CK  = CK;
  assign \DFF_691.CK  = CK;
  assign \DFF_692.CK  = CK;
  assign \DFF_693.CK  = CK;
  assign \DFF_694.CK  = CK;
  assign \DFF_695.CK  = CK;
  assign \DFF_695.D  = \DFF_1352.Q ;
  assign \DFF_696.CK  = CK;
  assign \DFF_697.CK  = CK;
  assign \DFF_698.CK  = CK;
  assign \DFF_698.D  = \DFF_600.Q ;
  assign \DFF_699.CK  = CK;
  assign \DFF_7.CK  = CK;
  assign \DFF_7.D  = \DFF_109.Q ;
  assign \DFF_70.CK  = CK;
  assign \DFF_700.CK  = CK;
  assign \DFF_701.CK  = CK;
  assign \DFF_702.CK  = CK;
  assign \DFF_703.CK  = CK;
  assign \DFF_704.CK  = CK;
  assign \DFF_704.D  = \DFF_1049.Q ;
  assign \DFF_705.CK  = CK;
  assign \DFF_706.CK  = CK;
  assign \DFF_707.CK  = CK;
  assign \DFF_708.CK  = CK;
  assign \DFF_709.CK  = CK;
  assign \DFF_71.CK  = CK;
  assign \DFF_710.CK  = CK;
  assign \DFF_711.CK  = CK;
  assign \DFF_712.CK  = CK;
  assign \DFF_713.CK  = CK;
  assign \DFF_714.CK  = CK;
  assign \DFF_715.CK  = CK;
  assign \DFF_716.CK  = CK;
  assign \DFF_717.CK  = CK;
  assign \DFF_718.CK  = CK;
  assign \DFF_719.CK  = CK;
  assign \DFF_72.CK  = CK;
  assign \DFF_720.CK  = CK;
  assign \DFF_721.CK  = CK;
  assign \DFF_722.CK  = CK;
  assign \DFF_723.CK  = CK;
  assign \DFF_724.CK  = CK;
  assign \DFF_725.CK  = CK;
  assign \DFF_726.CK  = CK;
  assign \DFF_727.CK  = CK;
  assign \DFF_728.CK  = CK;
  assign \DFF_729.CK  = CK;
  assign \DFF_73.CK  = CK;
  assign \DFF_730.CK  = CK;
  assign \DFF_731.CK  = CK;
  assign \DFF_732.CK  = CK;
  assign \DFF_733.CK  = CK;
  assign \DFF_734.CK  = CK;
  assign \DFF_735.CK  = CK;
  assign \DFF_736.CK  = CK;
  assign \DFF_737.CK  = CK;
  assign \DFF_737.D  = \DFF_110.Q ;
  assign \DFF_738.CK  = CK;
  assign \DFF_739.CK  = CK;
  assign \DFF_74.CK  = CK;
  assign \DFF_740.CK  = CK;
  assign \DFF_741.CK  = CK;
  assign \DFF_742.CK  = CK;
  assign \DFF_743.CK  = CK;
  assign \DFF_744.CK  = CK;
  assign \DFF_745.CK  = CK;
  assign \DFF_746.CK  = CK;
  assign \DFF_747.CK  = CK;
  assign \DFF_748.CK  = CK;
  assign \DFF_749.CK  = CK;
  assign \DFF_75.CK  = CK;
  assign \DFF_750.CK  = CK;
  assign \DFF_751.CK  = CK;
  assign \DFF_752.CK  = CK;
  assign \DFF_753.CK  = CK;
  assign \DFF_754.CK  = CK;
  assign \DFF_755.CK  = CK;
  assign \DFF_756.CK  = CK;
  assign \DFF_757.CK  = CK;
  assign \DFF_758.CK  = CK;
  assign \DFF_759.CK  = CK;
  assign \DFF_76.CK  = CK;
  assign \DFF_76.D  = \DFF_856.Q ;
  assign \DFF_760.CK  = CK;
  assign \DFF_761.CK  = CK;
  assign \DFF_762.CK  = CK;
  assign \DFF_763.CK  = CK;
  assign \DFF_764.CK  = CK;
  assign \DFF_764.D  = \DFF_380.Q ;
  assign \DFF_765.CK  = CK;
  assign \DFF_765.D  = \DFF_616.Q ;
  assign \DFF_766.CK  = CK;
  assign \DFF_767.CK  = CK;
  assign \DFF_768.CK  = CK;
  assign \DFF_769.CK  = CK;
  assign \DFF_77.CK  = CK;
  assign \DFF_770.CK  = CK;
  assign \DFF_771.CK  = CK;
  assign \DFF_772.CK  = CK;
  assign \DFF_773.CK  = CK;
  assign \DFF_774.CK  = CK;
  assign \DFF_775.CK  = CK;
  assign \DFF_776.CK  = CK;
  assign \DFF_777.CK  = CK;
  assign \DFF_778.CK  = CK;
  assign \DFF_779.CK  = CK;
  assign \DFF_78.CK  = CK;
  assign \DFF_780.CK  = CK;
  assign \DFF_780.D  = \DFF_836.Q ;
  assign \DFF_781.CK  = CK;
  assign \DFF_782.CK  = CK;
  assign \DFF_783.CK  = CK;
  assign \DFF_783.D  = \DFF_1262.Q ;
  assign \DFF_784.CK  = CK;
  assign \DFF_785.CK  = CK;
  assign \DFF_785.D  = \DFF_181.Q ;
  assign \DFF_786.CK  = CK;
  assign \DFF_787.CK  = CK;
  assign \DFF_788.CK  = CK;
  assign \DFF_789.CK  = CK;
  assign \DFF_79.CK  = CK;
  assign \DFF_790.CK  = CK;
  assign \DFF_791.CK  = CK;
  assign \DFF_791.D  = \DFF_185.Q ;
  assign \DFF_792.CK  = CK;
  assign \DFF_793.CK  = CK;
  assign \DFF_794.CK  = CK;
  assign \DFF_795.CK  = CK;
  assign \DFF_796.CK  = CK;
  assign \DFF_797.CK  = CK;
  assign \DFF_797.D  = \DFF_326.Q ;
  assign \DFF_798.CK  = CK;
  assign \DFF_798.D  = \DFF_269.Q ;
  assign \DFF_799.CK  = CK;
  assign \DFF_8.CK  = CK;
  assign \DFF_80.CK  = CK;
  assign \DFF_800.CK  = CK;
  assign \DFF_801.CK  = CK;
  assign \DFF_802.CK  = CK;
  assign \DFF_803.CK  = CK;
  assign \DFF_804.CK  = CK;
  assign \DFF_805.CK  = CK;
  assign \DFF_806.CK  = CK;
  assign \DFF_806.D  = \DFF_1158.Q ;
  assign \DFF_807.CK  = CK;
  assign \DFF_808.CK  = CK;
  assign \DFF_809.CK  = CK;
  assign \DFF_81.CK  = CK;
  assign \DFF_81.D  = \DFF_220.Q ;
  assign \DFF_810.CK  = CK;
  assign \DFF_810.D  = \DFF_830.Q ;
  assign \DFF_811.CK  = CK;
  assign \DFF_812.CK  = CK;
  assign \DFF_813.CK  = CK;
  assign \DFF_814.CK  = CK;
  assign \DFF_815.CK  = CK;
  assign \DFF_816.CK  = CK;
  assign \DFF_817.CK  = CK;
  assign \DFF_817.D  = \DFF_1256.Q ;
  assign \DFF_818.CK  = CK;
  assign \DFF_819.CK  = CK;
  assign \DFF_82.CK  = CK;
  assign \DFF_820.CK  = CK;
  assign \DFF_821.CK  = CK;
  assign \DFF_822.CK  = CK;
  assign \DFF_823.CK  = CK;
  assign \DFF_824.CK  = CK;
  assign \DFF_825.CK  = CK;
  assign \DFF_826.CK  = CK;
  assign \DFF_827.CK  = CK;
  assign \DFF_828.CK  = CK;
  assign \DFF_828.D  = \DFF_339.Q ;
  assign \DFF_829.CK  = CK;
  assign \DFF_83.CK  = CK;
  assign \DFF_830.CK  = CK;
  assign \DFF_831.CK  = CK;
  assign \DFF_832.CK  = CK;
  assign \DFF_833.CK  = CK;
  assign \DFF_834.CK  = CK;
  assign \DFF_835.CK  = CK;
  assign \DFF_836.CK  = CK;
  assign \DFF_836.D  = \DFF_971.Q ;
  assign \DFF_837.CK  = CK;
  assign \DFF_838.CK  = CK;
  assign \DFF_839.CK  = CK;
  assign \DFF_84.CK  = CK;
  assign \DFF_840.CK  = CK;
  assign \DFF_841.CK  = CK;
  assign \DFF_842.CK  = CK;
  assign \DFF_842.D  = \DFF_824.Q ;
  assign \DFF_843.CK  = CK;
  assign \DFF_844.CK  = CK;
  assign \DFF_845.CK  = CK;
  assign \DFF_846.CK  = CK;
  assign \DFF_847.CK  = CK;
  assign \DFF_848.CK  = CK;
  assign \DFF_848.D  = \DFF_1087.Q ;
  assign \DFF_849.CK  = CK;
  assign \DFF_85.CK  = CK;
  assign \DFF_850.CK  = CK;
  assign \DFF_851.CK  = CK;
  assign \DFF_852.CK  = CK;
  assign \DFF_853.CK  = CK;
  assign \DFF_854.CK  = CK;
  assign \DFF_855.CK  = CK;
  assign \DFF_856.CK  = CK;
  assign \DFF_856.D  = \DFF_1155.Q ;
  assign \DFF_857.CK  = CK;
  assign \DFF_858.CK  = CK;
  assign \DFF_859.CK  = CK;
  assign \DFF_86.CK  = CK;
  assign \DFF_860.CK  = CK;
  assign \DFF_861.CK  = CK;
  assign \DFF_862.CK  = CK;
  assign \DFF_863.CK  = CK;
  assign \DFF_864.CK  = CK;
  assign \DFF_865.CK  = CK;
  assign \DFF_866.CK  = CK;
  assign \DFF_867.CK  = CK;
  assign \DFF_868.CK  = CK;
  assign \DFF_869.CK  = CK;
  assign \DFF_87.CK  = CK;
  assign \DFF_870.CK  = CK;
  assign \DFF_871.CK  = CK;
  assign \DFF_872.CK  = CK;
  assign \DFF_873.CK  = CK;
  assign \DFF_873.D  = \DFF_34.Q ;
  assign \DFF_874.CK  = CK;
  assign \DFF_875.CK  = CK;
  assign \DFF_876.CK  = CK;
  assign \DFF_877.CK  = CK;
  assign \DFF_878.CK  = CK;
  assign \DFF_879.CK  = CK;
  assign \DFF_88.CK  = CK;
  assign \DFF_880.CK  = CK;
  assign \DFF_881.CK  = CK;
  assign \DFF_882.CK  = CK;
  assign \DFF_883.CK  = CK;
  assign \DFF_884.CK  = CK;
  assign \DFF_885.CK  = CK;
  assign \DFF_885.D  = \DFF_992.Q ;
  assign \DFF_886.CK  = CK;
  assign \DFF_887.CK  = CK;
  assign \DFF_888.CK  = CK;
  assign \DFF_889.CK  = CK;
  assign \DFF_89.CK  = CK;
  assign \DFF_890.CK  = CK;
  assign \DFF_891.CK  = CK;
  assign \DFF_892.CK  = CK;
  assign \DFF_893.CK  = CK;
  assign \DFF_894.CK  = CK;
  assign \DFF_895.CK  = CK;
  assign \DFF_896.CK  = CK;
  assign \DFF_897.CK  = CK;
  assign \DFF_898.CK  = CK;
  assign \DFF_898.D  = \DFF_905.Q ;
  assign \DFF_899.CK  = CK;
  assign \DFF_9.CK  = CK;
  assign \DFF_90.CK  = CK;
  assign \DFF_900.CK  = CK;
  assign \DFF_901.CK  = CK;
  assign \DFF_902.CK  = CK;
  assign \DFF_903.CK  = CK;
  assign \DFF_904.CK  = CK;
  assign \DFF_905.CK  = CK;
  assign \DFF_905.D  = \DFF_970.Q ;
  assign \DFF_906.CK  = CK;
  assign \DFF_906.D  = \DFF_927.Q ;
  assign \DFF_907.CK  = CK;
  assign \DFF_908.CK  = CK;
  assign \DFF_909.CK  = CK;
  assign \DFF_909.D  = \DFF_480.Q ;
  assign \DFF_91.CK  = CK;
  assign \DFF_910.CK  = CK;
  assign \DFF_911.CK  = CK;
  assign \DFF_912.CK  = CK;
  assign \DFF_913.CK  = CK;
  assign \DFF_914.CK  = CK;
  assign \DFF_915.CK  = CK;
  assign \DFF_916.CK  = CK;
  assign \DFF_917.CK  = CK;
  assign \DFF_918.CK  = CK;
  assign \DFF_919.CK  = CK;
  assign \DFF_92.CK  = CK;
  assign \DFF_920.CK  = CK;
  assign \DFF_921.CK  = CK;
  assign \DFF_922.CK  = CK;
  assign \DFF_923.CK  = CK;
  assign \DFF_924.CK  = CK;
  assign \DFF_925.CK  = CK;
  assign \DFF_926.CK  = CK;
  assign \DFF_927.CK  = CK;
  assign \DFF_927.D  = \DFF_655.Q ;
  assign \DFF_928.CK  = CK;
  assign \DFF_929.CK  = CK;
  assign \DFF_93.CK  = CK;
  assign \DFF_930.CK  = CK;
  assign \DFF_931.CK  = CK;
  assign \DFF_932.CK  = CK;
  assign \DFF_933.CK  = CK;
  assign \DFF_934.CK  = CK;
  assign \DFF_935.CK  = CK;
  assign \DFF_936.CK  = CK;
  assign \DFF_937.CK  = CK;
  assign \DFF_938.CK  = CK;
  assign \DFF_939.CK  = CK;
  assign \DFF_94.CK  = CK;
  assign \DFF_940.CK  = CK;
  assign \DFF_941.CK  = CK;
  assign \DFF_942.CK  = CK;
  assign \DFF_942.D  = \DFF_468.Q ;
  assign \DFF_943.CK  = CK;
  assign \DFF_944.CK  = CK;
  assign \DFF_944.D  = \DFF_418.Q ;
  assign \DFF_945.CK  = CK;
  assign \DFF_946.CK  = CK;
  assign \DFF_947.CK  = CK;
  assign \DFF_948.CK  = CK;
  assign \DFF_949.CK  = CK;
  assign \DFF_95.CK  = CK;
  assign \DFF_950.CK  = CK;
  assign \DFF_951.CK  = CK;
  assign \DFF_952.CK  = CK;
  assign \DFF_953.CK  = CK;
  assign \DFF_954.CK  = CK;
  assign \DFF_955.CK  = CK;
  assign \DFF_956.CK  = CK;
  assign \DFF_957.CK  = CK;
  assign \DFF_958.CK  = CK;
  assign \DFF_959.CK  = CK;
  assign \DFF_96.CK  = CK;
  assign \DFF_960.CK  = CK;
  assign \DFF_961.CK  = CK;
  assign \DFF_962.CK  = CK;
  assign \DFF_963.CK  = CK;
  assign \DFF_964.CK  = CK;
  assign \DFF_965.CK  = CK;
  assign \DFF_966.CK  = CK;
  assign \DFF_967.CK  = CK;
  assign \DFF_968.CK  = CK;
  assign \DFF_969.CK  = CK;
  assign \DFF_97.CK  = CK;
  assign \DFF_970.CK  = CK;
  assign \DFF_970.D  = \DFF_1119.Q ;
  assign \DFF_971.CK  = CK;
  assign \DFF_971.D  = \DFF_163.Q ;
  assign \DFF_972.CK  = CK;
  assign \DFF_973.CK  = CK;
  assign \DFF_974.CK  = CK;
  assign \DFF_975.CK  = CK;
  assign \DFF_976.CK  = CK;
  assign \DFF_977.CK  = CK;
  assign \DFF_978.CK  = CK;
  assign \DFF_979.CK  = CK;
  assign \DFF_98.CK  = CK;
  assign \DFF_980.CK  = CK;
  assign \DFF_981.CK  = CK;
  assign \DFF_981.D  = \DFF_672.Q ;
  assign \DFF_982.CK  = CK;
  assign \DFF_983.CK  = CK;
  assign \DFF_984.CK  = CK;
  assign \DFF_985.CK  = CK;
  assign \DFF_986.CK  = CK;
  assign \DFF_987.CK  = CK;
  assign \DFF_988.CK  = CK;
  assign \DFF_989.CK  = CK;
  assign \DFF_99.CK  = CK;
  assign \DFF_990.CK  = CK;
  assign \DFF_990.D  = \DFF_327.Q ;
  assign \DFF_991.CK  = CK;
  assign \DFF_991.D  = \DFF_1345.Q ;
  assign \DFF_992.CK  = CK;
  assign \DFF_992.D  = \DFF_485.Q ;
  assign \DFF_993.CK  = CK;
  assign \DFF_994.CK  = CK;
  assign \DFF_995.CK  = CK;
  assign \DFF_995.D  = \DFF_1219.Q ;
  assign \DFF_996.CK  = CK;
  assign \DFF_997.CK  = CK;
  assign \DFF_997.D  = \DFF_178.Q ;
  assign \DFF_998.CK  = CK;
  assign \DFF_999.CK  = CK;
  assign I13708 = g23612;
  assign I13847 = g35;
  assign I13968 = \DFF_411.Q ;
  assign I13979 = \DFF_551.Q ;
  assign I13990 = \DFF_351.Q ;
  assign I13995 = \DFF_1390.Q ;
  assign I14033 = \DFF_1389.Q ;
  assign I14046 = \DFF_619.Q ;
  assign I14050 = \DFF_1222.Q ;
  assign I14054 = \DFF_761.Q ;
  assign I14079 = g5;
  assign I14119 = \DFF_434.Q ;
  assign I14222 = g53;
  assign I14241 = g54;
  assign I14267 = \DFF_1204.Q ;
  assign I14271 = g56;
  assign I14301 = g57;
  assign I14326 = \DFF_994.Q ;
  assign I14381 = \DFF_828.Q ;
  assign I14409 = \DFF_481.Q ;
  assign I14455 = \DFF_512.Q ;
  assign I14475 = \DFF_790.Q ;
  assign I14505 = \DFF_1229.Q ;
  assign I14537 = \DFF_355.Q ;
  assign I14550 = \DFF_547.Q ;
  assign I14567 = \DFF_1080.Q ;
  assign I14584 = \DFF_1020.Q ;
  assign I14593 = \DFF_428.Q ;
  assign I14679 = g64;
  assign I14742 = g90;
  assign I14773 = g91;
  assign I14797 = g72;
  assign I14823 = \DFF_343.Q ;
  assign I14827 = g73;
  assign I14836 = g113;
  assign I14839 = g124;
  assign I14862 = \DFF_395.Q ;
  assign I14866 = g114;
  assign I14893 = g92;
  assign I14896 = g99;
  assign I14902 = g115;
  assign I14905 = g125;
  assign I14932 = g84;
  assign I14935 = g100;
  assign I14967 = g126;
  assign I14970 = g127;
  assign I14999 = g116;
  assign I15030 = g134;
  assign I15033 = g23612;
  assign I15070 = g120;
  assign I15073 = g135;
  assign I15162 = g44;
  assign I15205 = \DFF_489.Q ;
  assign I15223 = \DFF_448.Q ;
  assign I15250 = \DFF_576.Q ;
  assign I15382 = \DFF_865.Q ;
  assign I15448 = g5;
  assign I15474 = g36;
  assign I15533 = g64;
  assign I15550 = g35;
  assign I15556 = g90;
  assign I15564 = g91;
  assign I15569 = g72;
  assign I15577 = g35;
  assign I15587 = g73;
  assign I15590 = g113;
  assign I15593 = g124;
  assign I15600 = g35;
  assign I15609 = g114;
  assign I15617 = g92;
  assign I15620 = g99;
  assign I15623 = g115;
  assign I15626 = g125;
  assign I15633 = g84;
  assign I15636 = g100;
  assign I15647 = g126;
  assign I15650 = g127;
  assign I15667 = g116;
  assign I15682 = g134;
  assign I15702 = g120;
  assign I15705 = g135;
  assign I15727 = \DFF_434.Q ;
  assign I15736 = g44;
  assign I15773 = g35;
  assign I15782 = g35;
  assign I15788 = g35;
  assign I15811 = \DFF_514.Q ;
  assign I15814 = \DFF_206.Q ;
  assign I15821 = \DFF_477.Q ;
  assign I15831 = g23190;
  assign I15834 = \DFF_829.Q ;
  assign I15843 = \DFF_150.Q ;
  assign I15846 = \DFF_621.Q ;
  assign I15862 = \DFF_1322.Q ;
  assign I15869 = \DFF_1012.Q ;
  assign I15878 = \DFF_420.Q ;
  assign I15893 = g35;
  assign I15906 = g35;
  assign I15915 = g35;
  assign I15918 = \DFF_448.Q ;
  assign I15921 = \DFF_448.Q ;
  assign I15929 = g35;
  assign I15932 = \DFF_448.Q ;
  assign I15942 = \DFF_448.Q ;
  assign I15954 = \DFF_448.Q ;
  assign I15981 = \DFF_994.Q ;
  assign I15987 = \DFF_448.Q ;
  assign I16028 = \DFF_448.Q ;
  assign I16040 = g35;
  assign I16057 = g35;
  assign I16077 = g35;
  assign I16090 = g35;
  assign I16102 = g35;
  assign I16117 = g35;
  assign I16120 = \DFF_961.Q ;
  assign I16135 = g35;
  assign I16150 = g35;
  assign I16163 = \DFF_1181.Q ;
  assign I16289 = \DFF_379.Q ;
  assign I16438 = g53;
  assign I16452 = g54;
  assign I16460 = g35;
  assign I16468 = \DFF_796.Q ;
  assign I16471 = \DFF_489.Q ;
  assign I16476 = g35;
  assign I16479 = g35;
  assign I16486 = g56;
  assign I16489 = \DFF_1424.Q ;
  assign I16492 = \DFF_576.Q ;
  assign I16498 = g35;
  assign I16502 = g35;
  assign I16512 = \DFF_1111.Q ;
  assign I16521 = g35;
  assign I16526 = g35;
  assign I16535 = g57;
  assign I16538 = \DFF_743.Q ;
  assign I16555 = g35;
  assign I16564 = \DFF_417.Q ;
  assign I16579 = \DFF_434.Q ;
  assign I16593 = \DFF_1220.Q ;
  assign I16596 = \DFF_865.Q ;
  assign I16610 = \DFF_434.Q ;
  assign I16613 = g35;
  assign I16651 = \DFF_304.Q ;
  assign I16660 = \DFF_434.Q ;
  assign I16663 = \DFF_434.Q ;
  assign I16688 = \DFF_434.Q ;
  assign I16709 = g35;
  assign I16775 = g23612;
  assign I17008 = g36;
  assign I17094 = \DFF_1424.Q ;
  assign I17098 = g35;
  assign I17101 = g35;
  assign I17104 = g35;
  assign I17108 = g35;
  assign I17111 = g35;
  assign I17114 = \DFF_1111.Q ;
  assign I17118 = g35;
  assign I17121 = g35;
  assign I17125 = g35;
  assign I17128 = g35;
  assign I17131 = \DFF_743.Q ;
  assign I17136 = g35;
  assign I17140 = g35;
  assign I17143 = \DFF_417.Q ;
  assign I17148 = \DFF_1220.Q ;
  assign I17154 = g35;
  assign I17159 = g35;
  assign I17166 = \DFF_304.Q ;
  assign I17173 = g35;
  assign I17181 = g35;
  assign I17188 = g35;
  assign I17198 = g35;
  assign I17207 = g35;
  assign I17228 = g35;
  assign I17249 = g35;
  assign I17276 = g35;
  assign I17355 = g35;
  assign I17374 = g35;
  assign I17392 = g35;
  assign I17401 = g35;
  assign I17420 = g35;
  assign I17425 = g35;
  assign I17436 = g35;
  assign I17442 = g35;
  assign I17456 = g35;
  assign I17471 = g35;
  assign I17488 = g35;
  assign I17491 = g35;
  assign I17507 = g35;
  assign I17590 = g35;
  assign I17609 = \DFF_994.Q ;
  assign I17612 = \DFF_514.Q ;
  assign I17615 = \DFF_206.Q ;
  assign I17633 = \DFF_477.Q ;
  assign I17636 = g53;
  assign I17639 = g35;
  assign I17650 = \DFF_829.Q ;
  assign I17653 = g54;
  assign I17658 = g35;
  assign I17661 = g35;
  assign I17668 = \DFF_150.Q ;
  assign I17671 = \DFF_621.Q ;
  assign I17675 = g35;
  assign I17679 = g35;
  assign I17695 = g56;
  assign I17699 = g35;
  assign I17704 = g35;
  assign I17723 = g35;
  assign I17747 = \DFF_1322.Q ;
  assign I17750 = g57;
  assign I17763 = g35;
  assign I17780 = \DFF_1012.Q ;
  assign I17808 = \DFF_420.Q ;
  assign I17976 = g35;
  assign I18003 = g35;
  assign I18006 = g35;
  assign I18009 = g35;
  assign I18028 = g35;
  assign I18031 = g35;
  assign I18034 = g35;
  assign I18048 = g35;
  assign I18051 = g35;
  assign I18071 = g35;
  assign I18078 = g35;
  assign I18083 = g35;
  assign I18089 = g35;
  assign I18101 = g35;
  assign I18104 = g35;
  assign I18120 = g35;
  assign I18125 = g35;
  assign I18131 = g35;
  assign I18135 = g35;
  assign I18143 = g35;
  assign I18151 = g35;
  assign I18154 = g35;
  assign I18165 = g35;
  assign I18168 = g35;
  assign I18177 = g35;
  assign I18180 = g35;
  assign I18214 = g64;
  assign I18221 = g35;
  assign I18224 = \DFF_961.Q ;
  assign I18238 = g35;
  assign I18245 = g23612;
  assign I18248 = g90;
  assign I18252 = g35;
  assign I18259 = g91;
  assign I18262 = \DFF_1181.Q ;
  assign I18265 = g35;
  assign I18270 = g35;
  assign I18280 = g72;
  assign I18285 = g35;
  assign I18301 = g73;
  assign I18307 = g113;
  assign I18310 = g124;
  assign I18313 = g35;
  assign I18320 = g35;
  assign I18323 = g35;
  assign I18341 = \DFF_489.Q ;
  assign I18344 = g114;
  assign I18350 = g35;
  assign I18364 = g92;
  assign I18367 = g99;
  assign I18373 = g115;
  assign I18376 = \DFF_576.Q ;
  assign I18379 = g125;
  assign I18382 = g35;
  assign I18398 = g35;
  assign I18408 = g84;
  assign I18411 = g100;
  assign I18434 = g35;
  assign I18443 = g126;
  assign I18446 = g127;
  assign I18469 = g35;
  assign I18476 = \DFF_379.Q ;
  assign I18479 = g116;
  assign I18482 = g35;
  assign I18518 = g35;
  assign I18523 = \DFF_865.Q ;
  assign I18526 = g134;
  assign I18571 = g120;
  assign I18574 = g135;
  assign I18674 = g44;
  assign I18810 = g35;
  assign I18822 = g35;
  assign I18829 = g35;
  assign I18832 = g35;
  assign I18839 = g35;
  assign I18842 = g35;
  assign I18849 = g35;
  assign I18852 = g35;
  assign I18855 = g35;
  assign I18858 = g35;
  assign I18861 = \DFF_796.Q ;
  assign I18865 = g35;
  assign I18868 = g35;
  assign I18872 = g35;
  assign I18875 = g35;
  assign I18879 = g23190;
  assign I19384 = g36;
  assign I19661 = g35;
  assign I19707 = \DFF_865.Q ;
  assign I19719 = \DFF_576.Q ;
  assign I19756 = g35;
  assign I19772 = g35;
  assign I19786 = g35;
  assign I19796 = g35;
  assign I19813 = g35;
  assign I19927 = \DFF_489.Q ;
  assign I20216 = g35;
  assign I20529 = g35;
  assign I20542 = g35;
  assign I20562 = g35;
  assign I20584 = g35;
  assign I20690 = g35;
  assign I20846 = g35;
  assign I20895 = g35;
  assign I20913 = g35;
  assign I20937 = g35;
  assign I21006 = g35;
  assign I21033 = g23612;
  assign I21036 = g23612;
  assign I21067 = g35;
  assign I21100 = \DFF_994.Q ;
  assign I21115 = g35;
  assign I21181 = g35;
  assign I21189 = g35;
  assign I21199 = g35;
  assign I21210 = g35;
  assign I21222 = g23190;
  assign I21810 = g35;
  assign I21922 = g35;
  assign I21934 = g35;
  assign I22031 = g35;
  assign I22177 = \DFF_994.Q ;
  assign I22180 = \DFF_994.Q ;
  assign I22745 = \DFF_489.Q ;
  assign I22748 = \DFF_489.Q ;
  assign I22785 = \DFF_576.Q ;
  assign I22788 = \DFF_576.Q ;
  assign I22886 = \DFF_865.Q ;
  assign I22889 = \DFF_865.Q ;
  assign I24920 = g23612;
  assign I26195 = \DFF_994.Q ;
  assign I26479 = g23612;
  assign I26503 = \DFF_489.Q ;
  assign I26508 = \DFF_576.Q ;
  assign I26516 = \DFF_865.Q ;
  assign I26705 = g23612;
  assign I26880 = \DFF_994.Q ;
  assign I26925 = g32185;
  assign I27232 = \DFF_489.Q ;
  assign I27253 = \DFF_576.Q ;
  assign I27314 = \DFF_865.Q ;
  assign I27579 = g23612;
  assign I27730 = \DFF_489.Q ;
  assign I27735 = \DFF_576.Q ;
  assign I27749 = \DFF_865.Q ;
  assign I28349 = \DFF_994.Q ;
  assign I28576 = g32185;
  assign I28582 = \DFF_994.Q ;
  assign I28588 = \DFF_489.Q ;
  assign I28591 = \DFF_576.Q ;
  assign I28594 = \DFF_865.Q ;
  assign I29371 = g32185;
  assign g1 = \DFF_1411.Q ;
  assign g10003 = \DFF_1005.Q ;
  assign g1002 = \DFF_788.Q ;
  assign g10029 = \DFF_1301.Q ;
  assign g10031 = \DFF_1033.Q ;
  assign g10061 = \DFF_198.Q ;
  assign g1008 = \DFF_979.Q ;
  assign g10087 = \DFF_1272.Q ;
  assign g101 = \DFF_417.Q ;
  assign g10107 = \DFF_654.Q ;
  assign g10122 = \DFF_739.Q ;
  assign g10139 = g23612;
  assign g10141 = \DFF_1044.Q ;
  assign g10142 = \DFF_357.Q ;
  assign g1018 = \DFF_421.Q ;
  assign g10198 = \DFF_1059.Q ;
  assign g102 = \DFF_357.Q ;
  assign g10216 = \DFF_132.Q ;
  assign g10230 = \DFF_125.Q ;
  assign g10233 = \DFF_724.Q ;
  assign g1024 = \DFF_70.Q ;
  assign g10272 = \DFF_796.Q ;
  assign g10273 = \DFF_489.Q ;
  assign g10287 = \DFF_1424.Q ;
  assign g10288 = \DFF_736.Q ;
  assign g10295 = \DFF_54.Q ;
  assign g1030 = \DFF_368.Q ;
  assign g10306 = \DFF_1265.Q ;
  assign g10318 = g23190;
  assign g10319 = \DFF_1111.Q ;
  assign g10323 = \DFF_245.Q ;
  assign g10347 = \DFF_1411.Q ;
  assign g10348 = \DFF_1411.Q ;
  assign g10349 = \DFF_919.Q ;
  assign g10350 = \DFF_96.Q ;
  assign g10351 = \DFF_629.Q ;
  assign g10352 = \DFF_47.Q ;
  assign g10353 = \DFF_143.Q ;
  assign g10354 = \DFF_1019.Q ;
  assign g10355 = \DFF_758.Q ;
  assign g10356 = \DFF_1144.Q ;
  assign g10357 = \DFF_698.Q ;
  assign g10358 = \DFF_754.Q ;
  assign g10359 = \DFF_211.Q ;
  assign g1036 = \DFF_131.Q ;
  assign g10360 = \DFF_990.Q ;
  assign g10361 = \DFF_445.Q ;
  assign g10362 = \DFF_1319.Q ;
  assign g10363 = \DFF_650.Q ;
  assign g10366 = \DFF_443.Q ;
  assign g10367 = \DFF_1076.Q ;
  assign g10368 = \DFF_697.Q ;
  assign g10369 = \DFF_196.Q ;
  assign g10370 = \DFF_498.Q ;
  assign g10371 = \DFF_536.Q ;
  assign g10372 = \DFF_180.Q ;
  assign g10373 = \DFF_535.Q ;
  assign g10374 = \DFF_657.Q ;
  assign g10375 = \DFF_517.Q ;
  assign g10376 = \DFF_540.Q ;
  assign g10377 = \DFF_857.Q ;
  assign g10378 = \DFF_144.Q ;
  assign g10379 = \DFF_767.Q ;
  assign g10380 = \DFF_1411.Q ;
  assign g10381 = \DFF_349.Q ;
  assign g10382 = \DFF_26.Q ;
  assign g10383 = \DFF_807.Q ;
  assign g10384 = \DFF_549.Q ;
  assign g10385 = \DFF_615.Q ;
  assign g10386 = \DFF_607.Q ;
  assign g10387 = \DFF_922.Q ;
  assign g10388 = \DFF_1311.Q ;
  assign g10389 = \DFF_609.Q ;
  assign g10390 = \DFF_207.Q ;
  assign g10391 = \DFF_1006.Q ;
  assign g10392 = \DFF_350.Q ;
  assign g10393 = \DFF_313.Q ;
  assign g10394 = \DFF_78.Q ;
  assign g10395 = \DFF_684.Q ;
  assign g10396 = \DFF_439.Q ;
  assign g10397 = \DFF_449.Q ;
  assign g10398 = \DFF_1078.Q ;
  assign g10399 = \DFF_132.Q ;
  assign g10400 = \DFF_190.Q ;
  assign g10401 = \DFF_1283.Q ;
  assign g10402 = \DFF_556.Q ;
  assign g10403 = \DFF_1205.Q ;
  assign g10404 = \DFF_80.Q ;
  assign g10405 = \DFF_429.Q ;
  assign g10406 = \DFF_459.Q ;
  assign g10407 = \DFF_249.Q ;
  assign g10408 = \DFF_75.Q ;
  assign g10409 = \DFF_118.Q ;
  assign g1041 = \DFF_486.Q ;
  assign g10410 = \DFF_138.Q ;
  assign g10411 = \DFF_493.Q ;
  assign g10412 = \DFF_64.Q ;
  assign g10413 = \DFF_878.Q ;
  assign g10414 = \DFF_266.Q ;
  assign g10415 = \DFF_714.Q ;
  assign g10420 = \DFF_244.Q ;
  assign g10427 = \DFF_1005.Q ;
  assign g10428 = \DFF_1068.Q ;
  assign g1046 = \DFF_1144.Q ;
  assign g10473 = \DFF_141.Q ;
  assign g10489 = \DFF_1098.Q ;
  assign g10490 = \DFF_734.Q ;
  assign g10497 = \DFF_198.Q ;
  assign g10499 = \DFF_934.Q ;
  assign g10500 = \DFF_185.Q ;
  assign g10518 = \DFF_289.Q ;
  assign g10519 = \DFF_925.Q ;
  assign g1052 = \DFF_261.Q ;
  assign g10527 = \DFF_1072.Q ;
  assign g10540 = \DFF_393.Q ;
  assign g10541 = \DFF_410.Q ;
  assign g1056 = \DFF_1207.Q ;
  assign g10564 = \DFF_104.Q ;
  assign g10581 = \DFF_1273.Q ;
  assign g10582 = \DFF_748.Q ;
  assign g10588 = g25114;
  assign g106 = \DFF_1059.Q ;
  assign g1061 = \DFF_1133.Q ;
  assign g10615 = g25259;
  assign g10664 = \DFF_853.Q ;
  assign g1070 = \DFF_277.Q ;
  assign g1075 = \DFF_711.Q ;
  assign g1079 = \DFF_643.Q ;
  assign g10795 = \DFF_331.Q ;
  assign g10823 = g26801;
  assign g1083 = \DFF_1122.Q ;
  assign g1087 = \DFF_295.Q ;
  assign g10877 = g12833;
  assign g1094 = \DFF_1382.Q ;
  assign g10960 = \DFF_1122.Q ;
  assign g10980 = \DFF_1110.Q ;
  assign g1099 = \DFF_98.Q ;
  assign g110 = \DFF_379.Q ;
  assign g11011 = \DFF_24.Q ;
  assign g11017 = \DFF_1092.Q ;
  assign g1105 = \DFF_296.Q ;
  assign g111 = \DFF_1220.Q ;
  assign g1111 = \DFF_1290.Q ;
  assign g11136 = \DFF_724.Q ;
  assign g1116 = \DFF_600.Q ;
  assign g112 = \DFF_1181.Q ;
  assign g11237 = \DFF_1425.Q ;
  assign g1124 = \DFF_921.Q ;
  assign g1129 = \DFF_1046.Q ;
  assign g11290 = g23002;
  assign g11317 = \DFF_724.Q ;
  assign g11349 = \DFF_819.Q ;
  assign g1135 = \DFF_137.Q ;
  assign g11388 = \DFF_1420.Q ;
  assign g1141 = \DFF_1274.Q ;
  assign g11418 = \DFF_1001.Q ;
  assign g11447 = \DFF_1234.Q ;
  assign g1146 = \DFF_580.Q ;
  assign g1152 = \DFF_1094.Q ;
  assign g1157 = \DFF_675.Q ;
  assign g11678 = \DFF_1081.Q ;
  assign g117 = \DFF_125.Q ;
  assign g11705 = \DFF_1379.Q ;
  assign g11706 = \DFF_853.Q ;
  assign g1171 = \DFF_214.Q ;
  assign g11714 = \DFF_271.Q ;
  assign g11720 = \DFF_1084.Q ;
  assign g11721 = \DFF_135.Q ;
  assign g11735 = \DFF_538.Q ;
  assign g11736 = \DFF_199.Q ;
  assign g11741 = \DFF_656.Q ;
  assign g11744 = \DFF_746.Q ;
  assign g11753 = \DFF_664.Q ;
  assign g11754 = \DFF_587.Q ;
  assign g11762 = \DFF_35.Q ;
  assign g11769 = \DFF_5.Q ;
  assign g11770 = \DFF_389.Q ;
  assign g11772 = \DFF_853.Q ;
  assign g1178 = \DFF_133.Q ;
  assign g11790 = \DFF_962.Q ;
  assign g11793 = \DFF_746.Q ;
  assign g11796 = \DFF_120.Q ;
  assign g11820 = \DFF_962.Q ;
  assign g11823 = \DFF_962.Q ;
  assign g11826 = \DFF_746.Q ;
  assign g11829 = \DFF_845.Q ;
  assign g1183 = \DFF_563.Q ;
  assign g11832 = \DFF_54.Q ;
  assign g11833 = \DFF_784.Q ;
  assign g11842 = \DFF_934.Q ;
  assign g11845 = \DFF_1078.Q ;
  assign g11852 = \DFF_893.Q ;
  assign g11855 = \DFF_962.Q ;
  assign g11861 = \DFF_245.Q ;
  assign g11872 = \DFF_962.Q ;
  assign g11875 = \DFF_893.Q ;
  assign g11878 = \DFF_746.Q ;
  assign g11884 = \DFF_473.Q ;
  assign g1189 = \DFF_208.Q ;
  assign g11894 = \DFF_962.Q ;
  assign g11897 = \DFF_962.Q ;
  assign g11900 = \DFF_845.Q ;
  assign g11917 = \DFF_893.Q ;
  assign g11920 = \DFF_962.Q ;
  assign g11929 = \DFF_1301.Q ;
  assign g1193 = \DFF_1237.Q ;
  assign g11931 = \DFF_1033.Q ;
  assign g11941 = \DFF_893.Q ;
  assign g11966 = \DFF_654.Q ;
  assign g11986 = \DFF_1044.Q ;
  assign g11987 = \DFF_357.Q ;
  assign g1199 = \DFF_936.Q ;
  assign g12039 = \DFF_1059.Q ;
  assign g1205 = \DFF_90.Q ;
  assign g12077 = \DFF_132.Q ;
  assign g121 = \DFF_1033.Q ;
  assign g12108 = \DFF_125.Q ;
  assign g1211 = \DFF_1103.Q ;
  assign g1216 = \DFF_363.Q ;
  assign g12183 = \DFF_489.Q ;
  assign g12184 = \DFF_515.Q ;
  assign g1221 = \DFF_1057.Q ;
  assign g12238 = \DFF_165.Q ;
  assign g1227 = \DFF_339.Q ;
  assign g12300 = \DFF_46.Q ;
  assign g1233 = \DFF_185.Q ;
  assign g12350 = \DFF_30.Q ;
  assign g1236 = \DFF_791.Q ;
  assign g12367 = g23612;
  assign g12368 = \DFF_752.Q ;
  assign g1239 = \DFF_1308.Q ;
  assign g12399 = \DFF_1084.Q ;
  assign g1242 = \DFF_828.Q ;
  assign g12422 = \DFF_554.Q ;
  assign g12430 = g23652;
  assign g12440 = \DFF_115.Q ;
  assign g1246 = \DFF_343.Q ;
  assign g12470 = \DFF_1158.Q ;
  assign g12477 = \DFF_828.Q ;
  assign g1249 = \DFF_871.Q ;
  assign g12490 = \DFF_1272.Q ;
  assign g1252 = \DFF_901.Q ;
  assign g1256 = \DFF_431.Q ;
  assign g1259 = \DFF_954.Q ;
  assign g1263 = \DFF_454.Q ;
  assign g12640 = g23759;
  assign g1266 = \DFF_1017.Q ;
  assign g1270 = \DFF_913.Q ;
  assign g12729 = g25167;
  assign g12738 = \DFF_598.Q ;
  assign g1274 = \DFF_1109.Q ;
  assign g1277 = \DFF_754.Q ;
  assign g12778 = \DFF_141.Q ;
  assign g12779 = \DFF_575.Q ;
  assign g128 = \DFF_132.Q ;
  assign g1280 = \DFF_1117.Q ;
  assign g12804 = \DFF_599.Q ;
  assign g12805 = \DFF_519.Q ;
  assign g12823 = \DFF_407.Q ;
  assign g1283 = \DFF_323.Q ;
  assign g12830 = \DFF_1320.Q ;
  assign g12831 = \DFF_916.Q ;
  assign g1287 = \DFF_932.Q ;
  assign g12875 = \DFF_615.Q ;
  assign g1291 = \DFF_948.Q ;
  assign g12919 = \DFF_339.Q ;
  assign g12923 = \DFF_1275.Q ;
  assign g12952 = \DFF_934.Q ;
  assign g1296 = \DFF_195.Q ;
  assign g1300 = \DFF_1323.Q ;
  assign g13036 = \DFF_434.Q ;
  assign g13037 = \DFF_434.Q ;
  assign g13039 = \DFF_616.Q ;
  assign g13049 = \DFF_1352.Q ;
  assign g13051 = g6748;
  assign g1306 = \DFF_1131.Q ;
  assign g13061 = \DFF_434.Q ;
  assign g13062 = \DFF_434.Q ;
  assign g13068 = \DFF_1087.Q ;
  assign g13070 = g6749;
  assign g13082 = \DFF_434.Q ;
  assign g13085 = \DFF_1119.Q ;
  assign g13087 = g6750;
  assign g13099 = \DFF_163.Q ;
  assign g13106 = \DFF_434.Q ;
  assign g1311 = \DFF_1292.Q ;
  assign g13117 = \DFF_434.Q ;
  assign g1312 = \DFF_1039.Q ;
  assign g13138 = g26801;
  assign g13174 = \DFF_339.Q ;
  assign g13189 = \DFF_1275.Q ;
  assign g1319 = \DFF_1092.Q ;
  assign g1322 = \DFF_990.Q ;
  assign g13259 = \DFF_600.Q ;
  assign g13272 = \DFF_327.Q ;
  assign g13302 = g6751;
  assign g1333 = \DFF_408.Q ;
  assign g1339 = \DFF_67.Q ;
  assign g13412 = g6752;
  assign g1345 = \DFF_1153.Q ;
  assign g13484 = \DFF_434.Q ;
  assign g13494 = g6753;
  assign g13505 = \DFF_434.Q ;
  assign g1351 = \DFF_1343.Q ;
  assign g13510 = g23002;
  assign g13522 = \DFF_434.Q ;
  assign g136 = \DFF_489.Q ;
  assign g1361 = \DFF_577.Q ;
  assign g1367 = \DFF_1227.Q ;
  assign g1373 = \DFF_316.Q ;
  assign g1379 = \DFF_1419.Q ;
  assign g1384 = \DFF_66.Q ;
  assign g13856 = \DFF_1425.Q ;
  assign g13865 = \DFF_76.Q ;
  assign g13881 = \DFF_369.Q ;
  assign g1389 = \DFF_211.Q ;
  assign g13895 = \DFF_529.Q ;
  assign g13906 = \DFF_662.Q ;
  assign g13926 = \DFF_468.Q ;
  assign g1395 = \DFF_1008.Q ;
  assign g13966 = \DFF_401.Q ;
  assign g1399 = \DFF_937.Q ;
  assign g1404 = \DFF_740.Q ;
  assign g14096 = \DFF_152.Q ;
  assign g14125 = \DFF_404.Q ;
  assign g1413 = \DFF_614.Q ;
  assign g14147 = \DFF_380.Q ;
  assign g14149 = \DFF_448.Q ;
  assign g14150 = \DFF_448.Q ;
  assign g14167 = \DFF_764.Q ;
  assign g14169 = \DFF_448.Q ;
  assign g14173 = g6744;
  assign g1418 = \DFF_422.Q ;
  assign g14183 = \DFF_448.Q ;
  assign g14184 = \DFF_448.Q ;
  assign g14189 = \DFF_585.Q ;
  assign g14191 = \DFF_448.Q ;
  assign g14198 = g6745;
  assign g142 = \DFF_359.Q ;
  assign g14201 = \DFF_561.Q ;
  assign g14203 = \DFF_448.Q ;
  assign g14205 = \DFF_448.Q ;
  assign g14217 = \DFF_1106.Q ;
  assign g14219 = \DFF_448.Q ;
  assign g1422 = \DFF_146.Q ;
  assign g14255 = \DFF_448.Q ;
  assign g1426 = \DFF_1110.Q ;
  assign g14277 = \DFF_1078.Q ;
  assign g1430 = \DFF_372.Q ;
  assign g14308 = g23612;
  assign g14332 = g23652;
  assign g14357 = g6746;
  assign g14359 = \DFF_828.Q ;
  assign g1437 = \DFF_169.Q ;
  assign g14385 = \DFF_1301.Q ;
  assign g14386 = \DFF_1033.Q ;
  assign g1442 = \DFF_182.Q ;
  assign g14421 = \DFF_1155.Q ;
  assign g14441 = \DFF_654.Q ;
  assign g14443 = g23759;
  assign g14451 = \DFF_34.Q ;
  assign g1448 = \DFF_403.Q ;
  assign g14509 = \DFF_1044.Q ;
  assign g14510 = \DFF_357.Q ;
  assign g14518 = \DFF_642.Q ;
  assign g1454 = \DFF_193.Q ;
  assign g14562 = g6747;
  assign g14563 = g25114;
  assign g14564 = \DFF_1059.Q ;
  assign g14582 = \DFF_132.Q ;
  assign g1459 = \DFF_327.Q ;
  assign g14597 = \DFF_537.Q ;
  assign g146 = \DFF_1060.Q ;
  assign g14609 = \DFF_125.Q ;
  assign g14635 = \DFF_1262.Q ;
  assign g14639 = g25167;
  assign g14662 = \DFF_655.Q ;
  assign g1467 = \DFF_424.Q ;
  assign g14673 = \DFF_1102.Q ;
  assign g14676 = \DFF_489.Q ;
  assign g14694 = \DFF_1335.Q ;
  assign g14705 = \DFF_905.Q ;
  assign g1472 = \DFF_595.Q ;
  assign g14738 = \DFF_326.Q ;
  assign g14749 = \DFF_836.Q ;
  assign g14779 = \DFF_188.Q ;
  assign g1478 = \DFF_774.Q ;
  assign g14790 = \DFF_141.Q ;
  assign g14828 = \DFF_806.Q ;
  assign g1484 = \DFF_720.Q ;
  assign g14873 = g25259;
  assign g1489 = \DFF_822.Q ;
  assign g14912 = \DFF_748.Q ;
  assign g1495 = \DFF_167.Q ;
  assign g150 = \DFF_582.Q ;
  assign g1500 = \DFF_60.Q ;
  assign g15078 = \DFF_680.D ;
  assign g15079 = \DFF_391.D ;
  assign g15083 = \DFF_611.D ;
  assign g15084 = \DFF_1101.D ;
  assign g1514 = \DFF_1148.Q ;
  assign g1521 = \DFF_1407.Q ;
  assign g1526 = \DFF_717.Q ;
  assign g153 = \DFF_409.Q ;
  assign g1532 = \DFF_202.Q ;
  assign g1536 = \DFF_1159.Q ;
  assign g1542 = \DFF_1189.Q ;
  assign g1548 = \DFF_1371.Q ;
  assign g1554 = \DFF_1194.Q ;
  assign g1559 = \DFF_1313.Q ;
  assign g1564 = \DFF_375.Q ;
  assign g157 = \DFF_318.Q ;
  assign g1570 = \DFF_1275.Q ;
  assign g1576 = \DFF_1072.Q ;
  assign g1579 = \DFF_171.Q ;
  assign g1582 = \DFF_334.Q ;
  assign g1585 = \DFF_481.Q ;
  assign g1589 = \DFF_395.Q ;
  assign g1592 = \DFF_1054.Q ;
  assign g15932 = \DFF_934.Q ;
  assign g16 = \DFF_355.Q ;
  assign g160 = \DFF_555.Q ;
  assign g1600 = \DFF_32.Q ;
  assign g1604 = \DFF_246.Q ;
  assign g1608 = \DFF_564.Q ;
  assign g1612 = \DFF_1180.Q ;
  assign g1616 = \DFF_735.Q ;
  assign g1620 = \DFF_864.Q ;
  assign g16216 = \DFF_357.Q ;
  assign g16228 = \DFF_1059.Q ;
  assign g1624 = \DFF_1064.Q ;
  assign g16284 = g23002;
  assign g16300 = \DFF_132.Q ;
  assign g1632 = \DFF_164.Q ;
  assign g16320 = g35;
  assign g1636 = \DFF_1127.Q ;
  assign g164 = \DFF_1339.Q ;
  assign g1644 = \DFF_1089.Q ;
  assign g1648 = \DFF_1344.Q ;
  assign g16530 = g35;
  assign g16540 = \DFF_748.Q ;
  assign g1657 = \DFF_794.Q ;
  assign g16579 = g23190;
  assign g16580 = g6753;
  assign g16603 = \DFF_1293.Q ;
  assign g16609 = g35;
  assign g16624 = \DFF_1354.Q ;
  assign g16627 = \DFF_220.Q ;
  assign g16631 = g35;
  assign g16632 = g35;
  assign g1664 = \DFF_342.Q ;
  assign g16643 = g6752;
  assign g16644 = g6748;
  assign g16656 = \DFF_81.Q ;
  assign g16659 = \DFF_181.Q ;
  assign g16661 = g35;
  assign g16676 = g6749;
  assign g16677 = \DFF_1033.Q ;
  assign g1668 = \DFF_646.Q ;
  assign g16686 = \DFF_1359.Q ;
  assign g16693 = \DFF_785.Q ;
  assign g16695 = g35;
  assign g16708 = g6750;
  assign g16709 = \DFF_125.Q ;
  assign g16718 = \DFF_1038.Q ;
  assign g16722 = \DFF_1300.Q ;
  assign g16726 = g35;
  assign g16727 = g35;
  assign g16738 = g6747;
  assign g16744 = \DFF_942.Q ;
  assign g16748 = \DFF_1219.Q ;
  assign g16750 = g35;
  assign g16767 = g6744;
  assign g1677 = \DFF_1069.Q ;
  assign g16775 = \DFF_305.Q ;
  assign g168 = \DFF_533.Q ;
  assign g1682 = \DFF_293.Q ;
  assign g1687 = \DFF_1266.Q ;
  assign g16872 = g6745;
  assign g16873 = g6746;
  assign g16874 = \DFF_856.Q ;
  assign g1691 = \DFF_1281.Q ;
  assign g16920 = \DFF_1425.Q ;
  assign g16924 = \DFF_873.Q ;
  assign g16955 = \DFF_367.Q ;
  assign g16958 = g26801;
  assign g1696 = \DFF_583.Q ;
  assign g16960 = \DFF_1044.Q ;
  assign g16963 = g6751;
  assign g16968 = g26801;
  assign g1700 = \DFF_446.Q ;
  assign g17010 = \DFF_1078.Q ;
  assign g1706 = \DFF_212.Q ;
  assign g17085 = g26801;
  assign g17088 = \DFF_654.Q ;
  assign g1710 = \DFF_1277.Q ;
  assign g1714 = \DFF_33.Q ;
  assign g17141 = \DFF_1301.Q ;
  assign g17155 = g25114;
  assign g17157 = g35;
  assign g17197 = g25167;
  assign g1720 = \DFF_1226.Q ;
  assign g17216 = g35;
  assign g17221 = \DFF_489.Q ;
  assign g1724 = \DFF_1418.Q ;
  assign g17242 = g35;
  assign g1728 = \DFF_272.Q ;
  assign g17291 = \DFF_711.Q ;
  assign g17292 = g27831;
  assign g17301 = g35;
  assign g17316 = \DFF_643.Q ;
  assign g17320 = \DFF_422.Q ;
  assign g17325 = \DFF_141.Q ;
  assign g1736 = \DFF_41.Q ;
  assign g17366 = g35;
  assign g174 = \DFF_292.Q ;
  assign g1740 = \DFF_1258.Q ;
  assign g17400 = \DFF_1122.Q ;
  assign g17404 = \DFF_146.Q ;
  assign g17408 = g23612;
  assign g17410 = g35;
  assign g17411 = g35;
  assign g17423 = \DFF_1110.Q ;
  assign g17429 = g25259;
  assign g17431 = g23652;
  assign g1744 = \DFF_16.Q ;
  assign g17465 = g35;
  assign g17466 = g35;
  assign g17470 = g35;
  assign g17471 = g35;
  assign g1748 = \DFF_306.Q ;
  assign g17487 = \DFF_828.Q ;
  assign g17489 = g35;
  assign g17491 = g35;
  assign g17512 = g35;
  assign g17519 = \DFF_906.Q ;
  assign g1752 = \DFF_173.Q ;
  assign g1756 = \DFF_1137.Q ;
  assign g17577 = \DFF_566.Q ;
  assign g17580 = \DFF_263.Q ;
  assign g17590 = g23759;
  assign g1760 = \DFF_552.Q ;
  assign g17604 = \DFF_101.Q ;
  assign g17607 = \DFF_110.Q ;
  assign g17639 = \DFF_360.Q ;
  assign g17646 = \DFF_737.Q ;
  assign g17649 = \DFF_315.Q ;
  assign g17674 = \DFF_927.Q ;
  assign g17678 = \DFF_783.Q ;
  assign g1768 = \DFF_984.Q ;
  assign g17685 = \DFF_123.Q ;
  assign g17688 = \DFF_1248.Q ;
  assign g17711 = \DFF_117.Q ;
  assign g17715 = \DFF_279.Q ;
  assign g1772 = \DFF_500.Q ;
  assign g17722 = \DFF_1185.Q ;
  assign g17733 = g26801;
  assign g17739 = \DFF_797.Q ;
  assign g17743 = \DFF_898.Q ;
  assign g17760 = \DFF_474.Q ;
  assign g17764 = \DFF_780.Q ;
  assign g17778 = \DFF_1196.Q ;
  assign g17782 = g26801;
  assign g17787 = \DFF_765.Q ;
  assign g1779 = \DFF_567.Q ;
  assign g17794 = g35;
  assign g17813 = \DFF_695.Q ;
  assign g17819 = \DFF_848.Q ;
  assign g1783 = \DFF_1037.Q ;
  assign g17845 = \DFF_970.Q ;
  assign g17871 = \DFF_971.Q ;
  assign g1792 = \DFF_1375.Q ;
  assign g1798 = \DFF_153.Q ;
  assign g1802 = \DFF_18.Q ;
  assign g18088 = g23190;
  assign g18092 = g6753;
  assign g18093 = g6752;
  assign g18094 = g6748;
  assign g18095 = g6749;
  assign g18096 = g6750;
  assign g18097 = g6747;
  assign g18098 = g6744;
  assign g18099 = g6745;
  assign g18100 = g6751;
  assign g18101 = g6746;
  assign g1811 = \DFF_1167.Q ;
  assign g1816 = \DFF_435.Q ;
  assign g182 = \DFF_1045.Q ;
  assign g1821 = \DFF_1114.Q ;
  assign g18215 = \DFF_800.D ;
  assign g18216 = \DFF_999.D ;
  assign g1825 = \DFF_977.Q ;
  assign g18273 = \DFF_1292.D ;
  assign g18274 = \DFF_1353.D ;
  assign g1830 = \DFF_1051.Q ;
  assign g1834 = \DFF_1243.Q ;
  assign g1840 = \DFF_649.Q ;
  assign g18421 = \DFF_680.D ;
  assign g18422 = \DFF_391.D ;
  assign g1844 = \DFF_814.Q ;
  assign g1848 = \DFF_1075.Q ;
  assign g18527 = \DFF_611.D ;
  assign g18528 = \DFF_1101.D ;
  assign g1854 = \DFF_882.Q ;
  assign g1858 = \DFF_1163.Q ;
  assign g18597 = \DFF_1381.D ;
  assign g18598 = g21727;
  assign g1862 = \DFF_111.Q ;
  assign g18695 = \DFF_501.D ;
  assign g18696 = \DFF_200.D ;
  assign g1870 = \DFF_973.Q ;
  assign g18726 = \DFF_1402.D ;
  assign g18727 = \DFF_1165.D ;
  assign g1874 = \DFF_1172.Q ;
  assign g1878 = \DFF_1422.Q ;
  assign g1882 = \DFF_2.Q ;
  assign g18827 = g35;
  assign g18828 = g35;
  assign g18829 = g35;
  assign g18830 = g35;
  assign g18831 = g35;
  assign g18832 = g35;
  assign g1886 = \DFF_968.Q ;
  assign g18874 = g35;
  assign g18875 = g35;
  assign g18876 = g35;
  assign g18877 = g35;
  assign g18878 = g35;
  assign g18880 = g35;
  assign g18881 = \DFF_934.Q ;
  assign g18882 = \DFF_934.Q ;
  assign g18883 = g35;
  assign g18884 = g35;
  assign g18885 = g35;
  assign g18886 = g35;
  assign g18887 = g35;
  assign g18888 = g35;
  assign g18889 = g35;
  assign g18891 = g35;
  assign g18892 = g35;
  assign g18894 = g35;
  assign g18895 = g35;
  assign g18896 = g35;
  assign g18897 = g35;
  assign g18898 = \DFF_417.Q ;
  assign g1890 = \DFF_504.Q ;
  assign g18903 = g35;
  assign g18904 = g35;
  assign g18905 = g35;
  assign g18907 = g35;
  assign g18908 = g35;
  assign g18911 = \DFF_1424.Q ;
  assign g18916 = g35;
  assign g18917 = g35;
  assign g18926 = g23759;
  assign g18929 = g35;
  assign g18931 = g35;
  assign g18932 = g35;
  assign g18938 = g35;
  assign g18939 = g35;
  assign g1894 = \DFF_705.Q ;
  assign g18940 = g23652;
  assign g18944 = g35;
  assign g18945 = g35;
  assign g18946 = g35;
  assign g18947 = g35;
  assign g18952 = g35;
  assign g18953 = g35;
  assign g18954 = g92;
  assign g18975 = g35;
  assign g18976 = g35;
  assign g18977 = g35;
  assign g18978 = g35;
  assign g18979 = g35;
  assign g18980 = g35;
  assign g18983 = g35;
  assign g18984 = g100;
  assign g18988 = g35;
  assign g18989 = g35;
  assign g18990 = g35;
  assign g18991 = g35;
  assign g19 = \DFF_1229.Q ;
  assign g1902 = \DFF_1202.Q ;
  assign g1906 = \DFF_759.Q ;
  assign g19067 = g35;
  assign g19068 = g35;
  assign g191 = \DFF_842.Q ;
  assign g1913 = \DFF_1009.Q ;
  assign g19144 = g35;
  assign g1917 = \DFF_174.Q ;
  assign g19208 = g35;
  assign g1926 = \DFF_103.Q ;
  assign g19273 = g35;
  assign g19276 = g35;
  assign g1932 = \DFF_1063.Q ;
  assign g19330 = g113;
  assign g19334 = \DFF_1207.Q ;
  assign g19343 = g35;
  assign g19345 = g134;
  assign g19351 = g35;
  assign g19352 = g35;
  assign g19357 = \DFF_937.Q ;
  assign g1936 = \DFF_620.Q ;
  assign g19360 = g35;
  assign g19365 = g35;
  assign g19366 = g35;
  assign g19368 = g35;
  assign g19370 = g35;
  assign g19373 = g35;
  assign g19376 = g127;
  assign g19379 = g124;
  assign g19385 = g35;
  assign g19386 = g35;
  assign g19387 = g35;
  assign g19389 = g116;
  assign g19394 = g35;
  assign g19395 = g35;
  assign g19396 = g35;
  assign g19397 = g35;
  assign g19398 = g35;
  assign g19399 = g35;
  assign g194 = \DFF_824.Q ;
  assign g19409 = g35;
  assign g19410 = g35;
  assign g19411 = g35;
  assign g19412 = g35;
  assign g19414 = g35;
  assign g19415 = g35;
  assign g19416 = g35;
  assign g19417 = g64;
  assign g19421 = g35;
  assign g19429 = g35;
  assign g19431 = g35;
  assign g19432 = g35;
  assign g19433 = g35;
  assign g19434 = g35;
  assign g19435 = g35;
  assign g19437 = g35;
  assign g19438 = g35;
  assign g19439 = g35;
  assign g19440 = g35;
  assign g19443 = g35;
  assign g19445 = g35;
  assign g19446 = g23190;
  assign g1945 = \DFF_772.Q ;
  assign g19451 = g35;
  assign g19452 = g35;
  assign g19454 = g35;
  assign g19458 = g23612;
  assign g19468 = g35;
  assign g19469 = g35;
  assign g19470 = g35;
  assign g19471 = g35;
  assign g19472 = g35;
  assign g19473 = g35;
  assign g19476 = g35;
  assign g19477 = g35;
  assign g19478 = g35;
  assign g19479 = g35;
  assign g19480 = g35;
  assign g19481 = g35;
  assign g19482 = g35;
  assign g19489 = g35;
  assign g19490 = g35;
  assign g19491 = g35;
  assign g19492 = g35;
  assign g19493 = g35;
  assign g19494 = g35;
  assign g19498 = g35;
  assign g19499 = g35;
  assign g1950 = \DFF_455.Q ;
  assign g19503 = g35;
  assign g19504 = g35;
  assign g19505 = g35;
  assign g19517 = g35;
  assign g19519 = g35;
  assign g19520 = g35;
  assign g19523 = g35;
  assign g19526 = g35;
  assign g19527 = g35;
  assign g19528 = g35;
  assign g19529 = g35;
  assign g19531 = g35;
  assign g19532 = g35;
  assign g19537 = g35;
  assign g19538 = g35;
  assign g19539 = g35;
  assign g19541 = g35;
  assign g19542 = g35;
  assign g19543 = g35;
  assign g19544 = g35;
  assign g1955 = \DFF_832.Q ;
  assign g19552 = g35;
  assign g19553 = g35;
  assign g19554 = g35;
  assign g19558 = g35;
  assign g19559 = g35;
  assign g19565 = g35;
  assign g19566 = g35;
  assign g19567 = g35;
  assign g19569 = g35;
  assign g19570 = g35;
  assign g19573 = g35;
  assign g19574 = g35;
  assign g19577 = g35;
  assign g19579 = g35;
  assign g19580 = g35;
  assign g19586 = g35;
  assign g1959 = \DFF_777.Q ;
  assign g19600 = g35;
  assign g19602 = g35;
  assign g19603 = g35;
  assign g19606 = g120;
  assign g19612 = g35;
  assign g19617 = g35;
  assign g19618 = g35;
  assign g19620 = g72;
  assign g19626 = g114;
  assign g19629 = g35;
  assign g19630 = g35;
  assign g19633 = g35;
  assign g19634 = g35;
  assign g19635 = g35;
  assign g19636 = g35;
  assign g19638 = g73;
  assign g1964 = \DFF_1216.Q ;
  assign g19644 = \DFF_796.Q ;
  assign g19649 = g35;
  assign g19650 = g35;
  assign g19652 = g35;
  assign g19653 = g35;
  assign g19654 = g35;
  assign g19657 = g35;
  assign g19658 = g35;
  assign g19659 = g35;
  assign g19662 = g125;
  assign g19666 = \DFF_961.Q ;
  assign g19670 = g35;
  assign g19672 = g35;
  assign g19673 = g35;
  assign g19675 = g35;
  assign g19676 = g35;
  assign g19677 = g35;
  assign g19678 = g35;
  assign g19679 = g35;
  assign g1968 = \DFF_42.Q ;
  assign g19682 = g35;
  assign g19683 = g35;
  assign g19685 = g35;
  assign g19686 = g35;
  assign g19687 = g35;
  assign g19688 = g35;
  assign g19689 = g35;
  assign g19690 = g35;
  assign g19694 = \DFF_621.Q ;
  assign g19695 = g35;
  assign g19696 = g35;
  assign g19697 = g35;
  assign g19698 = g35;
  assign g19709 = g35;
  assign g19710 = g35;
  assign g19711 = g35;
  assign g19712 = g35;
  assign g19713 = g35;
  assign g19714 = g35;
  assign g19718 = g35;
  assign g19719 = g35;
  assign g19730 = g35;
  assign g19731 = g35;
  assign g19732 = g35;
  assign g19733 = g35;
  assign g19734 = g35;
  assign g19737 = g35;
  assign g19739 = g35;
  assign g1974 = \DFF_912.Q ;
  assign g19741 = g35;
  assign g19742 = g35;
  assign g19743 = g35;
  assign g19744 = g35;
  assign g19745 = g35;
  assign g19747 = g35;
  assign g19748 = g35;
  assign g19750 = g35;
  assign g19753 = g35;
  assign g19754 = g35;
  assign g19755 = g35;
  assign g19757 = g90;
  assign g19760 = g35;
  assign g19761 = g35;
  assign g19762 = g35;
  assign g19763 = g35;
  assign g19765 = g35;
  assign g19766 = g35;
  assign g19769 = g35;
  assign g19770 = g35;
  assign g19771 = g35;
  assign g19772 = g35;
  assign g19773 = g135;
  assign g19776 = g35;
  assign g19777 = g35;
  assign g19779 = g35;
  assign g1978 = \DFF_1179.Q ;
  assign g19780 = g35;
  assign g19781 = g35;
  assign g19783 = g35;
  assign g19785 = g35;
  assign g19786 = g35;
  assign g19787 = g35;
  assign g19789 = g35;
  assign g19790 = g35;
  assign g19794 = g35;
  assign g19798 = g35;
  assign g19799 = g35;
  assign g19800 = g35;
  assign g1982 = \DFF_1184.Q ;
  assign g19852 = g35;
  assign g19860 = g35;
  assign g19861 = g35;
  assign g19862 = \DFF_828.Q ;
  assign g19865 = g35;
  assign g19872 = g35;
  assign g19878 = g35;
  assign g1988 = \DFF_1369.Q ;
  assign g19881 = g35;
  assign g19885 = g35;
  assign g199 = \DFF_715.Q ;
  assign g19902 = g35;
  assign g19905 = g35;
  assign g19912 = g35;
  assign g19915 = g35;
  assign g1992 = \DFF_520.Q ;
  assign g19930 = g35;
  assign g19931 = g35;
  assign g19947 = g35;
  assign g19950 = g35;
  assign g19952 = g35;
  assign g1996 = \DFF_1413.Q ;
  assign g19960 = g35;
  assign g19961 = g35;
  assign g19963 = g35;
  assign g19964 = g35;
  assign g19979 = g35;
  assign g19980 = g35;
  assign g19996 = g35;
  assign g19998 = g35;
  assign g20004 = g35;
  assign g20005 = g35;
  assign g20006 = g35;
  assign g20008 = g35;
  assign g20009 = g35;
  assign g20010 = g35;
  assign g20025 = g35;
  assign g20026 = g35;
  assign g20028 = \DFF_1111.Q ;
  assign g20036 = g35;
  assign g20037 = g35;
  assign g20038 = g35;
  assign g2004 = \DFF_1394.Q ;
  assign g20040 = g35;
  assign g20041 = \DFF_1220.Q ;
  assign g20049 = \DFF_1425.Q ;
  assign g20050 = \DFF_1425.Q ;
  assign g20052 = g35;
  assign g20053 = g35;
  assign g20054 = g35;
  assign g20057 = g35;
  assign g20058 = g35;
  assign g20059 = g35;
  assign g20064 = g35;
  assign g20066 = g35;
  assign g20067 = g35;
  assign g20071 = g35;
  assign g20072 = g35;
  assign g20079 = g35;
  assign g2008 = \DFF_255.Q ;
  assign g20080 = g35;
  assign g20087 = g35;
  assign g20088 = g35;
  assign g20089 = g35;
  assign g20090 = g35;
  assign g20091 = g35;
  assign g20096 = g35;
  assign g20097 = g44;
  assign g20101 = g35;
  assign g20102 = g35;
  assign g20103 = g35;
  assign g20104 = g35;
  assign g20105 = g35;
  assign g20106 = g35;
  assign g20110 = g35;
  assign g20113 = g35;
  assign g2012 = \DFF_924.Q ;
  assign g20128 = g35;
  assign g20129 = g35;
  assign g20130 = g35;
  assign g20132 = g35;
  assign g20144 = g35;
  assign g20145 = g35;
  assign g20146 = g35;
  assign g20147 = g35;
  assign g20153 = g35;
  assign g20157 = g35;
  assign g20158 = g35;
  assign g20159 = g35;
  assign g2016 = \DFF_465.Q ;
  assign g20164 = g35;
  assign g20166 = g35;
  assign g20167 = g35;
  assign g20168 = g35;
  assign g20178 = g35;
  assign g20179 = g35;
  assign g20180 = g35;
  assign g20182 = g35;
  assign g20190 = g35;
  assign g20191 = g35;
  assign g20194 = g35;
  assign g20195 = g35;
  assign g20197 = g35;
  assign g2020 = \DFF_641.Q ;
  assign g20204 = g57;
  assign g20207 = g35;
  assign g20208 = g35;
  assign g20209 = g35;
  assign g20210 = g35;
  assign g20211 = g35;
  assign g20213 = g35;
  assign g20229 = g35;
  assign g20231 = g35;
  assign g20232 = g35;
  assign g20233 = g35;
  assign g20235 = g35;
  assign g20238 = g35;
  assign g20239 = g35;
  assign g2024 = \DFF_809.Q ;
  assign g20240 = g35;
  assign g20242 = g53;
  assign g20247 = g35;
  assign g20265 = g35;
  assign g20266 = g35;
  assign g20267 = g35;
  assign g20268 = g35;
  assign g20270 = g35;
  assign g20273 = g35;
  assign g20274 = g35;
  assign g20275 = g35;
  assign g20277 = g56;
  assign g2028 = \DFF_1070.Q ;
  assign g203 = \DFF_96.Q ;
  assign g20320 = g35;
  assign g20321 = g35;
  assign g20322 = g35;
  assign g20323 = g35;
  assign g20324 = g35;
  assign g20325 = g35;
  assign g20326 = g35;
  assign g20327 = g35;
  assign g20329 = g35;
  assign g2036 = \DFF_862.Q ;
  assign g20372 = g35;
  assign g20373 = g35;
  assign g20374 = g35;
  assign g20379 = g35;
  assign g20380 = g35;
  assign g20381 = g35;
  assign g20382 = g35;
  assign g20383 = g35;
  assign g20384 = g35;
  assign g20385 = g35;
  assign g20386 = g35;
  assign g20387 = g35;
  assign g20389 = g35;
  assign g2040 = \DFF_671.Q ;
  assign g20432 = g35;
  assign g20433 = g35;
  assign g20434 = g35;
  assign g20435 = g35;
  assign g20441 = g35;
  assign g20442 = g35;
  assign g20443 = g35;
  assign g20444 = g35;
  assign g20445 = g35;
  assign g20446 = g35;
  assign g20447 = g35;
  assign g20448 = g35;
  assign g20449 = g35;
  assign g20450 = g35;
  assign g20451 = g35;
  assign g20452 = g35;
  assign g2047 = \DFF_472.Q ;
  assign g20494 = g35;
  assign g20495 = g35;
  assign g20496 = g35;
  assign g20497 = g35;
  assign g20498 = g35;
  assign g20499 = g35;
  assign g20500 = g35;
  assign g20501 = g35;
  assign g20502 = g35;
  assign g20503 = g35;
  assign g20504 = g35;
  assign g20505 = g35;
  assign g20506 = g35;
  assign g20507 = g35;
  assign g20508 = g35;
  assign g20509 = g35;
  assign g2051 = \DFF_1236.Q ;
  assign g20510 = g35;
  assign g20511 = g35;
  assign g20512 = g35;
  assign g20513 = g35;
  assign g20514 = g35;
  assign g20515 = g35;
  assign g20523 = g35;
  assign g20524 = g35;
  assign g20525 = g35;
  assign g20526 = g35;
  assign g20527 = g35;
  assign g20528 = g35;
  assign g20529 = g35;
  assign g20530 = g35;
  assign g20532 = g35;
  assign g20533 = g35;
  assign g20534 = g35;
  assign g20535 = g35;
  assign g20536 = g35;
  assign g20537 = g35;
  assign g20538 = g35;
  assign g20539 = g35;
  assign g20541 = g35;
  assign g20542 = g35;
  assign g20543 = g35;
  assign g20544 = g35;
  assign g20545 = g35;
  assign g20546 = g35;
  assign g20547 = g35;
  assign g20548 = g35;
  assign g20549 = g35;
  assign g20551 = g35;
  assign g20552 = g35;
  assign g20553 = g35;
  assign g20554 = g35;
  assign g20555 = g35;
  assign g20556 = g35;
  assign g20557 = \DFF_1078.Q ;
  assign g20558 = \DFF_1078.Q ;
  assign g20560 = g35;
  assign g20561 = g35;
  assign g20562 = g35;
  assign g20563 = g35;
  assign g20564 = g35;
  assign g20565 = g35;
  assign g20566 = g35;
  assign g20567 = g35;
  assign g20568 = g35;
  assign g20569 = g35;
  assign g20570 = g35;
  assign g20571 = g35;
  assign g20573 = g35;
  assign g20574 = g35;
  assign g20575 = g35;
  assign g20576 = g35;
  assign g20577 = g35;
  assign g20578 = g35;
  assign g20579 = g35;
  assign g20580 = g35;
  assign g20582 = g35;
  assign g20583 = g35;
  assign g20584 = g35;
  assign g20585 = g35;
  assign g20586 = g35;
  assign g20587 = g35;
  assign g20588 = g35;
  assign g20589 = g35;
  assign g20590 = g35;
  assign g20591 = g35;
  assign g20592 = g35;
  assign g20593 = g35;
  assign g20594 = g35;
  assign g20597 = g35;
  assign g20598 = g35;
  assign g20599 = g35;
  assign g2060 = \DFF_1295.Q ;
  assign g20600 = g35;
  assign g20601 = g35;
  assign g20603 = g35;
  assign g20604 = g35;
  assign g20605 = g35;
  assign g20606 = g35;
  assign g20607 = g35;
  assign g20608 = g35;
  assign g20609 = g35;
  assign g20610 = g35;
  assign g20611 = g35;
  assign g20612 = g35;
  assign g20613 = g35;
  assign g20614 = g35;
  assign g20615 = g35;
  assign g20616 = g35;
  assign g20617 = g35;
  assign g20618 = g35;
  assign g20622 = g35;
  assign g20623 = g35;
  assign g20624 = g35;
  assign g20625 = g35;
  assign g20626 = g35;
  assign g20627 = g35;
  assign g20629 = g35;
  assign g20630 = g35;
  assign g20631 = g35;
  assign g20632 = g35;
  assign g20633 = g35;
  assign g20634 = g35;
  assign g20635 = g35;
  assign g20636 = g35;
  assign g20637 = g35;
  assign g20638 = g35;
  assign g20639 = g35;
  assign g20640 = g35;
  assign g20641 = g35;
  assign g20642 = g35;
  assign g20648 = g35;
  assign g20649 = g35;
  assign g20650 = g35;
  assign g20651 = g35;
  assign g20652 = \DFF_1301.Q ;
  assign g20653 = \DFF_1301.Q ;
  assign g20654 = \DFF_1033.Q ;
  assign g20655 = \DFF_1033.Q ;
  assign g20656 = g35;
  assign g20657 = g35;
  assign g20659 = g35;
  assign g2066 = \DFF_1093.Q ;
  assign g20660 = g35;
  assign g20661 = g35;
  assign g20662 = g35;
  assign g20663 = g35;
  assign g20664 = g35;
  assign g20665 = g35;
  assign g20666 = g35;
  assign g20667 = g35;
  assign g20668 = g35;
  assign g20669 = g35;
  assign g20670 = g35;
  assign g20671 = g35;
  assign g20672 = g35;
  assign g20673 = g35;
  assign g20674 = g35;
  assign g20679 = g35;
  assign g20680 = g35;
  assign g20681 = g35;
  assign g20682 = g28753;
  assign g20695 = g25114;
  assign g20696 = g35;
  assign g20697 = g35;
  assign g20698 = g35;
  assign g20699 = g35;
  assign g2070 = \DFF_996.Q ;
  assign g20700 = g35;
  assign g20701 = g35;
  assign g20702 = g35;
  assign g20703 = g35;
  assign g20704 = g35;
  assign g20706 = g35;
  assign g20707 = g35;
  assign g20708 = g35;
  assign g20709 = g35;
  assign g20710 = g35;
  assign g20711 = g35;
  assign g20712 = g35;
  assign g20713 = g35;
  assign g20714 = g35;
  assign g20715 = g35;
  assign g20716 = g35;
  assign g20732 = g35;
  assign g20737 = g35;
  assign g20738 = g35;
  assign g20763 = \DFF_654.Q ;
  assign g20764 = \DFF_654.Q ;
  assign g20766 = g35;
  assign g20767 = g35;
  assign g20768 = g35;
  assign g20769 = g35;
  assign g20770 = g35;
  assign g20771 = g35;
  assign g20772 = g35;
  assign g20774 = g35;
  assign g20775 = g35;
  assign g20776 = g35;
  assign g20777 = g35;
  assign g20778 = g35;
  assign g20779 = g35;
  assign g20780 = g35;
  assign g2079 = \DFF_1310.Q ;
  assign g2084 = \DFF_1376.Q ;
  assign g20852 = g35;
  assign g20853 = g35;
  assign g20869 = g35;
  assign g20874 = g35;
  assign g2089 = \DFF_77.Q ;
  assign g20899 = \DFF_1044.Q ;
  assign g209 = \DFF_956.Q ;
  assign g20900 = \DFF_1044.Q ;
  assign g20901 = \DFF_357.Q ;
  assign g20902 = \DFF_357.Q ;
  assign g20903 = g35;
  assign g20904 = g35;
  assign g20909 = g35;
  assign g20910 = g35;
  assign g20911 = g35;
  assign g20912 = g35;
  assign g20913 = g35;
  assign g20914 = g35;
  assign g20916 = g35;
  assign g20917 = g35;
  assign g20918 = g35;
  assign g20919 = g35;
  assign g20920 = g35;
  assign g20921 = g35;
  assign g20923 = g35;
  assign g2093 = \DFF_1129.Q ;
  assign g20978 = g35;
  assign g2098 = \DFF_964.Q ;
  assign g20993 = g35;
  assign g20994 = g35;
  assign g21010 = g35;
  assign g2102 = \DFF_888.Q ;
  assign g21036 = g25167;
  assign g21048 = g35;
  assign g21049 = g35;
  assign g21050 = g35;
  assign g21051 = g35;
  assign g21052 = g35;
  assign g21053 = g35;
  assign g21054 = g35;
  assign g21055 = g35;
  assign g21056 = g35;
  assign g21057 = g35;
  assign g21058 = g35;
  assign g21059 = g35;
  assign g21060 = g35;
  assign g21068 = g35;
  assign g21069 = g35;
  assign g2108 = \DFF_1086.Q ;
  assign g2112 = \DFF_322.Q ;
  assign g21123 = g35;
  assign g21138 = g35;
  assign g21139 = g35;
  assign g21155 = g35;
  assign g21156 = g91;
  assign g2116 = \DFF_1261.Q ;
  assign g21160 = g126;
  assign g21175 = g26801;
  assign g21176 = \DFF_1059.Q ;
  assign g21177 = \DFF_1059.Q ;
  assign g21178 = g35;
  assign g21179 = g35;
  assign g21180 = g35;
  assign g21181 = g35;
  assign g21182 = g35;
  assign g21183 = g35;
  assign g21184 = g35;
  assign g21185 = g35;
  assign g21189 = g35;
  assign g21204 = g35;
  assign g21205 = g35;
  assign g2122 = \DFF_264.Q ;
  assign g21221 = g35;
  assign g21222 = g115;
  assign g21225 = g99;
  assign g21228 = \DFF_379.Q ;
  assign g21245 = \DFF_132.Q ;
  assign g21246 = \DFF_132.Q ;
  assign g21247 = g35;
  assign g21248 = g35;
  assign g21249 = g35;
  assign g21252 = g35;
  assign g2126 = \DFF_1213.Q ;
  assign g21267 = g35;
  assign g21268 = g35;
  assign g21269 = \DFF_743.Q ;
  assign g21270 = \DFF_125.Q ;
  assign g21271 = \DFF_125.Q ;
  assign g21274 = g35;
  assign g21275 = g35;
  assign g21279 = g35;
  assign g21281 = \DFF_206.Q ;
  assign g21282 = \DFF_141.Q ;
  assign g21286 = g35;
  assign g21291 = \DFF_420.Q ;
  assign g21292 = \DFF_489.Q ;
  assign g21293 = \DFF_489.Q ;
  assign g21295 = g35;
  assign g21299 = \DFF_1012.Q ;
  assign g2130 = \DFF_507.Q ;
  assign g21300 = g25259;
  assign g21304 = g35;
  assign g21305 = g35;
  assign g21308 = g84;
  assign g21329 = \DFF_1322.Q ;
  assign g21336 = g35;
  assign g21337 = g35;
  assign g21343 = \DFF_150.Q ;
  assign g21346 = g35;
  assign g21349 = g35;
  assign g21352 = \DFF_829.Q ;
  assign g21355 = g35;
  assign g21358 = \DFF_477.Q ;
  assign g21362 = g35;
  assign g21366 = g23002;
  assign g21369 = \DFF_514.Q ;
  assign g21370 = g54;
  assign g21379 = g35;
  assign g2138 = \DFF_941.Q ;
  assign g21380 = g35;
  assign g21381 = g35;
  assign g21383 = g35;
  assign g21395 = g35;
  assign g21396 = g35;
  assign g21397 = g35;
  assign g21398 = g35;
  assign g21399 = g35;
  assign g21400 = g35;
  assign g21406 = g35;
  assign g21407 = g35;
  assign g21408 = g35;
  assign g21409 = g35;
  assign g21410 = g35;
  assign g21411 = g35;
  assign g21412 = g35;
  assign g21414 = g35;
  assign g21418 = g35;
  assign g21421 = g35;
  assign g21422 = g35;
  assign g21423 = g35;
  assign g21424 = g35;
  assign g21425 = g35;
  assign g21426 = g35;
  assign g21427 = g35;
  assign g21428 = g35;
  assign g21431 = g35;
  assign g21434 = \DFF_1181.Q ;
  assign g2145 = \DFF_445.Q ;
  assign g21451 = g27831;
  assign g21454 = g35;
  assign g21455 = g35;
  assign g21456 = g35;
  assign g21457 = g35;
  assign g21458 = g35;
  assign g21461 = g35;
  assign g21463 = \DFF_304.Q ;
  assign g21466 = g35;
  assign g21467 = g35;
  assign g215 = \DFF_612.Q ;
  assign g2151 = \DFF_680.Q ;
  assign g21511 = g35;
  assign g2152 = \DFF_391.Q ;
  assign g2153 = \DFF_769.Q ;
  assign g21560 = g35;
  assign g21561 = g35;
  assign g21604 = g35;
  assign g21607 = g35;
  assign g21608 = g35;
  assign g21609 = g35;
  assign g2161 = \DFF_1231.Q ;
  assign g21610 = g35;
  assign g2165 = \DFF_1096.Q ;
  assign g21665 = \DFF_748.Q ;
  assign g21669 = \DFF_748.Q ;
  assign g21673 = \DFF_748.Q ;
  assign g21677 = \DFF_748.Q ;
  assign g21681 = \DFF_748.Q ;
  assign g21685 = \DFF_748.Q ;
  assign g21689 = \DFF_748.Q ;
  assign g2169 = \DFF_1030.Q ;
  assign g21693 = \DFF_748.Q ;
  assign g21697 = \DFF_748.Q ;
  assign g21698 = g36;
  assign g21722 = \DFF_800.D ;
  assign g21723 = \DFF_999.D ;
  assign g21724 = \DFF_1292.D ;
  assign g21725 = \DFF_1353.D ;
  assign g21726 = \DFF_1381.D ;
  assign g2173 = \DFF_1026.Q ;
  assign g2177 = \DFF_204.Q ;
  assign g218 = \DFF_1061.Q ;
  assign g2181 = \DFF_1135.Q ;
  assign g2185 = \DFF_993.Q ;
  assign g21891 = \DFF_389.D ;
  assign g21892 = \DFF_1387.D ;
  assign g21893 = \DFF_1190.D ;
  assign g21894 = \DFF_73.D ;
  assign g21895 = \DFF_215.D ;
  assign g21896 = \DFF_831.D ;
  assign g21897 = \DFF_1384.D ;
  assign g21898 = \DFF_1027.D ;
  assign g21899 = \DFF_858.D ;
  assign g21900 = \DFF_739.D ;
  assign g21901 = \DFF_1234.D ;
  assign g21902 = \DFF_501.D ;
  assign g21903 = \DFF_200.D ;
  assign g21904 = \DFF_1402.D ;
  assign g21905 = \DFF_1165.D ;
  assign g2193 = \DFF_570.Q ;
  assign g2197 = \DFF_1141.Q ;
  assign g22 = \DFF_748.Q ;
  assign g2204 = \DFF_658.Q ;
  assign g2208 = \DFF_889.Q ;
  assign g22144 = g35;
  assign g22146 = g35;
  assign g22147 = g35;
  assign g22148 = g35;
  assign g22153 = g35;
  assign g22154 = g35;
  assign g22155 = g35;
  assign g22156 = g35;
  assign g22166 = g35;
  assign g22167 = g35;
  assign g22168 = g35;
  assign g22169 = g35;
  assign g2217 = \DFF_1091.Q ;
  assign g22170 = g35;
  assign g22173 = g84;
  assign g22176 = g35;
  assign g22177 = g35;
  assign g22178 = g35;
  assign g22179 = g35;
  assign g22180 = g35;
  assign g22181 = g35;
  assign g22182 = g72;
  assign g22192 = g35;
  assign g22194 = g84;
  assign g22197 = g35;
  assign g22198 = g35;
  assign g22199 = g35;
  assign g222 = \DFF_258.Q ;
  assign g22200 = g35;
  assign g22201 = g35;
  assign g22202 = g73;
  assign g22210 = g84;
  assign g22213 = g35;
  assign g22214 = g35;
  assign g22215 = g35;
  assign g22220 = g84;
  assign g22223 = g35;
  assign g22224 = g35;
  assign g22227 = g35;
  assign g2223 = \DFF_462.Q ;
  assign g2227 = \DFF_1047.Q ;
  assign g22300 = g84;
  assign g22303 = g35;
  assign g22305 = g35;
  assign g22317 = g35;
  assign g22330 = g35;
  assign g22338 = g35;
  assign g22339 = g35;
  assign g22341 = g35;
  assign g22358 = g35;
  assign g2236 = \DFF_37.Q ;
  assign g22360 = g72;
  assign g22409 = g73;
  assign g2241 = \DFF_374.Q ;
  assign g22455 = g35;
  assign g22456 = g35;
  assign g2246 = \DFF_1050.Q ;
  assign g22493 = g35;
  assign g22494 = g35;
  assign g22495 = g35;
  assign g225 = \DFF_382.Q ;
  assign g2250 = \DFF_1328.Q ;
  assign g22519 = g35;
  assign g22520 = g35;
  assign g22526 = g35;
  assign g22528 = g35;
  assign g22542 = g35;
  assign g22543 = g35;
  assign g2255 = \DFF_301.Q ;
  assign g2259 = \DFF_232.Q ;
  assign g22593 = g35;
  assign g22635 = g35;
  assign g22647 = g53;
  assign g2265 = \DFF_903.Q ;
  assign g22658 = g54;
  assign g22683 = g56;
  assign g2269 = \DFF_841.Q ;
  assign g22698 = \DFF_743.Q ;
  assign g22721 = g57;
  assign g2273 = \DFF_835.Q ;
  assign g22758 = g35;
  assign g22763 = g113;
  assign g2279 = \DFF_558.Q ;
  assign g2283 = \DFF_1031.Q ;
  assign g22830 = g35;
  assign g22840 = g35;
  assign g22841 = g35;
  assign g22847 = g35;
  assign g22854 = g35;
  assign g22855 = g35;
  assign g22856 = g35;
  assign g22865 = g35;
  assign g22866 = g35;
  assign g22867 = g35;
  assign g22868 = g35;
  assign g2287 = \DFF_209.Q ;
  assign g22882 = g35;
  assign g22883 = g35;
  assign g22884 = g35;
  assign g22898 = g35;
  assign g22903 = g35;
  assign g22906 = g35;
  assign g22907 = g35;
  assign g22922 = g35;
  assign g22923 = g25259;
  assign g22926 = g35;
  assign g22935 = g35;
  assign g22936 = g35;
  assign g2295 = \DFF_65.Q ;
  assign g22973 = g35;
  assign g22974 = g35;
  assign g22975 = g35;
  assign g22976 = g25167;
  assign g22979 = g35;
  assign g22981 = g35;
  assign g22985 = g35;
  assign g22986 = g35;
  assign g22987 = g35;
  assign g22988 = g35;
  assign g22989 = g35;
  assign g2299 = \DFF_4.Q ;
  assign g22995 = g35;
  assign g22996 = g35;
  assign g22997 = g35;
  assign g22998 = g35;
  assign g22999 = g35;
  assign g23000 = g35;
  assign g23001 = g35;
  assign g23003 = g23002;
  assign g23004 = g35;
  assign g23005 = g35;
  assign g23011 = g35;
  assign g23012 = g35;
  assign g23013 = g35;
  assign g23014 = g35;
  assign g23015 = g35;
  assign g23016 = g35;
  assign g23017 = g35;
  assign g23018 = g35;
  assign g23019 = \DFF_748.Q ;
  assign g23020 = \DFF_748.Q ;
  assign g23021 = g35;
  assign g23022 = g35;
  assign g23026 = g35;
  assign g23027 = g35;
  assign g23028 = g35;
  assign g23029 = g35;
  assign g2303 = \DFF_1247.Q ;
  assign g23030 = g35;
  assign g23031 = g35;
  assign g23032 = \DFF_304.Q ;
  assign g23041 = \DFF_748.Q ;
  assign g23046 = g35;
  assign g23057 = g35;
  assign g23058 = g35;
  assign g23059 = g35;
  assign g23060 = \DFF_748.Q ;
  assign g23061 = g35;
  assign g23066 = g35;
  assign g2307 = \DFF_457.Q ;
  assign g23084 = \DFF_748.Q ;
  assign g23085 = \DFF_748.Q ;
  assign g23086 = g35;
  assign g2311 = \DFF_625.Q ;
  assign g23111 = g35;
  assign g23128 = g35;
  assign g23138 = g35;
  assign g2315 = \DFF_469.Q ;
  assign g23152 = g35;
  assign g23170 = \DFF_748.Q ;
  assign g23189 = \DFF_748.Q ;
  assign g2319 = \DFF_387.Q ;
  assign g23191 = g23190;
  assign g23196 = g35;
  assign g232 = \DFF_496.Q ;
  assign g23203 = \DFF_748.Q ;
  assign g23214 = g35;
  assign g23215 = g35;
  assign g23216 = g35;
  assign g23221 = g35;
  assign g23222 = g35;
  assign g23226 = g35;
  assign g23227 = g35;
  assign g23228 = g35;
  assign g23232 = g64;
  assign g23233 = g35;
  assign g23235 = g35;
  assign g23236 = g35;
  assign g23237 = g35;
  assign g23238 = g35;
  assign g23242 = g35;
  assign g23243 = g35;
  assign g23245 = g35;
  assign g23246 = g35;
  assign g23247 = g35;
  assign g23248 = g35;
  assign g23249 = g35;
  assign g23250 = g35;
  assign g23253 = g35;
  assign g23256 = g35;
  assign g23257 = g35;
  assign g23258 = g35;
  assign g23259 = g35;
  assign g23260 = g35;
  assign g23263 = g90;
  assign g23264 = g35;
  assign g2327 = \DFF_1240.Q ;
  assign g23270 = g35;
  assign g23271 = g35;
  assign g23272 = g35;
  assign g23273 = g35;
  assign g23274 = g35;
  assign g23277 = g91;
  assign g23278 = g35;
  assign g23279 = g35;
  assign g23282 = g35;
  assign g23283 = g35;
  assign g23284 = g35;
  assign g23289 = g35;
  assign g23290 = g35;
  assign g23291 = g35;
  assign g23299 = g72;
  assign g23300 = g35;
  assign g23301 = g35;
  assign g23302 = g35;
  assign g23303 = g35;
  assign g23304 = g35;
  assign g23305 = g35;
  assign g23306 = g35;
  assign g23307 = g35;
  assign g2331 = \DFF_1010.Q ;
  assign g23312 = g35;
  assign g23313 = g35;
  assign g23320 = g73;
  assign g23321 = g113;
  assign g23322 = g124;
  assign g23323 = g35;
  assign g23332 = g35;
  assign g23333 = g35;
  assign g23334 = g35;
  assign g23335 = g35;
  assign g23336 = g35;
  assign g23337 = g35;
  assign g23338 = g35;
  assign g23339 = g35;
  assign g23340 = g35;
  assign g23347 = g114;
  assign g23350 = g35;
  assign g23351 = g35;
  assign g23352 = g35;
  assign g23353 = g35;
  assign g23354 = g35;
  assign g23355 = g35;
  assign g23356 = g35;
  assign g23359 = g92;
  assign g23360 = g99;
  assign g23361 = g115;
  assign g23362 = g125;
  assign g23375 = g35;
  assign g23376 = g35;
  assign g23377 = g35;
  assign g23378 = g35;
  assign g2338 = \DFF_943.Q ;
  assign g23384 = g84;
  assign g23385 = g100;
  assign g23388 = g35;
  assign g23390 = g35;
  assign g23394 = g126;
  assign g23395 = g127;
  assign g23398 = g35;
  assign g23399 = g35;
  assign g23403 = g116;
  assign g23406 = g35;
  assign g23408 = g35;
  assign g23409 = g35;
  assign g23410 = g35;
  assign g23414 = g134;
  assign g23417 = g35;
  assign g23418 = g35;
  assign g23419 = g35;
  assign g2342 = \DFF_297.Q ;
  assign g23420 = g35;
  assign g23421 = g35;
  assign g23422 = g35;
  assign g23426 = g120;
  assign g23427 = g135;
  assign g23429 = g35;
  assign g23431 = g35;
  assign g23432 = g35;
  assign g23433 = g35;
  assign g23434 = g35;
  assign g23435 = g35;
  assign g23440 = g25114;
  assign g23443 = g35;
  assign g23446 = g35;
  assign g23447 = g35;
  assign g23448 = g35;
  assign g23449 = g35;
  assign g23450 = g44;
  assign g23452 = g35;
  assign g23453 = \DFF_141.Q ;
  assign g23456 = g35;
  assign g23459 = g35;
  assign g23460 = g35;
  assign g23461 = g35;
  assign g23473 = g35;
  assign g23476 = g35;
  assign g23477 = g35;
  assign g23478 = g35;
  assign g23479 = g35;
  assign g23482 = g35;
  assign g23483 = g35;
  assign g23485 = g35;
  assign g23486 = g35;
  assign g23487 = g35;
  assign g23488 = g35;
  assign g23489 = g35;
  assign g23490 = g35;
  assign g23491 = g35;
  assign g23492 = g35;
  assign g23493 = g35;
  assign g23499 = g35;
  assign g23500 = g35;
  assign g23501 = g35;
  assign g23502 = g35;
  assign g23503 = g35;
  assign g23504 = g35;
  assign g23505 = g35;
  assign g23506 = g35;
  assign g23507 = g35;
  assign g23508 = g35;
  assign g23509 = g35;
  assign g2351 = \DFF_681.Q ;
  assign g23510 = g35;
  assign g23515 = g35;
  assign g23516 = g35;
  assign g23517 = g35;
  assign g23518 = g35;
  assign g23519 = g35;
  assign g23520 = g35;
  assign g23521 = g35;
  assign g23522 = g35;
  assign g23523 = g35;
  assign g23524 = g35;
  assign g23525 = g35;
  assign g23526 = g35;
  assign g23527 = g35;
  assign g23528 = g35;
  assign g23534 = g84;
  assign g23537 = g35;
  assign g23538 = g35;
  assign g23539 = g35;
  assign g23541 = g35;
  assign g23542 = g35;
  assign g23543 = g35;
  assign g23544 = g35;
  assign g23545 = g35;
  assign g23546 = g35;
  assign g23547 = g35;
  assign g23548 = g35;
  assign g23549 = g35;
  assign g23555 = g84;
  assign g23558 = g35;
  assign g23559 = g35;
  assign g23565 = g35;
  assign g23566 = g35;
  assign g23567 = g35;
  assign g23568 = g35;
  assign g23569 = g35;
  assign g2357 = \DFF_1337.Q ;
  assign g23570 = g35;
  assign g23571 = g35;
  assign g23582 = g84;
  assign g23585 = g35;
  assign g23589 = g35;
  assign g23607 = g35;
  assign g23608 = g35;
  assign g23609 = g35;
  assign g2361 = \DFF_1233.Q ;
  assign g23610 = g35;
  assign g23611 = g35;
  assign g23613 = g23612;
  assign g23629 = g35;
  assign g23647 = g35;
  assign g23648 = g35;
  assign g23649 = g35;
  assign g23653 = g23652;
  assign g23665 = g35;
  assign g23683 = \DFF_828.Q ;
  assign g23684 = \DFF_828.Q ;
  assign g23698 = g35;
  assign g2370 = \DFF_406.Q ;
  assign g23732 = g35;
  assign g23749 = g35;
  assign g2375 = \DFF_795.Q ;
  assign g23760 = g23759;
  assign g23767 = g35;
  assign g23768 = g35;
  assign g23769 = g35;
  assign g23777 = g27831;
  assign g23787 = g35;
  assign g23788 = g35;
  assign g23792 = g35;
  assign g23793 = g35;
  assign g23794 = g35;
  assign g2380 = \DFF_637.Q ;
  assign g23812 = g35;
  assign g23813 = g35;
  assign g23814 = g35;
  assign g23815 = g35;
  assign g23819 = g35;
  assign g23820 = g35;
  assign g23821 = g35;
  assign g23823 = g26801;
  assign g23838 = g35;
  assign g23839 = g35;
  assign g2384 = \DFF_804.Q ;
  assign g23840 = g35;
  assign g23841 = g35;
  assign g23842 = g35;
  assign g23843 = g35;
  assign g23847 = g35;
  assign g23848 = g35;
  assign g23849 = g35;
  assign g23858 = g35;
  assign g23859 = g35;
  assign g23860 = g35;
  assign g23861 = g35;
  assign g23862 = g35;
  assign g23863 = g35;
  assign g23864 = g35;
  assign g23868 = g35;
  assign g23869 = g35;
  assign g23870 = g23612;
  assign g23874 = g35;
  assign g23875 = g35;
  assign g23876 = g35;
  assign g23877 = g35;
  assign g23878 = g35;
  assign g23879 = g35;
  assign g23880 = g35;
  assign g23881 = g35;
  assign g23882 = g35;
  assign g23886 = g35;
  assign g23887 = g35;
  assign g23888 = g35;
  assign g2389 = \DFF_928.Q ;
  assign g23893 = g35;
  assign g23894 = g35;
  assign g23895 = g35;
  assign g23896 = g35;
  assign g23897 = g35;
  assign g23898 = g35;
  assign g23899 = g35;
  assign g239 = \DFF_362.Q ;
  assign g23902 = g35;
  assign g23903 = g35;
  assign g23904 = g35;
  assign g23905 = g35;
  assign g23906 = g35;
  assign g23907 = g35;
  assign g23912 = g35;
  assign g23913 = g35;
  assign g23914 = g35;
  assign g23915 = g35;
  assign g23916 = g35;
  assign g23922 = g35;
  assign g23923 = g35;
  assign g23924 = g35;
  assign g23925 = g35;
  assign g23926 = g35;
  assign g23927 = g35;
  assign g23928 = g35;
  assign g23929 = g35;
  assign g2393 = \DFF_571.Q ;
  assign g23930 = g35;
  assign g23935 = g35;
  assign g23936 = g35;
  assign g23937 = g35;
  assign g23938 = g35;
  assign g23939 = g35;
  assign g23940 = g35;
  assign g23941 = g35;
  assign g23942 = g35;
  assign g23943 = g35;
  assign g23944 = g35;
  assign g23945 = g35;
  assign g23946 = g35;
  assign g23947 = g35;
  assign g23952 = g35;
  assign g23953 = g35;
  assign g23954 = g28753;
  assign g23961 = g35;
  assign g23962 = g35;
  assign g23963 = g35;
  assign g23964 = g35;
  assign g23965 = g35;
  assign g23966 = g35;
  assign g23967 = g35;
  assign g23968 = g35;
  assign g23969 = g35;
  assign g23970 = g35;
  assign g23982 = g35;
  assign g23983 = g35;
  assign g23984 = g35;
  assign g23985 = g35;
  assign g23986 = g35;
  assign g23987 = g35;
  assign g23988 = g35;
  assign g2399 = \DFF_216.Q ;
  assign g23992 = g35;
  assign g23993 = g35;
  assign g23994 = g35;
  assign g23995 = g35;
  assign g23999 = g35;
  assign g24000 = g35;
  assign g24003 = g35;
  assign g24010 = g35;
  assign g24013 = g35;
  assign g24017 = g35;
  assign g2403 = \DFF_444.Q ;
  assign g2407 = \DFF_1034.Q ;
  assign g2413 = \DFF_1276.Q ;
  assign g24151 = 1'b1;
  assign g24152 = \DFF_748.Q ;
  assign g24153 = \DFF_748.Q ;
  assign g24154 = \DFF_748.Q ;
  assign g24155 = \DFF_748.Q ;
  assign g24156 = \DFF_748.Q ;
  assign g24157 = \DFF_748.Q ;
  assign g24158 = \DFF_748.Q ;
  assign g24159 = \DFF_748.Q ;
  assign g24160 = \DFF_748.Q ;
  assign g24161 = g53;
  assign g24162 = g54;
  assign g24163 = g56;
  assign g24164 = g57;
  assign g24165 = g64;
  assign g24166 = g72;
  assign g24167 = g73;
  assign g24168 = g84;
  assign g24169 = g90;
  assign g2417 = \DFF_499.Q ;
  assign g24170 = g91;
  assign g24171 = g92;
  assign g24172 = g99;
  assign g24173 = g100;
  assign g24174 = g113;
  assign g24175 = g114;
  assign g24176 = g115;
  assign g24177 = g116;
  assign g24178 = g120;
  assign g24179 = g124;
  assign g24180 = g125;
  assign g24181 = g126;
  assign g24182 = g127;
  assign g24183 = g134;
  assign g24184 = g135;
  assign g24185 = g44;
  assign g24200 = \DFF_1053.D ;
  assign g24201 = \DFF_601.D ;
  assign g24202 = \DFF_1108.D ;
  assign g24203 = \DFF_542.D ;
  assign g24204 = \DFF_972.D ;
  assign g24205 = \DFF_324.D ;
  assign g24206 = \DFF_239.D ;
  assign g24207 = \DFF_544.D ;
  assign g24208 = \DFF_510.D ;
  assign g24209 = \DFF_237.D ;
  assign g2421 = \DFF_1143.Q ;
  assign g24210 = \DFF_252.D ;
  assign g24211 = \DFF_597.D ;
  assign g24212 = \DFF_752.D ;
  assign g24213 = \DFF_515.D ;
  assign g24214 = \DFF_667.D ;
  assign g24215 = \DFF_872.D ;
  assign g24216 = \DFF_23.D ;
  assign g24229 = \DFF_908.D ;
  assign g24231 = \DFF_880.D ;
  assign g24232 = \DFF_24.D ;
  assign g24233 = \DFF_580.D ;
  assign g24234 = \DFF_1094.D ;
  assign g24235 = \DFF_98.D ;
  assign g24236 = \DFF_133.D ;
  assign g24237 = \DFF_208.D ;
  assign g24238 = \DFF_711.D ;
  assign g24239 = \DFF_185.D ;
  assign g24240 = \DFF_675.D ;
  assign g24241 = \DFF_1207.D ;
  assign g24242 = \DFF_339.D ;
  assign g24243 = \DFF_606.D ;
  assign g24244 = \DFF_90.D ;
  assign g24245 = \DFF_343.D ;
  assign g24246 = \DFF_1057.D ;
  assign g24247 = \DFF_871.D ;
  assign g24248 = \DFF_1092.D ;
  assign g24249 = \DFF_822.D ;
  assign g24250 = \DFF_167.D ;
  assign g24251 = \DFF_182.D ;
  assign g24252 = \DFF_1407.D ;
  assign g24253 = \DFF_202.D ;
  assign g24254 = \DFF_422.D ;
  assign g24255 = \DFF_1072.D ;
  assign g24256 = \DFF_60.D ;
  assign g24257 = \DFF_937.D ;
  assign g24258 = \DFF_1275.D ;
  assign g24259 = \DFF_67.D ;
  assign g24260 = \DFF_1371.D ;
  assign g24261 = \DFF_395.D ;
  assign g24262 = \DFF_375.D ;
  assign g24263 = \DFF_962.D ;
  assign g24264 = \DFF_126.D ;
  assign g24265 = \DFF_448.D ;
  assign g24266 = \DFF_843.D ;
  assign g24267 = \DFF_819.D ;
  assign g24268 = \DFF_538.D ;
  assign g24269 = \DFF_224.D ;
  assign g24270 = \DFF_840.D ;
  assign g24271 = \DFF_1420.D ;
  assign g24272 = \DFF_664.D ;
  assign g24273 = \DFF_1214.D ;
  assign g24274 = \DFF_39.D ;
  assign g24275 = \DFF_1001.D ;
  assign g24276 = \DFF_5.D ;
  assign g24277 = \DFF_423.D ;
  assign g24278 = \DFF_347.D ;
  assign g24279 = \DFF_919.D ;
  assign g24280 = \DFF_210.D ;
  assign g24281 = \DFF_203.D ;
  assign g24282 = \DFF_349.D ;
  assign g2429 = \DFF_930.Q ;
  assign g24298 = \DFF_1305.D ;
  assign g2433 = \DFF_273.Q ;
  assign g24334 = \DFF_934.D ;
  assign g24335 = \DFF_607.D ;
  assign g24336 = \DFF_165.D ;
  assign g24337 = \DFF_141.D ;
  assign g24338 = \DFF_1400.D ;
  assign g24339 = \DFF_1285.D ;
  assign g24340 = \DFF_46.D ;
  assign g24341 = \DFF_599.D ;
  assign g24342 = \DFF_1162.D ;
  assign g24343 = \DFF_1404.D ;
  assign g24344 = \DFF_30.D ;
  assign g24345 = \DFF_1320.D ;
  assign g24346 = \DFF_543.D ;
  assign g24347 = \DFF_731.D ;
  assign g24348 = \DFF_554.D ;
  assign g24349 = \DFF_1005.D ;
  assign g24350 = \DFF_251.D ;
  assign g24351 = \DFF_1188.D ;
  assign g24352 = \DFF_1158.D ;
  assign g24353 = \DFF_198.D ;
  assign g24354 = \DFF_1130.D ;
  assign g24355 = \DFF_683.D ;
  assign g24356 = g35;
  assign g24358 = g35;
  assign g24359 = g35;
  assign g24360 = g35;
  assign g24364 = g35;
  assign g24365 = g35;
  assign g24366 = g35;
  assign g24367 = g35;
  assign g24368 = g35;
  assign g2437 = \DFF_887.Q ;
  assign g24375 = g35;
  assign g24376 = g35;
  assign g24377 = g35;
  assign g24379 = g35;
  assign g24386 = g35;
  assign g24394 = g35;
  assign g24405 = g35;
  assign g24407 = g35;
  assign g2441 = \DFF_1171.Q ;
  assign g24417 = \DFF_934.Q ;
  assign g24418 = g35;
  assign g24419 = g35;
  assign g24424 = g35;
  assign g24425 = g35;
  assign g24426 = g35;
  assign g24428 = g35;
  assign g24429 = g35;
  assign g24431 = g35;
  assign g24438 = g35;
  assign g2445 = \DFF_1025.Q ;
  assign g24452 = g35;
  assign g2449 = \DFF_959.Q ;
  assign g24490 = g35;
  assign g2453 = \DFF_1331.Q ;
  assign g24575 = \DFF_1220.D ;
  assign g246 = \DFF_346.Q ;
  assign g2461 = \DFF_425.Q ;
  assign g24619 = \DFF_1111.D ;
  assign g2465 = \DFF_265.Q ;
  assign g2472 = \DFF_1254.Q ;
  assign g24759 = \DFF_994.Q ;
  assign g2476 = \DFF_793.Q ;
  assign g24819 = g72;
  assign g24836 = g72;
  assign g2485 = \DFF_148.Q ;
  assign g24850 = g72;
  assign g24866 = g73;
  assign g24869 = g72;
  assign g24891 = \DFF_1425.Q ;
  assign g24893 = g73;
  assign g2491 = \DFF_1028.Q ;
  assign g24911 = g72;
  assign g24920 = g73;
  assign g2495 = \DFF_886.Q ;
  assign g25027 = g72;
  assign g2504 = \DFF_989.Q ;
  assign g25051 = g72;
  assign g25064 = g73;
  assign g25067 = \DFF_161.Q ;
  assign g25073 = g26801;
  assign g25084 = \DFF_177.Q ;
  assign g25085 = \DFF_766.Q ;
  assign g2509 = \DFF_1115.Q ;
  assign g25102 = \DFF_1157.Q ;
  assign g25103 = \DFF_231.Q ;
  assign g25115 = g25114;
  assign g25123 = \DFF_677.Q ;
  assign g25124 = \DFF_276.Q ;
  assign g2514 = \DFF_442.Q ;
  assign g25140 = g35;
  assign g25142 = \DFF_1193.Q ;
  assign g25143 = \DFF_721.Q ;
  assign g25158 = g35;
  assign g25159 = \DFF_855.Q ;
  assign g25168 = g25167;
  assign g25171 = g35;
  assign g2518 = \DFF_726.Q ;
  assign g25180 = \DFF_1078.Q ;
  assign g25185 = g35;
  assign g25198 = g35;
  assign g25206 = \DFF_489.Q ;
  assign g25214 = g35;
  assign g25219 = \DFF_141.Q ;
  assign g25220 = \DFF_141.Q ;
  assign g25221 = \DFF_576.Q ;
  assign g25222 = g28753;
  assign g2523 = \DFF_818.Q ;
  assign g25231 = g35;
  assign g25232 = g35;
  assign g25240 = \DFF_1301.Q ;
  assign g25241 = \DFF_1033.Q ;
  assign g25248 = g35;
  assign g25249 = g35;
  assign g25250 = g113;
  assign g25260 = g25259;
  assign g25266 = g35;
  assign g25267 = g35;
  assign g2527 = \DFF_1395.Q ;
  assign g25272 = \DFF_654.Q ;
  assign g25286 = g35;
  assign g25287 = g35;
  assign g25288 = g35;
  assign g25289 = g35;
  assign g25296 = \DFF_1044.Q ;
  assign g25297 = \DFF_357.Q ;
  assign g25298 = \DFF_865.Q ;
  assign g25324 = g35;
  assign g25325 = g35;
  assign g25326 = g35;
  assign g2533 = \DFF_1268.Q ;
  assign g25369 = g35;
  assign g2537 = \DFF_488.Q ;
  assign g25370 = g35;
  assign g25380 = \DFF_1059.Q ;
  assign g25409 = g35;
  assign g2541 = \DFF_768.Q ;
  assign g25410 = g35;
  assign g25423 = g27831;
  assign g25424 = \DFF_132.Q ;
  assign g25448 = g31521;
  assign g25451 = g35;
  assign g25452 = g35;
  assign g25465 = \DFF_125.Q ;
  assign g2547 = \DFF_6.Q ;
  assign g25480 = g35;
  assign g25481 = g35;
  assign g255 = \DFF_771.Q ;
  assign g25505 = g35;
  assign g25506 = g35;
  assign g2551 = \DFF_825.Q ;
  assign g25513 = \DFF_489.Q ;
  assign g25517 = g35;
  assign g25523 = g35;
  assign g25524 = g35;
  assign g25525 = g35;
  assign g25528 = g35;
  assign g25531 = g31665;
  assign g25533 = g35;
  assign g25537 = g31656;
  assign g25538 = g35;
  assign g25544 = g35;
  assign g25546 = g35;
  assign g25547 = g35;
  assign g25548 = g35;
  assign g2555 = \DFF_713.Q ;
  assign g25552 = g35;
  assign g25553 = g35;
  assign g25554 = g35;
  assign g25555 = g35;
  assign g25558 = g35;
  assign g25560 = g35;
  assign g25561 = g35;
  assign g25563 = g35;
  assign g25566 = g35;
  assign g25582 = 1'b1;
  assign g25583 = 1'b1;
  assign g25584 = 1'b1;
  assign g25585 = 1'b1;
  assign g25586 = 1'b1;
  assign g25587 = 1'b1;
  assign g25588 = 1'b1;
  assign g25589 = 1'b1;
  assign g25590 = 1'b1;
  assign g25591 = \DFF_612.D ;
  assign g25592 = \DFF_824.D ;
  assign g25593 = \DFF_956.D ;
  assign g25594 = \DFF_128.D ;
  assign g25595 = \DFF_269.D ;
  assign g25596 = \DFF_1232.D ;
  assign g25597 = \DFF_1161.D ;
  assign g25598 = \DFF_1393.D ;
  assign g25599 = \DFF_96.D ;
  assign g25600 = \DFF_533.D ;
  assign g25601 = \DFF_292.D ;
  assign g25602 = \DFF_1045.D ;
  assign g25603 = \DFF_427.D ;
  assign g25604 = \DFF_10.D ;
  assign g25605 = \DFF_652.D ;
  assign g25606 = \DFF_629.D ;
  assign g25607 = \DFF_11.D ;
  assign g25608 = \DFF_430.D ;
  assign g25609 = \DFF_786.D ;
  assign g25610 = \DFF_622.D ;
  assign g25611 = \DFF_447.D ;
  assign g25612 = \DFF_591.D ;
  assign g25613 = \DFF_88.D ;
  assign g25614 = \DFF_900.D ;
  assign g25615 = \DFF_866.D ;
  assign g25616 = \DFF_988.D ;
  assign g25617 = \DFF_870.D ;
  assign g25618 = \DFF_525.D ;
  assign g25619 = \DFF_113.D ;
  assign g25620 = \DFF_908.D ;
  assign g25621 = \DFF_94.D ;
  assign g25622 = \DFF_283.D ;
  assign g25623 = \DFF_979.D ;
  assign g25624 = \DFF_486.D ;
  assign g25625 = \DFF_261.D ;
  assign g25626 = \DFF_1136.D ;
  assign g25627 = \DFF_416.D ;
  assign g25628 = \DFF_1103.D ;
  assign g25629 = \DFF_363.D ;
  assign g2563 = \DFF_61.Q ;
  assign g25630 = \DFF_1017.D ;
  assign g25631 = \DFF_1039.D ;
  assign g25632 = \DFF_1343.D ;
  assign g25633 = \DFF_66.D ;
  assign g25634 = \DFF_1008.D ;
  assign g25635 = \DFF_1323.D ;
  assign g25636 = \DFF_1131.D ;
  assign g25637 = \DFF_1194.D ;
  assign g25638 = \DFF_1313.D ;
  assign g25639 = \DFF_893.D ;
  assign g25640 = \DFF_126.D ;
  assign g25641 = \DFF_448.D ;
  assign g25642 = \DFF_843.D ;
  assign g25643 = \DFF_1318.D ;
  assign g25644 = \DFF_827.D ;
  assign g25645 = \DFF_775.D ;
  assign g25646 = \DFF_1156.D ;
  assign g25647 = \DFF_1076.D ;
  assign g25648 = \DFF_317.D ;
  assign g25649 = \DFF_1256.D ;
  assign g25650 = \DFF_259.D ;
  assign g25651 = \DFF_205.D ;
  assign g25652 = \DFF_1249.D ;
  assign g25653 = \DFF_1342.D ;
  assign g25654 = \DFF_356.D ;
  assign g25655 = \DFF_222.D ;
  assign g25656 = \DFF_124.D ;
  assign g25657 = \DFF_578.D ;
  assign g25658 = \DFF_801.D ;
  assign g25659 = \DFF_1168.D ;
  assign g25660 = \DFF_437.D ;
  assign g25661 = \DFF_180.D ;
  assign g25662 = \DFF_830.D ;
  assign g25663 = \DFF_1414.D ;
  assign g25664 = \DFF_1298.D ;
  assign g25665 = \DFF_805.D ;
  assign g25666 = \DFF_1405.D ;
  assign g25667 = \DFF_589.D ;
  assign g25668 = \DFF_29.D ;
  assign g25669 = \DFF_243.D ;
  assign g2567 = \DFF_727.Q ;
  assign g25670 = \DFF_1134.D ;
  assign g25671 = \DFF_495.D ;
  assign g25672 = \DFF_701.D ;
  assign g25673 = \DFF_939.D ;
  assign g25674 = \DFF_523.D ;
  assign g25675 = \DFF_540.D ;
  assign g25676 = \DFF_147.D ;
  assign g25677 = \DFF_460.D ;
  assign g25678 = \DFF_478.D ;
  assign g25679 = \DFF_405.D ;
  assign g25680 = \DFF_631.D ;
  assign g25681 = \DFF_1360.D ;
  assign g25682 = \DFF_1383.D ;
  assign g25683 = \DFF_1260.D ;
  assign g25684 = \DFF_87.D ;
  assign g25685 = \DFF_891.D ;
  assign g25686 = \DFF_1324.D ;
  assign g25687 = \DFF_1361.D ;
  assign g25688 = \DFF_527.D ;
  assign g25689 = \DFF_434.D ;
  assign g25690 = \DFF_1204.D ;
  assign g25691 = \DFF_685.D ;
  assign g25692 = \DFF_1305.D ;
  assign g25693 = \DFF_178.D ;
  assign g25694 = \DFF_672.D ;
  assign g25695 = \DFF_722.D ;
  assign g25696 = \DFF_883.D ;
  assign g25697 = \DFF_248.D ;
  assign g25698 = \DFF_1217.D ;
  assign g25699 = \DFF_1078.D ;
  assign g25700 = \DFF_678.D ;
  assign g25701 = \DFF_545.D ;
  assign g25702 = \DFF_1065.D ;
  assign g25703 = \DFF_366.D ;
  assign g25704 = \DFF_288.D ;
  assign g25705 = \DFF_1370.D ;
  assign g25706 = \DFF_1398.D ;
  assign g25707 = \DFF_1284.D ;
  assign g25708 = \DFF_926.D ;
  assign g25709 = \DFF_285.D ;
  assign g2571 = \DFF_1097.Q ;
  assign g25710 = \DFF_605.D ;
  assign g25711 = \DFF_354.D ;
  assign g25712 = \DFF_691.D ;
  assign g25713 = \DFF_556.D ;
  assign g25714 = \DFF_630.D ;
  assign g25715 = \DFF_503.D ;
  assign g25716 = \DFF_539.D ;
  assign g25717 = \DFF_1392.D ;
  assign g25718 = \DFF_668.D ;
  assign g25719 = \DFF_875.D ;
  assign g25720 = \DFF_388.D ;
  assign g25721 = \DFF_310.D ;
  assign g25722 = \DFF_651.D ;
  assign g25723 = \DFF_415.D ;
  assign g25724 = \DFF_636.D ;
  assign g25725 = \DFF_869.D ;
  assign g25726 = \DFF_438.D ;
  assign g25727 = \DFF_459.D ;
  assign g25728 = \DFF_85.D ;
  assign g25729 = \DFF_376.D ;
  assign g25730 = \DFF_396.D ;
  assign g25731 = \DFF_329.D ;
  assign g25732 = \DFF_572.D ;
  assign g25733 = \DFF_1306.D ;
  assign g25734 = \DFF_1332.D ;
  assign g25735 = \DFF_1198.D ;
  assign g25736 = \DFF_14.D ;
  assign g25737 = \DFF_1142.D ;
  assign g25738 = \DFF_1287.D ;
  assign g25739 = \DFF_344.D ;
  assign g25740 = \DFF_978.D ;
  assign g25741 = \DFF_138.D ;
  assign g25742 = \DFF_1316.D ;
  assign g25743 = \DFF_86.D ;
  assign g25744 = \DFF_838.D ;
  assign g25745 = \DFF_1048.D ;
  assign g25746 = \DFF_596.D ;
  assign g25747 = \DFF_400.D ;
  assign g25748 = \DFF_275.D ;
  assign g25749 = \DFF_287.D ;
  assign g2575 = \DFF_960.Q ;
  assign g25750 = \DFF_300.D ;
  assign g25751 = \DFF_3.D ;
  assign g25752 = \DFF_969.D ;
  assign g25753 = \DFF_1062.D ;
  assign g25754 = \DFF_1183.D ;
  assign g25755 = \DFF_266.D ;
  assign g25756 = \DFF_861.D ;
  assign g25757 = \DFF_371.D ;
  assign g25758 = \DFF_732.D ;
  assign g25759 = \DFF_1279.D ;
  assign g25760 = \DFF_907.D ;
  assign g25761 = \DFF_755.D ;
  assign g25762 = \DFF_1154.D ;
  assign g25763 = \DFF_332.D ;
  assign g25764 = \DFF_1055.D ;
  assign g25768 = \DFF_1336.Q ;
  assign g25771 = \DFF_489.Q ;
  assign g25775 = \DFF_1289.Q ;
  assign g25782 = \DFF_1282.Q ;
  assign g2579 = \DFF_890.Q ;
  assign g2583 = \DFF_1380.Q ;
  assign g25831 = \DFF_196.Q ;
  assign g25850 = \DFF_657.Q ;
  assign g25866 = \DFF_144.Q ;
  assign g2587 = \DFF_623.Q ;
  assign g25903 = \DFF_934.Q ;
  assign g2595 = \DFF_487.Q ;
  assign g25986 = \DFF_190.Q ;
  assign g2599 = \DFF_402.Q ;
  assign g26019 = \DFF_80.Q ;
  assign g26048 = \DFF_75.Q ;
  assign g2606 = \DFF_594.Q ;
  assign g26079 = \DFF_64.Q ;
  assign g26088 = \DFF_498.Q ;
  assign g2610 = \DFF_189.Q ;
  assign g26105 = g72;
  assign g26131 = g73;
  assign g26187 = g27831;
  assign g2619 = \DFF_562.Q ;
  assign g262 = \DFF_648.Q ;
  assign g2625 = \DFF_581.Q ;
  assign g26257 = \DFF_1340.Q ;
  assign g26260 = g23002;
  assign g26274 = \DFF_507.Q ;
  assign g26279 = \DFF_974.Q ;
  assign g26287 = \DFF_941.Q ;
  assign g2629 = \DFF_505.Q ;
  assign g26292 = \DFF_1067.Q ;
  assign g26294 = \DFF_1041.Q ;
  assign g26301 = \DFF_445.Q ;
  assign g26304 = \DFF_1270.Q ;
  assign g26312 = \DFF_1319.Q ;
  assign g26337 = g23190;
  assign g2638 = \DFF_1082.Q ;
  assign g2643 = \DFF_820.Q ;
  assign g2648 = \DFF_682.Q ;
  assign g26510 = \DFF_1425.Q ;
  assign g2652 = \DFF_568.Q ;
  assign g2657 = \DFF_45.Q ;
  assign g2661 = \DFF_1368.Q ;
  assign g2667 = \DFF_702.Q ;
  assign g2671 = \DFF_1071.Q ;
  assign g2675 = \DFF_933.Q ;
  assign g26802 = g26801;
  assign g2681 = \DFF_1267.Q ;
  assign g26811 = g23612;
  assign g26814 = g23652;
  assign g26817 = \DFF_828.Q ;
  assign g26818 = g28753;
  assign g26820 = g31521;
  assign g26824 = g23759;
  assign g26825 = \DFF_1078.Q ;
  assign g26829 = \DFF_69.Q ;
  assign g26833 = \DFF_236.Q ;
  assign g26834 = \DFF_1301.Q ;
  assign g26835 = \DFF_1033.Q ;
  assign g26838 = \DFF_608.Q ;
  assign g26839 = \DFF_706.Q ;
  assign g26840 = g113;
  assign g26842 = \DFF_1357.Q ;
  assign g26843 = \DFF_654.Q ;
  assign g26846 = \DFF_994.Q ;
  assign g26847 = \DFF_881.Q ;
  assign g26848 = \DFF_1151.Q ;
  assign g26849 = \DFF_1125.Q ;
  assign g2685 = \DFF_1140.Q ;
  assign g26850 = \DFF_1044.Q ;
  assign g26851 = \DFF_357.Q ;
  assign g26853 = \DFF_1301.Q ;
  assign g26854 = \DFF_1035.Q ;
  assign g26855 = \DFF_311.Q ;
  assign g26856 = g31656;
  assign g26858 = \DFF_1403.Q ;
  assign g26859 = \DFF_1059.Q ;
  assign g26860 = g31665;
  assign g26862 = \DFF_132.Q ;
  assign g26864 = \DFF_15.Q ;
  assign g26869 = g32185;
  assign g26870 = \DFF_125.Q ;
  assign g26880 = \DFF_760.D ;
  assign g26881 = \DFF_48.D ;
  assign g26882 = \DFF_1329.D ;
  assign g26883 = \DFF_753.D ;
  assign g26884 = \DFF_532.D ;
  assign g26885 = \DFF_1149.D ;
  assign g26886 = \DFF_756.D ;
  assign g26887 = \DFF_1269.D ;
  assign g26888 = \DFF_709.D ;
  assign g26889 = \DFF_1059.D ;
  assign g2689 = \DFF_1067.Q ;
  assign g26890 = \DFF_686.D ;
  assign g26891 = \DFF_240.D ;
  assign g26892 = \DFF_294.D ;
  assign g26893 = \DFF_654.D ;
  assign g26894 = \DFF_353.D ;
  assign g26895 = \DFF_728.D ;
  assign g26896 = \DFF_1044.D ;
  assign g26897 = \DFF_194.D ;
  assign g26898 = \DFF_524.D ;
  assign g26899 = \DFF_278.D ;
  assign g269 = \DFF_541.Q ;
  assign g26900 = \DFF_585.D ;
  assign g26901 = \DFF_382.D ;
  assign g26902 = \DFF_771.D ;
  assign g26903 = \DFF_496.D ;
  assign g26904 = \DFF_648.D ;
  assign g26905 = \DFF_362.D ;
  assign g26906 = \DFF_541.D ;
  assign g26907 = \DFF_346.D ;
  assign g26908 = \DFF_1164.D ;
  assign g26909 = \DFF_669.D ;
  assign g26910 = \DFF_799.D ;
  assign g26911 = \DFF_1099.D ;
  assign g26912 = \DFF_963.D ;
  assign g26913 = \DFF_1144.D ;
  assign g26914 = \DFF_1133.D ;
  assign g26915 = \DFF_296.D ;
  assign g26916 = \DFF_1046.D ;
  assign g26917 = \DFF_137.D ;
  assign g26918 = \DFF_1237.D ;
  assign g26919 = \DFF_1117.D ;
  assign g26920 = \DFF_211.D ;
  assign g26921 = \DFF_740.D ;
  assign g26922 = \DFF_403.D ;
  assign g26923 = \DFF_595.D ;
  assign g26924 = \DFF_774.D ;
  assign g26925 = \DFF_1159.D ;
  assign g26926 = \DFF_746.D ;
  assign g26927 = \DFF_1036.D ;
  assign g26928 = \DFF_1223.D ;
  assign g26929 = \DFF_946.D ;
  assign g26930 = \DFF_811.D ;
  assign g26931 = \DFF_763.D ;
  assign g26932 = \DFF_470.D ;
  assign g26933 = \DFF_534.D ;
  assign g26934 = \DFF_1104.D ;
  assign g26935 = \DFF_126.D ;
  assign g26936 = \DFF_448.D ;
  assign g26937 = \DFF_843.D ;
  assign g26938 = \DFF_860.D ;
  assign g26939 = \DFF_1230.D ;
  assign g26940 = \DFF_282.D ;
  assign g26941 = \DFF_527.D ;
  assign g26942 = \DFF_434.D ;
  assign g26943 = \DFF_1204.D ;
  assign g26944 = \DFF_1299.D ;
  assign g26945 = \DFF_1073.D ;
  assign g26946 = \DFF_234.D ;
  assign g26947 = \DFF_250.D ;
  assign g26948 = \DFF_1146.D ;
  assign g26949 = \DFF_482.D ;
  assign g26950 = \DFF_980.D ;
  assign g26951 = \DFF_159.D ;
  assign g26952 = \DFF_1221.D ;
  assign g26953 = \DFF_929.D ;
  assign g26954 = \DFF_1225.D ;
  assign g26955 = \DFF_348.D ;
  assign g26956 = \DFF_692.D ;
  assign g26957 = \DFF_490.D ;
  assign g26958 = \DFF_1411.D ;
  assign g26959 = \DFF_530.D ;
  assign g26960 = \DFF_184.D ;
  assign g26961 = \DFF_383.D ;
  assign g26962 = \DFF_911.D ;
  assign g26963 = \DFF_129.D ;
  assign g26964 = \DFF_1415.D ;
  assign g26965 = \DFF_1397.D ;
  assign g26966 = \DFF_121.D ;
  assign g26967 = \DFF_491.D ;
  assign g26968 = \DFF_808.D ;
  assign g26969 = \DFF_724.D ;
  assign g2697 = \DFF_1270.Q ;
  assign g26970 = \DFF_436.D ;
  assign g26971 = \DFF_79.D ;
  assign g27013 = \DFF_934.Q ;
  assign g2704 = \DFF_1319.Q ;
  assign g2710 = \DFF_611.Q ;
  assign g2711 = \DFF_1101.Q ;
  assign g2712 = \DFF_843.Q ;
  assign g27121 = \DFF_489.Q ;
  assign g2715 = \DFF_962.Q ;
  assign g2719 = \DFF_893.Q ;
  assign g2724 = \DFF_746.Q ;
  assign g2729 = \DFF_845.Q ;
  assign g27320 = g28753;
  assign g2735 = \DFF_1364.Q ;
  assign g2741 = \DFF_1080.Q ;
  assign g27438 = \DFF_1425.Q ;
  assign g2748 = \DFF_1020.Q ;
  assign g27511 = \DFF_748.D ;
  assign g27527 = g23002;
  assign g2756 = \DFF_428.Q ;
  assign g27576 = \DFF_1111.D ;
  assign g27585 = \DFF_1220.D ;
  assign g2759 = \DFF_951.Q ;
  assign g2763 = \DFF_451.Q ;
  assign g27662 = g31521;
  assign g2767 = \DFF_1036.Q ;
  assign g27675 = \DFF_1078.Q ;
  assign g27678 = \DFF_1242.Q ;
  assign g27686 = \DFF_948.Q ;
  assign g27698 = g25114;
  assign g27708 = \DFF_1301.Q ;
  assign g27709 = \DFF_1033.Q ;
  assign g2771 = \DFF_1.Q ;
  assign g27736 = \DFF_654.Q ;
  assign g27737 = g25167;
  assign g2775 = \DFF_1288.Q ;
  assign g27765 = \DFF_673.Q ;
  assign g27773 = \DFF_1044.Q ;
  assign g27774 = \DFF_357.Q ;
  assign g2779 = \DFF_1223.Q ;
  assign g278 = \DFF_128.Q ;
  assign g27822 = \DFF_767.Q ;
  assign g2783 = \DFF_319.Q ;
  assign g27832 = g27831;
  assign g2787 = \DFF_931.Q ;
  assign g27880 = \DFF_1059.Q ;
  assign g27881 = g31656;
  assign g2791 = \DFF_946.Q ;
  assign g27928 = \DFF_141.Q ;
  assign g27929 = g31665;
  assign g27930 = \DFF_132.Q ;
  assign g2795 = \DFF_811.Q ;
  assign g27956 = \DFF_125.Q ;
  assign g27961 = g25259;
  assign g27967 = \DFF_489.Q ;
  assign g2799 = \DFF_763.Q ;
  assign g27993 = g23612;
  assign g27996 = g23652;
  assign g27998 = \DFF_828.Q ;
  assign g28 = \DFF_790.Q ;
  assign g28009 = g23759;
  assign g2803 = \DFF_1112.Q ;
  assign g28043 = \DFF_802.D ;
  assign g28044 = \DFF_1145.D ;
  assign g28045 = \DFF_506.D ;
  assign g28046 = \DFF_1042.D ;
  assign g28047 = \DFF_238.D ;
  assign g28048 = \DFF_1390.D ;
  assign g28049 = \DFF_1126.D ;
  assign g28050 = \DFF_656.D ;
  assign g28051 = \DFF_135.D ;
  assign g28052 = \DFF_573.D ;
  assign g28053 = \DFF_1250.D ;
  assign g28054 = \DFF_1365.D ;
  assign g28055 = \DFF_710.D ;
  assign g28056 = \DFF_1241.D ;
  assign g28057 = \DFF_788.D ;
  assign g28058 = \DFF_901.D ;
  assign g28059 = \DFF_1153.D ;
  assign g28060 = \DFF_845.D ;
  assign g28061 = \DFF_1377.D ;
  assign g28062 = \DFF_57.D ;
  assign g28063 = \DFF_697.D ;
  assign g28064 = \DFF_513.D ;
  assign g28065 = \DFF_1239.D ;
  assign g28066 = \DFF_535.D ;
  assign g28067 = \DFF_1385.D ;
  assign g28068 = \DFF_548.D ;
  assign g28069 = \DFF_857.D ;
  assign g2807 = \DFF_284.Q ;
  assign g28070 = \DFF_154.D ;
  assign g28071 = \DFF_1139.D ;
  assign g28072 = \DFF_689.D ;
  assign g28073 = \DFF_1187.D ;
  assign g28074 = \DFF_1083.D ;
  assign g28075 = \DFF_1152.D ;
  assign g28076 = \DFF_114.D ;
  assign g28077 = \DFF_247.D ;
  assign g28078 = \DFF_330.D ;
  assign g28079 = \DFF_527.D ;
  assign g28080 = \DFF_434.D ;
  assign g28081 = \DFF_1204.D ;
  assign g28082 = \DFF_813.D ;
  assign g28083 = \DFF_747.D ;
  assign g28084 = \DFF_254.D ;
  assign g28085 = \DFF_647.D ;
  assign g28086 = \DFF_837.D ;
  assign g28087 = \DFF_782.D ;
  assign g28088 = \DFF_1206.D ;
  assign g28089 = \DFF_574.D ;
  assign g28090 = \DFF_229.D ;
  assign g28091 = \DFF_1116.D ;
  assign g28092 = \DFF_1124.D ;
  assign g28093 = \DFF_132.D ;
  assign g28094 = \DFF_1367.D ;
  assign g28095 = \DFF_787.D ;
  assign g28096 = \DFF_1205.D ;
  assign g28097 = \DFF_1333.D ;
  assign g28098 = \DFF_466.D ;
  assign g28099 = \DFF_249.D ;
  assign g28100 = \DFF_821.D ;
  assign g28101 = \DFF_879.D ;
  assign g28102 = \DFF_493.D ;
  assign g28103 = \DFF_975.D ;
  assign g28104 = \DFF_1113.D ;
  assign g28105 = \DFF_714.D ;
  assign g2811 = \DFF_470.Q ;
  assign g28142 = \DFF_1078.Q ;
  assign g28147 = \DFF_1111.D ;
  assign g2815 = \DFF_302.Q ;
  assign g28155 = \DFF_1301.Q ;
  assign g28156 = \DFF_1220.D ;
  assign g28157 = \DFF_1033.Q ;
  assign g28161 = \DFF_654.Q ;
  assign g28162 = \DFF_1044.Q ;
  assign g28163 = \DFF_357.Q ;
  assign g28166 = \DFF_1059.Q ;
  assign g28173 = \DFF_132.Q ;
  assign g28181 = \DFF_125.Q ;
  assign g28184 = \DFF_489.Q ;
  assign g28187 = \DFF_748.D ;
  assign g2819 = \DFF_233.Q ;
  assign g2823 = \DFF_534.Q ;
  assign g28262 = \DFF_934.Q ;
  assign g2827 = \DFF_1104.Q ;
  assign g283 = \DFF_802.Q ;
  assign g2831 = \DFF_865.Q ;
  assign g2834 = \DFF_576.Q ;
  assign g28367 = g23002;
  assign g2837 = \DFF_126.Q ;
  assign g2841 = \DFF_448.Q ;
  assign g2844 = \DFF_69.Q ;
  assign g2848 = \DFF_364.Q ;
  assign g2852 = \DFF_236.Q ;
  assign g2856 = \DFF_1182.Q ;
  assign g2860 = \DFF_608.Q ;
  assign g2864 = \DFF_781.Q ;
  assign g28652 = g33894;
  assign g2868 = \DFF_1035.Q ;
  assign g287 = \DFF_745.Q ;
  assign g28709 = g31521;
  assign g2873 = \DFF_881.Q ;
  assign g28752 = g23612;
  assign g28754 = g28753;
  assign g28779 = g23652;
  assign g2878 = \DFF_749.Q ;
  assign g28819 = \DFF_828.Q ;
  assign g2882 = \DFF_757.Q ;
  assign g2886 = \DFF_242.Q ;
  assign g2890 = \DFF_1178.Q ;
  assign g28917 = g23759;
  assign g2894 = \DFF_1357.Q ;
  assign g28954 = g26801;
  assign g2898 = \DFF_223.Q ;
  assign g29013 = g31656;
  assign g2902 = \DFF_531.Q ;
  assign g29041 = \DFF_1425.Q ;
  assign g29042 = g25114;
  assign g29043 = g31665;
  assign g2907 = \DFF_15.Q ;
  assign g291 = \DFF_106.Q ;
  assign g2912 = \DFF_1336.Q ;
  assign g29147 = g25167;
  assign g2917 = \DFF_899.Q ;
  assign g29185 = \DFF_141.Q ;
  assign g29194 = \DFF_748.D ;
  assign g29195 = g25259;
  assign g29209 = \DFF_748.D ;
  assign g29210 = \DFF_1425.Q ;
  assign g29211 = \DFF_654.Q ;
  assign g29212 = \DFF_1044.Q ;
  assign g29213 = \DFF_1078.Q ;
  assign g29214 = \DFF_1301.Q ;
  assign g29215 = \DFF_357.Q ;
  assign g29216 = \DFF_1059.Q ;
  assign g29217 = \DFF_125.Q ;
  assign g29218 = \DFF_934.Q ;
  assign g29219 = \DFF_1033.Q ;
  assign g2922 = \DFF_1289.Q ;
  assign g29220 = \DFF_132.Q ;
  assign g29221 = \DFF_489.Q ;
  assign g29222 = \DFF_1315.D ;
  assign g29223 = \DFF_47.D ;
  assign g29224 = \DFF_560.D ;
  assign g29225 = \DFF_902.D ;
  assign g29226 = \DFF_112.D ;
  assign g29227 = \DFF_1019.D ;
  assign g29228 = \DFF_876.D ;
  assign g29229 = \DFF_1251.D ;
  assign g29230 = \DFF_303.D ;
  assign g29231 = \DFF_1382.D ;
  assign g29232 = \DFF_921.D ;
  assign g29233 = \DFF_1274.D ;
  assign g29234 = \DFF_1290.D ;
  assign g29235 = \DFF_431.D ;
  assign g29236 = \DFF_169.D ;
  assign g29237 = \DFF_424.D ;
  assign g29238 = \DFF_720.D ;
  assign g29239 = \DFF_193.D ;
  assign g29240 = \DFF_1069.D ;
  assign g29241 = \DFF_1281.D ;
  assign g29242 = \DFF_1167.D ;
  assign g29243 = \DFF_977.D ;
  assign g29244 = \DFF_772.D ;
  assign g29245 = \DFF_777.D ;
  assign g29246 = \DFF_1310.D ;
  assign g29247 = \DFF_1129.D ;
  assign g29248 = \DFF_37.D ;
  assign g29249 = \DFF_1328.D ;
  assign g29250 = \DFF_406.D ;
  assign g29251 = \DFF_804.D ;
  assign g29252 = \DFF_989.D ;
  assign g29253 = \DFF_726.D ;
  assign g29254 = \DFF_1082.D ;
  assign g29255 = \DFF_568.D ;
  assign g29256 = \DFF_1364.D ;
  assign g29257 = \DFF_1372.D ;
  assign g29258 = \DFF_1409.D ;
  assign g29259 = \DFF_1358.D ;
  assign g29260 = \DFF_1302.D ;
  assign g29261 = \DFF_696.D ;
  assign g29262 = \DFF_839.D ;
  assign g29263 = \DFF_58.D ;
  assign g29264 = \DFF_688.D ;
  assign g29265 = \DFF_341.D ;
  assign g29266 = \DFF_778.D ;
  assign g29267 = \DFF_955.D ;
  assign g29268 = \DFF_559.D ;
  assign g29269 = \DFF_546.D ;
  assign g2927 = \DFF_852.Q ;
  assign g29270 = \DFF_742.D ;
  assign g29271 = \DFF_693.D ;
  assign g29272 = \DFF_441.D ;
  assign g29273 = \DFF_274.D ;
  assign g29274 = \DFF_1195.D ;
  assign g29275 = \DFF_411.D ;
  assign g29276 = \DFF_350.D ;
  assign g29277 = \DFF_1425.D ;
  assign g29278 = \DFF_439.D ;
  assign g29279 = \DFF_221.D ;
  assign g29280 = \DFF_1346.D ;
  assign g29281 = \DFF_1121.D ;
  assign g29282 = \DFF_145.D ;
  assign g29283 = \DFF_456.D ;
  assign g29284 = \DFF_1211.D ;
  assign g29285 = \DFF_826.D ;
  assign g29286 = \DFF_1066.D ;
  assign g29287 = \DFF_1021.D ;
  assign g29288 = \DFF_1215.D ;
  assign g29289 = \DFF_1079.D ;
  assign g29290 = \DFF_1018.D ;
  assign g29291 = \DFF_918.D ;
  assign g29292 = \DFF_463.D ;
  assign g29293 = \DFF_679.D ;
  assign g29294 = \DFF_632.D ;
  assign g29295 = \DFF_361.D ;
  assign g29296 = \DFF_213.D ;
  assign g29297 = \DFF_1138.D ;
  assign g29298 = \DFF_170.D ;
  assign g29299 = \DFF_1203.D ;
  assign g29300 = \DFF_897.D ;
  assign g29301 = \DFF_52.D ;
  assign g29302 = \DFF_1004.D ;
  assign g29303 = \DFF_136.D ;
  assign g29304 = \DFF_694.D ;
  assign g29305 = \DFF_987.D ;
  assign g29306 = \DFF_433.D ;
  assign g29307 = \DFF_716.D ;
  assign g29308 = \DFF_1278.D ;
  assign g29309 = \DFF_644.D ;
  assign g29317 = \DFF_1220.D ;
  assign g2932 = \DFF_349.Q ;
  assign g2936 = \DFF_1282.Q ;
  assign g29368 = g23612;
  assign g29371 = g23652;
  assign g29374 = \DFF_828.Q ;
  assign g29379 = g23759;
  assign g294 = \DFF_83.Q ;
  assign g2941 = \DFF_155.Q ;
  assign g2946 = \DFF_858.Q ;
  assign g29491 = g31665;
  assign g29498 = g31656;
  assign g2950 = \DFF_1151.Q ;
  assign g2955 = \DFF_95.Q ;
  assign g2960 = \DFF_311.Q ;
  assign g2965 = \DFF_733.Q ;
  assign g2970 = \DFF_1403.Q ;
  assign g29744 = g32185;
  assign g2975 = \DFF_399.Q ;
  assign g298 = \DFF_700.Q ;
  assign g2980 = \DFF_197.Q ;
  assign g29814 = \DFF_748.D ;
  assign g2984 = \DFF_413.Q ;
  assign g2988 = \DFF_706.Q ;
  assign g2994 = \DFF_1125.Q ;
  assign g2999 = \DFF_1245.Q ;
  assign g30012 = g31521;
  assign g3003 = \DFF_1381.Q ;
  assign g3004 = \DFF_976.Q ;
  assign g30072 = g25114;
  assign g301 = \DFF_708.Q ;
  assign g3010 = \DFF_205.Q ;
  assign g30105 = g25167;
  assign g30116 = g23002;
  assign g30155 = \DFF_141.Q ;
  assign g3017 = \DFF_8.Q ;
  assign g30182 = g25259;
  assign g3021 = \DFF_725.Q ;
  assign g30218 = g27831;
  assign g30237 = g33894;
  assign g3025 = \DFF_592.Q ;
  assign g3029 = \DFF_521.Q ;
  assign g30295 = g26801;
  assign g30301 = \DFF_1111.D ;
  assign g30322 = g32185;
  assign g30327 = g23002;
  assign g30329 = g23612;
  assign g30330 = g23652;
  assign g30331 = g23759;
  assign g30332 = \DFF_828.Q ;
  assign g30333 = \DFF_1060.D ;
  assign g30334 = \DFF_863.D ;
  assign g30335 = \DFF_175.D ;
  assign g30336 = \DFF_280.D ;
  assign g30337 = \DFF_421.D ;
  assign g30338 = \DFF_214.D ;
  assign g30339 = \DFF_563.D ;
  assign g3034 = \DFF_834.Q ;
  assign g30340 = \DFF_936.D ;
  assign g30341 = \DFF_277.D ;
  assign g30342 = \DFF_954.D ;
  assign g30343 = \DFF_577.D ;
  assign g30344 = \DFF_1148.D ;
  assign g30345 = \DFF_717.D ;
  assign g30346 = \DFF_1189.D ;
  assign g30347 = \DFF_614.D ;
  assign g30348 = \DFF_164.D ;
  assign g30349 = \DFF_583.D ;
  assign g30350 = \DFF_446.D ;
  assign g30351 = \DFF_1226.D ;
  assign g30352 = \DFF_1418.D ;
  assign g30353 = \DFF_984.D ;
  assign g30354 = \DFF_1051.D ;
  assign g30355 = \DFF_1243.D ;
  assign g30356 = \DFF_882.D ;
  assign g30357 = \DFF_1163.D ;
  assign g30358 = \DFF_1202.D ;
  assign g30359 = \DFF_1216.D ;
  assign g30360 = \DFF_42.D ;
  assign g30361 = \DFF_1369.D ;
  assign g30362 = \DFF_520.D ;
  assign g30363 = \DFF_862.D ;
  assign g30364 = \DFF_964.D ;
  assign g30365 = \DFF_888.D ;
  assign g30366 = \DFF_264.D ;
  assign g30367 = \DFF_1213.D ;
  assign g30368 = \DFF_570.D ;
  assign g30369 = \DFF_301.D ;
  assign g30370 = \DFF_232.D ;
  assign g30371 = \DFF_558.D ;
  assign g30372 = \DFF_1031.D ;
  assign g30373 = \DFF_1240.D ;
  assign g30374 = \DFF_928.D ;
  assign g30375 = \DFF_571.D ;
  assign g30376 = \DFF_1276.D ;
  assign g30377 = \DFF_499.D ;
  assign g30378 = \DFF_425.D ;
  assign g30379 = \DFF_818.D ;
  assign g30380 = \DFF_1395.D ;
  assign g30381 = \DFF_6.D ;
  assign g30382 = \DFF_825.D ;
  assign g30383 = \DFF_487.D ;
  assign g30384 = \DFF_45.D ;
  assign g30385 = \DFF_1368.D ;
  assign g30386 = \DFF_1267.D ;
  assign g30387 = \DFF_1140.D ;
  assign g30388 = \DFF_1080.D ;
  assign g30389 = \DFF_1033.D ;
  assign g30390 = \DFF_125.D ;
  assign g30391 = \DFF_865.D ;
  assign g30392 = \DFF_576.D ;
  assign g30393 = \DFF_35.D ;
  assign g30394 = \DFF_1378.D ;
  assign g30395 = \DFF_1386.D ;
  assign g30396 = \DFF_1197.D ;
  assign g30397 = \DFF_1208.D ;
  assign g30398 = \DFF_1218.D ;
  assign g30399 = \DFF_1166.D ;
  assign g3040 = \DFF_176.Q ;
  assign g30400 = \DFF_1401.D ;
  assign g30401 = \DFF_640.D ;
  assign g30402 = \DFF_370.D ;
  assign g30403 = \DFF_225.D ;
  assign g30404 = \DFF_134.D ;
  assign g30405 = \DFF_9.D ;
  assign g30406 = \DFF_670.D ;
  assign g30407 = \DFF_1410.D ;
  assign g30408 = \DFF_1280.D ;
  assign g30409 = \DFF_1210.D ;
  assign g30410 = \DFF_1263.D ;
  assign g30411 = \DFF_645.D ;
  assign g30412 = \DFF_1351.D ;
  assign g30413 = \DFF_729.D ;
  assign g30414 = \DFF_120.D ;
  assign g30415 = \DFF_707.D ;
  assign g30416 = \DFF_12.D ;
  assign g30417 = \DFF_1259.D ;
  assign g30418 = \DFF_309.D ;
  assign g30419 = \DFF_227.D ;
  assign g30420 = \DFF_108.D ;
  assign g30421 = \DFF_321.D ;
  assign g30422 = \DFF_628.D ;
  assign g30423 = \DFF_633.D ;
  assign g30424 = \DFF_105.D ;
  assign g30425 = \DFF_1052.D ;
  assign g30426 = \DFF_1244.D ;
  assign g30427 = \DFF_72.D ;
  assign g30428 = \DFF_626.D ;
  assign g30429 = \DFF_102.D ;
  assign g30430 = \DFF_1177.D ;
  assign g30431 = \DFF_982.D ;
  assign g30432 = \DFF_19.D ;
  assign g30433 = \DFF_738.D ;
  assign g30434 = \DFF_1356.D ;
  assign g30435 = \DFF_784.D ;
  assign g30436 = \DFF_340.D ;
  assign g30437 = \DFF_1350.D ;
  assign g30438 = \DFF_312.D ;
  assign g30439 = \DFF_91.D ;
  assign g30440 = \DFF_479.D ;
  assign g30441 = \DFF_1128.D ;
  assign g30442 = \DFF_986.D ;
  assign g30443 = \DFF_917.D ;
  assign g30444 = \DFF_257.D ;
  assign g30445 = \DFF_868.D ;
  assign g30446 = \DFF_1160.D ;
  assign g30447 = \DFF_1013.D ;
  assign g30448 = \DFF_947.D ;
  assign g30449 = \DFF_1317.D ;
  assign g3045 = \DFF_618.Q ;
  assign g30450 = \DFF_550.D ;
  assign g30451 = \DFF_414.D ;
  assign g30452 = \DFF_590.D ;
  assign g30453 = \DFF_156.D ;
  assign g30454 = \DFF_1264.D ;
  assign g30455 = \DFF_253.D ;
  assign g30456 = \DFF_551.D ;
  assign g30457 = \DFF_116.D ;
  assign g30458 = \DFF_1399.D ;
  assign g30459 = \DFF_407.D ;
  assign g30460 = \DFF_638.D ;
  assign g30461 = \DFF_1325.D ;
  assign g30462 = \DFF_390.D ;
  assign g30463 = \DFF_602.D ;
  assign g30464 = \DFF_923.D ;
  assign g30465 = \DFF_1186.D ;
  assign g30466 = \DFF_13.D ;
  assign g30467 = \DFF_983.D ;
  assign g30468 = \DFF_773.D ;
  assign g30469 = \DFF_950.D ;
  assign g30470 = \DFF_1212.D ;
  assign g30471 = \DFF_1095.D ;
  assign g30472 = \DFF_659.D ;
  assign g30473 = \DFF_1406.D ;
  assign g30474 = \DFF_187.D ;
  assign g30475 = \DFF_497.D ;
  assign g30476 = \DFF_100.D ;
  assign g30477 = \DFF_1040.D ;
  assign g30478 = \DFF_750.D ;
  assign g30479 = \DFF_1363.D ;
  assign g30480 = \DFF_244.D ;
  assign g30481 = \DFF_333.D ;
  assign g30482 = \DFF_938.D ;
  assign g30483 = \DFF_151.D ;
  assign g30484 = \DFF_1007.D ;
  assign g30485 = \DFF_627.D ;
  assign g30486 = \DFF_476.D ;
  assign g30487 = \DFF_392.D ;
  assign g30488 = \DFF_895.D ;
  assign g30489 = \DFF_51.D ;
  assign g30490 = \DFF_71.D ;
  assign g30491 = \DFF_1355.D ;
  assign g30492 = \DFF_1297.D ;
  assign g30493 = \DFF_884.D ;
  assign g30494 = \DFF_44.D ;
  assign g30495 = \DFF_219.D ;
  assign g30496 = \DFF_55.D ;
  assign g30497 = \DFF_307.D ;
  assign g30498 = \DFF_84.D ;
  assign g30499 = \DFF_172.D ;
  assign g305 = \DFF_760.Q ;
  assign g3050 = \DFF_259.Q ;
  assign g30500 = \DFF_1423.D ;
  assign g30501 = \DFF_734.D ;
  assign g30502 = \DFF_267.D ;
  assign g30503 = \DFF_1291.D ;
  assign g30504 = \DFF_241.D ;
  assign g30505 = \DFF_17.D ;
  assign g30506 = \DFF_398.D ;
  assign g30507 = \DFF_1058.D ;
  assign g30508 = \DFF_920.D ;
  assign g30509 = \DFF_854.D ;
  assign g30510 = \DFF_192.D ;
  assign g30511 = \DFF_815.D ;
  assign g30512 = \DFF_1085.D ;
  assign g30513 = \DFF_949.D ;
  assign g30514 = \DFF_877.D ;
  assign g30515 = \DFF_1255.D ;
  assign g30516 = \DFF_471.D ;
  assign g30517 = \DFF_336.D ;
  assign g30518 = \DFF_526.D ;
  assign g30519 = \DFF_93.D ;
  assign g30520 = \DFF_1201.D ;
  assign g30521 = \DFF_183.D ;
  assign g30522 = \DFF_925.D ;
  assign g30523 = \DFF_579.D ;
  assign g30524 = \DFF_494.D ;
  assign g30525 = \DFF_945.D ;
  assign g30526 = \DFF_158.D ;
  assign g30527 = \DFF_1011.D ;
  assign g30528 = \DFF_179.D ;
  assign g30529 = \DFF_634.D ;
  assign g30530 = \DFF_483.D ;
  assign g30531 = \DFF_397.D ;
  assign g30532 = \DFF_904.D ;
  assign g30533 = \DFF_59.D ;
  assign g30534 = \DFF_82.D ;
  assign g30535 = \DFF_1366.D ;
  assign g30536 = \DFF_1307.D ;
  assign g30537 = \DFF_1123.D ;
  assign g30538 = \DFF_298.D ;
  assign g30539 = \DFF_337.D ;
  assign g30540 = \DFF_314.D ;
  assign g30541 = \DFF_92.D ;
  assign g30542 = \DFF_484.D ;
  assign g30543 = \DFF_410.D ;
  assign g30544 = \DFF_1174.D ;
  assign g30545 = \DFF_1032.D ;
  assign g30546 = \DFF_610.D ;
  assign g30547 = \DFF_1169.D ;
  assign g30548 = \DFF_957.D ;
  assign g30549 = \DFF_730.D ;
  assign g30550 = \DFF_1294.D ;
  assign g30551 = \DFF_588.D ;
  assign g30552 = \DFF_419.D ;
  assign g30553 = \DFF_345.D ;
  assign g30554 = \DFF_1120.D ;
  assign g30555 = \DFF_291.D ;
  assign g30556 = \DFF_617.D ;
  assign g30557 = \DFF_464.D ;
  assign g30558 = \DFF_378.D ;
  assign g30559 = \DFF_779.D ;
  assign g30560 = \DFF_967.D ;
  assign g30561 = \DFF_1175.D ;
  assign g30562 = \DFF_1024.D ;
  assign g30563 = \DFF_1348.D ;
  assign g30565 = \DFF_1111.D ;
  assign g3057 = \DFF_57.Q ;
  assign g30591 = \DFF_1220.D ;
  assign g3061 = \DFF_1377.Q ;
  assign g30610 = g25114;
  assign g3065 = \DFF_1249.Q ;
  assign g3068 = \DFF_1318.Q ;
  assign g3072 = \DFF_827.Q ;
  assign g30729 = g25167;
  assign g3080 = \DFF_775.Q ;
  assign g3085 = \DFF_1156.Q ;
  assign g3089 = \DFF_1076.Q ;
  assign g30917 = \DFF_141.Q ;
  assign g3092 = \DFF_317.Q ;
  assign g30928 = g25259;
  assign g30931 = g32185;
  assign g3096 = \DFF_1256.Q ;
  assign g31 = \DFF_512.Q ;
  assign g3100 = \DFF_166.Q ;
  assign g3103 = \DFF_817.Q ;
  assign g3106 = \DFF_1372.Q ;
  assign g311 = \DFF_48.Q ;
  assign g3111 = \DFF_124.Q ;
  assign g3115 = \DFF_1409.Q ;
  assign g3119 = \DFF_1342.Q ;
  assign g3125 = \DFF_1358.Q ;
  assign g3129 = \DFF_1302.Q ;
  assign g3133 = \DFF_696.Q ;
  assign g3139 = \DFF_356.Q ;
  assign g3143 = \DFF_222.Q ;
  assign g3147 = \DFF_839.Q ;
  assign g3151 = \DFF_196.Q ;
  assign g31522 = g31521;
  assign g3155 = \DFF_35.Q ;
  assign g31578 = g33894;
  assign g316 = \DFF_753.Q ;
  assign g3161 = \DFF_803.Q ;
  assign g31655 = g26801;
  assign g31657 = g31656;
  assign g31666 = g31665;
  assign g31667 = g28753;
  assign g3167 = \DFF_54.Q ;
  assign g3171 = \DFF_522.Q ;
  assign g3179 = \DFF_271.Q ;
  assign g31791 = g27831;
  assign g31860 = g25114;
  assign g31861 = \DFF_141.Q ;
  assign g31862 = g25259;
  assign g31863 = g25167;
  assign g31864 = \DFF_1339.D ;
  assign g31865 = \DFF_745.D ;
  assign g31866 = \DFF_1235.D ;
  assign g31867 = \DFF_28.D ;
  assign g31868 = \DFF_859.D ;
  assign g31869 = \DFF_70.D ;
  assign g3187 = \DFF_1378.Q ;
  assign g31870 = \DFF_454.D ;
  assign g31871 = \DFF_1227.D ;
  assign g31872 = \DFF_1020.D ;
  assign g31873 = \DFF_976.D ;
  assign g31874 = \DFF_592.D ;
  assign g31875 = \DFF_521.D ;
  assign g31876 = \DFF_834.D ;
  assign g31877 = \DFF_8.D ;
  assign g31878 = \DFF_176.D ;
  assign g31879 = \DFF_725.D ;
  assign g31880 = \DFF_36.D ;
  assign g31881 = \DFF_1170.D ;
  assign g31882 = \DFF_140.D ;
  assign g31883 = \DFF_586.D ;
  assign g31884 = \DFF_762.D ;
  assign g31885 = \DFF_1388.D ;
  assign g31886 = \DFF_217.D ;
  assign g31887 = \DFF_516.D ;
  assign g31888 = \DFF_1309.D ;
  assign g31889 = \DFF_1077.D ;
  assign g31890 = \DFF_335.D ;
  assign g31891 = \DFF_475.D ;
  assign g31892 = \DFF_381.D ;
  assign g31893 = \DFF_741.D ;
  assign g31894 = \DFF_351.D ;
  assign g31895 = \DFF_1272.D ;
  assign g31896 = \DFF_624.D ;
  assign g31897 = \DFF_1022.D ;
  assign g31898 = \DFF_1341.D ;
  assign g31899 = \DFF_386.D ;
  assign g319 = \DFF_1329.Q ;
  assign g31900 = \DFF_690.D ;
  assign g31901 = \DFF_1327.D ;
  assign g31902 = \DFF_432.D ;
  assign g31903 = \DFF_502.D ;
  assign g31904 = \DFF_1192.D ;
  assign g31905 = \DFF_191.D ;
  assign g31906 = \DFF_665.D ;
  assign g31907 = \DFF_518.D ;
  assign g31908 = \DFF_823.D ;
  assign g31909 = \DFF_557.D ;
  assign g3191 = \DFF_1386.Q ;
  assign g31910 = \DFF_639.D ;
  assign g31911 = \DFF_1132.D ;
  assign g31912 = \DFF_426.D ;
  assign g31913 = \DFF_1246.D ;
  assign g31914 = \DFF_1015.D ;
  assign g31915 = \DFF_260.D ;
  assign g31916 = \DFF_394.D ;
  assign g31917 = \DFF_308.D ;
  assign g31918 = \DFF_676.D ;
  assign g31919 = \DFF_851.D ;
  assign g31920 = \DFF_40.D ;
  assign g31921 = \DFF_712.D ;
  assign g31922 = \DFF_1321.D ;
  assign g31923 = \DFF_122.D ;
  assign g31924 = \DFF_97.D ;
  assign g31925 = \DFF_49.D ;
  assign g31926 = \DFF_230.D ;
  assign g31927 = \DFF_850.D ;
  assign g31928 = \DFF_1105.D ;
  assign g31929 = \DFF_940.D ;
  assign g31930 = \DFF_1056.D ;
  assign g31931 = \DFF_1147.D ;
  assign g31932 = \DFF_915.D ;
  assign g3195 = \DFF_1263.Q ;
  assign g3199 = \DFF_1197.Q ;
  assign g32021 = \DFF_1111.D ;
  assign g32024 = \DFF_1220.D ;
  assign g32027 = g26801;
  assign g3203 = \DFF_645.Q ;
  assign g3207 = \DFF_1208.Q ;
  assign g3211 = \DFF_1351.Q ;
  assign g3215 = \DFF_1218.Q ;
  assign g32186 = g32185;
  assign g3219 = \DFF_1166.Q ;
  assign g3223 = \DFF_1401.Q ;
  assign g3227 = \DFF_640.Q ;
  assign g3231 = \DFF_370.Q ;
  assign g3235 = \DFF_225.Q ;
  assign g32363 = g33894;
  assign g32381 = g27831;
  assign g3239 = \DFF_134.Q ;
  assign g324 = \DFF_1269.Q ;
  assign g32407 = g28753;
  assign g32429 = 1'b1;
  assign g3243 = \DFF_9.Q ;
  assign g32454 = 1'b1;
  assign g3247 = \DFF_670.Q ;
  assign g3251 = \DFF_1410.Q ;
  assign g3255 = \DFF_1280.Q ;
  assign g3259 = \DFF_1210.Q ;
  assign g3263 = \DFF_729.Q ;
  assign g3267 = \DFF_1293.Q ;
  assign g3274 = \DFF_1354.Q ;
  assign g3281 = \DFF_529.Q ;
  assign g3288 = \DFF_443.Q ;
  assign g329 = \DFF_1149.Q ;
  assign g32975 = g26801;
  assign g32976 = \DFF_582.D ;
  assign g32977 = \DFF_106.D ;
  assign g32978 = \DFF_162.D ;
  assign g32979 = \DFF_328.D ;
  assign g3298 = \DFF_1155.Q ;
  assign g32980 = \DFF_719.D ;
  assign g32981 = \DFF_149.D ;
  assign g32982 = \DFF_758.D ;
  assign g32983 = \DFF_368.D ;
  assign g32984 = \DFF_913.D ;
  assign g32985 = \DFF_754.D ;
  assign g32986 = \DFF_316.D ;
  assign g32987 = \DFF_1064.D ;
  assign g32988 = \DFF_1344.D ;
  assign g32989 = \DFF_794.D ;
  assign g32990 = \DFF_342.D ;
  assign g32991 = \DFF_552.D ;
  assign g32992 = \DFF_1037.D ;
  assign g32993 = \DFF_1375.D ;
  assign g32994 = \DFF_153.D ;
  assign g32995 = \DFF_705.D ;
  assign g32996 = \DFF_174.D ;
  assign g32997 = \DFF_103.D ;
  assign g32998 = \DFF_1063.D ;
  assign g32999 = \DFF_1070.D ;
  assign g33000 = \DFF_1236.D ;
  assign g33001 = \DFF_1295.D ;
  assign g33002 = \DFF_1093.D ;
  assign g33003 = \DFF_993.D ;
  assign g33004 = \DFF_889.D ;
  assign g33005 = \DFF_1091.D ;
  assign g33006 = \DFF_462.D ;
  assign g33007 = \DFF_387.D ;
  assign g33008 = \DFF_297.D ;
  assign g33009 = \DFF_681.D ;
  assign g33010 = \DFF_1337.D ;
  assign g33011 = \DFF_1331.D ;
  assign g33012 = \DFF_793.D ;
  assign g33013 = \DFF_148.D ;
  assign g33014 = \DFF_1028.D ;
  assign g33015 = \DFF_623.D ;
  assign g33016 = \DFF_189.D ;
  assign g33017 = \DFF_562.D ;
  assign g33018 = \DFF_581.D ;
  assign g33019 = \DFF_428.D ;
  assign g33020 = \DFF_618.D ;
  assign g33021 = \DFF_803.D ;
  assign g33022 = \DFF_54.D ;
  assign g33023 = \DFF_522.D ;
  assign g33024 = \DFF_271.D ;
  assign g33025 = \DFF_703.D ;
  assign g33026 = \DFF_27.D ;
  assign g33027 = \DFF_245.D ;
  assign g33028 = \DFF_1408.D ;
  assign g33029 = \DFF_199.D ;
  assign g3303 = \DFF_819.Q ;
  assign g33030 = \DFF_1334.D ;
  assign g33031 = \DFF_776.D ;
  assign g33032 = \DFF_473.D ;
  assign g33033 = \DFF_467.D ;
  assign g33034 = \DFF_587.D ;
  assign g33035 = \DFF_508.D ;
  assign g33036 = \DFF_268.D ;
  assign g33037 = \DFF_352.D ;
  assign g33038 = \DFF_744.D ;
  assign g33039 = \DFF_384.D ;
  assign g33040 = \DFF_1296.D ;
  assign g33041 = \DFF_1330.D ;
  assign g33042 = \DFF_226.D ;
  assign g33043 = \DFF_56.D ;
  assign g33044 = \DFF_1349.D ;
  assign g33045 = \DFF_816.D ;
  assign g33046 = \DFF_0.D ;
  assign g33047 = \DFF_1304.D ;
  assign g33048 = \DFF_1098.D ;
  assign g33049 = \DFF_68.D ;
  assign g33050 = \DFF_598.D ;
  assign g33051 = \DFF_1238.D ;
  assign g33052 = \DFF_958.D ;
  assign g33053 = \DFF_289.D ;
  assign g33054 = \DFF_910.D ;
  assign g33055 = \DFF_575.D ;
  assign g33056 = \DFF_1271.D ;
  assign g33057 = \DFF_723.D ;
  assign g33058 = \DFF_393.D ;
  assign g33059 = \DFF_385.D ;
  assign g33060 = \DFF_519.D ;
  assign g33061 = \DFF_998.D ;
  assign g33062 = \DFF_653.D ;
  assign g33063 = \DFF_104.D ;
  assign g33064 = \DFF_20.D ;
  assign g33065 = \DFF_916.D ;
  assign g33066 = \DFF_1257.D ;
  assign g33067 = \DFF_584.D ;
  assign g33068 = \DFF_1273.D ;
  assign g33069 = \DFF_1150.D ;
  assign g33070 = \DFF_1068.D ;
  assign g33076 = g33874;
  assign g33079 = \DFF_1220.D ;
  assign g33080 = \DFF_1220.D ;
  assign g3310 = \DFF_1038.Q ;
  assign g33120 = g27831;
  assign g33149 = \DFF_512.D ;
  assign g33164 = \DFF_790.D ;
  assign g3317 = \DFF_856.Q ;
  assign g33176 = \DFF_1229.D ;
  assign g33187 = \DFF_355.D ;
  assign g33197 = \DFF_547.D ;
  assign g33204 = \DFF_761.D ;
  assign g3321 = \DFF_76.Q ;
  assign g33212 = \DFF_1222.D ;
  assign g33219 = \DFF_619.D ;
  assign g33228 = g33894;
  assign g3325 = \DFF_1359.Q ;
  assign g33283 = g33659;
  assign g3329 = \DFF_1303.Q ;
  assign g333 = \DFF_532.Q ;
  assign g33318 = g33636;
  assign g33323 = g33935;
  assign g3333 = \DFF_697.Q ;
  assign g33354 = g31521;
  assign g33377 = g28753;
  assign g3338 = \DFF_538.Q ;
  assign g33388 = g31656;
  assign g33391 = g31665;
  assign g3343 = \DFF_224.Q ;
  assign g33435 = \DFF_1111.D ;
  assign g33436 = \DFF_1111.D ;
  assign g3347 = \DFF_840.Q ;
  assign g3352 = \DFF_1347.Q ;
  assign g33533 = g27831;
  assign g33534 = \DFF_409.D ;
  assign g33535 = \DFF_83.D ;
  assign g33536 = \DFF_708.D ;
  assign g33537 = \DFF_258.D ;
  assign g33538 = \DFF_1090.D ;
  assign g33539 = \DFF_157.D ;
  assign g33540 = \DFF_867.D ;
  assign g33541 = \DFF_131.D ;
  assign g33542 = \DFF_1109.D ;
  assign g33543 = \DFF_1419.D ;
  assign g33544 = \DFF_1054.D ;
  assign g33545 = \DFF_1127.D ;
  assign g33546 = \DFF_646.D ;
  assign g33547 = \DFF_1266.D ;
  assign g33548 = \DFF_212.D ;
  assign g33549 = \DFF_1277.D ;
  assign g3355 = \DFF_36.Q ;
  assign g33550 = \DFF_33.D ;
  assign g33551 = \DFF_1089.D ;
  assign g33552 = \DFF_272.D ;
  assign g33553 = \DFF_500.D ;
  assign g33554 = \DFF_18.D ;
  assign g33555 = \DFF_1114.D ;
  assign g33556 = \DFF_649.D ;
  assign g33557 = \DFF_814.D ;
  assign g33558 = \DFF_1075.D ;
  assign g33559 = \DFF_567.D ;
  assign g33560 = \DFF_111.D ;
  assign g33561 = \DFF_759.D ;
  assign g33562 = \DFF_620.D ;
  assign g33563 = \DFF_832.D ;
  assign g33564 = \DFF_912.D ;
  assign g33565 = \DFF_1179.D ;
  assign g33566 = \DFF_1184.D ;
  assign g33567 = \DFF_1009.D ;
  assign g33568 = \DFF_1413.D ;
  assign g33569 = \DFF_671.D ;
  assign g33570 = \DFF_996.D ;
  assign g33571 = \DFF_77.D ;
  assign g33572 = \DFF_1086.D ;
  assign g33573 = \DFF_322.D ;
  assign g33574 = \DFF_1261.D ;
  assign g33575 = \DFF_472.D ;
  assign g33576 = \DFF_769.D ;
  assign g33577 = \DFF_1141.D ;
  assign g33578 = \DFF_1047.D ;
  assign g33579 = \DFF_1050.D ;
  assign g33580 = \DFF_903.D ;
  assign g33581 = \DFF_841.D ;
  assign g33582 = \DFF_835.D ;
  assign g33583 = \DFF_658.D ;
  assign g33584 = \DFF_209.D ;
  assign g33585 = \DFF_1010.D ;
  assign g33586 = \DFF_1233.D ;
  assign g33587 = \DFF_637.D ;
  assign g33588 = \DFF_216.D ;
  assign g33589 = \DFF_444.D ;
  assign g33590 = \DFF_1034.D ;
  assign g33591 = \DFF_943.D ;
  assign g33592 = \DFF_1143.D ;
  assign g33593 = \DFF_265.D ;
  assign g33594 = \DFF_886.D ;
  assign g33595 = \DFF_442.D ;
  assign g33596 = \DFF_1268.D ;
  assign g33597 = \DFF_488.D ;
  assign g33598 = \DFF_768.D ;
  assign g33599 = \DFF_1254.D ;
  assign g336 = \DFF_756.Q ;
  assign g33600 = \DFF_713.D ;
  assign g33601 = \DFF_402.D ;
  assign g33602 = \DFF_505.D ;
  assign g33603 = \DFF_682.D ;
  assign g33604 = \DFF_702.D ;
  assign g33605 = \DFF_1071.D ;
  assign g33606 = \DFF_933.D ;
  assign g33607 = \DFF_594.D ;
  assign g33608 = \DFF_951.D ;
  assign g33609 = \DFF_1347.D ;
  assign g3361 = \DFF_805.Q ;
  assign g33610 = \DFF_443.D ;
  assign g33611 = \DFF_1312.D ;
  assign g33612 = \DFF_536.D ;
  assign g33613 = \DFF_286.D ;
  assign g33614 = \DFF_517.D ;
  assign g33615 = \DFF_201.D ;
  assign g33616 = \DFF_1345.D ;
  assign g33617 = \DFF_1362.D ;
  assign g33618 = \DFF_846.D ;
  assign g33619 = \DFF_449.D ;
  assign g33620 = \DFF_1252.D ;
  assign g33621 = \DFF_1283.D ;
  assign g33622 = \DFF_833.D ;
  assign g33623 = \DFF_429.D ;
  assign g33624 = \DFF_139.D ;
  assign g33625 = \DFF_118.D ;
  assign g33626 = \DFF_952.D ;
  assign g33627 = \DFF_878.D ;
  assign g33628 = g34221;
  assign g33631 = \DFF_619.D ;
  assign g33637 = g33636;
  assign g33638 = g31656;
  assign g33641 = \DFF_1222.D ;
  assign g33645 = g31665;
  assign g33648 = \DFF_761.D ;
  assign g33653 = \DFF_547.D ;
  assign g33660 = g33659;
  assign g33661 = \DFF_355.D ;
  assign g33665 = \DFF_1229.D ;
  assign g33670 = \DFF_790.D ;
  assign g3368 = \DFF_762.Q ;
  assign g33682 = \DFF_355.D ;
  assign g33688 = \DFF_355.D ;
  assign g33691 = \DFF_619.D ;
  assign g33696 = g28753;
  assign g33698 = \DFF_1222.D ;
  assign g33702 = \DFF_619.D ;
  assign g33705 = \DFF_761.D ;
  assign g33708 = \DFF_1222.D ;
  assign g33712 = \DFF_547.D ;
  assign g33713 = \DFF_761.D ;
  assign g33716 = \DFF_547.D ;
  assign g3372 = \DFF_217.Q ;
  assign g33726 = \DFF_790.D ;
  assign g33729 = \DFF_512.D ;
  assign g33736 = \DFF_355.D ;
  assign g33744 = \DFF_1229.D ;
  assign g33750 = \DFF_790.D ;
  assign g33755 = \DFF_512.D ;
  assign g3376 = \DFF_1170.Q ;
  assign g33761 = \DFF_619.D ;
  assign g33766 = \DFF_1222.D ;
  assign g33772 = \DFF_761.D ;
  assign g33778 = \DFF_547.D ;
  assign g33791 = g34201;
  assign g3380 = \DFF_140.Q ;
  assign g33800 = \DFF_761.D ;
  assign g33804 = g32185;
  assign g33806 = \DFF_1222.D ;
  assign g33813 = \DFF_619.D ;
  assign g33827 = \DFF_512.D ;
  assign g33839 = \DFF_790.D ;
  assign g33845 = \DFF_1229.D ;
  assign g3385 = \DFF_586.Q ;
  assign g33850 = \DFF_790.D ;
  assign g33875 = g33874;
  assign g33895 = g33894;
  assign g3391 = \DFF_1388.Q ;
  assign g33912 = \DFF_547.D ;
  assign g33916 = \DFF_761.D ;
  assign g33917 = \DFF_1222.D ;
  assign g33918 = \DFF_619.D ;
  assign g33920 = \DFF_547.D ;
  assign g33923 = g31521;
  assign g33926 = \DFF_1229.D ;
  assign g33928 = \DFF_790.D ;
  assign g33929 = \DFF_1229.D ;
  assign g33931 = \DFF_512.D ;
  assign g33932 = \DFF_790.D ;
  assign g33934 = \DFF_512.D ;
  assign g33936 = g33935;
  assign g33937 = \DFF_512.D ;
  assign g33945 = 1'b1;
  assign g33946 = 1'b1;
  assign g33947 = 1'b1;
  assign g33948 = 1'b1;
  assign g33949 = 1'b1;
  assign g33950 = 1'b1;
  assign g33959 = g28753;
  assign g3396 = \DFF_703.Q ;
  assign g33960 = \DFF_318.D ;
  assign g33961 = \DFF_700.D ;
  assign g33962 = \DFF_357.D ;
  assign g33963 = \DFF_143.D ;
  assign g33964 = \DFF_874.D ;
  assign g33965 = \DFF_74.D ;
  assign g33966 = \DFF_32.D ;
  assign g33967 = \DFF_564.D ;
  assign g33968 = \DFF_1180.D ;
  assign g33969 = \DFF_735.D ;
  assign g33970 = \DFF_864.D ;
  assign g33971 = \DFF_293.D ;
  assign g33972 = \DFF_246.D ;
  assign g33973 = \DFF_41.D ;
  assign g33974 = \DFF_16.D ;
  assign g33975 = \DFF_306.D ;
  assign g33976 = \DFF_173.D ;
  assign g33977 = \DFF_1137.D ;
  assign g33978 = \DFF_435.D ;
  assign g33979 = \DFF_1258.D ;
  assign g33980 = \DFF_973.D ;
  assign g33981 = \DFF_1422.D ;
  assign g33982 = \DFF_2.D ;
  assign g33983 = \DFF_968.D ;
  assign g33984 = \DFF_504.D ;
  assign g33985 = \DFF_455.D ;
  assign g33986 = \DFF_1172.D ;
  assign g33987 = \DFF_1394.D ;
  assign g33988 = \DFF_924.D ;
  assign g33989 = \DFF_465.D ;
  assign g33990 = \DFF_641.D ;
  assign g33991 = \DFF_809.D ;
  assign g33992 = \DFF_1376.D ;
  assign g33993 = \DFF_255.D ;
  assign g33994 = \DFF_1231.D ;
  assign g33995 = \DFF_1030.D ;
  assign g33996 = \DFF_1026.D ;
  assign g33997 = \DFF_204.D ;
  assign g33998 = \DFF_1135.D ;
  assign g33999 = \DFF_374.D ;
  assign g34 = \DFF_1074.Q ;
  assign g34000 = \DFF_1096.D ;
  assign g34001 = \DFF_65.D ;
  assign g34002 = \DFF_1247.D ;
  assign g34003 = \DFF_457.D ;
  assign g34004 = \DFF_625.D ;
  assign g34005 = \DFF_469.D ;
  assign g34006 = \DFF_795.D ;
  assign g34007 = \DFF_4.D ;
  assign g34008 = \DFF_930.D ;
  assign g34009 = \DFF_887.D ;
  assign g3401 = \DFF_1298.Q ;
  assign g34010 = \DFF_1171.D ;
  assign g34011 = \DFF_1025.D ;
  assign g34012 = \DFF_959.D ;
  assign g34013 = \DFF_1115.D ;
  assign g34014 = \DFF_273.D ;
  assign g34015 = \DFF_61.D ;
  assign g34016 = \DFF_1097.D ;
  assign g34017 = \DFF_960.D ;
  assign g34018 = \DFF_890.D ;
  assign g34019 = \DFF_1380.D ;
  assign g34020 = \DFF_820.D ;
  assign g34021 = \DFF_727.D ;
  assign g34022 = \DFF_451.D ;
  assign g34023 = \DFF_228.D ;
  assign g34024 = \DFF_1265.D ;
  assign g34025 = \DFF_331.D ;
  assign g34026 = \DFF_107.D ;
  assign g34027 = \DFF_699.D ;
  assign g34028 = \DFF_635.D ;
  assign g34029 = \DFF_894.D ;
  assign g34030 = \DFF_412.D ;
  assign g34031 = \DFF_62.D ;
  assign g34032 = \DFF_849.D ;
  assign g34033 = \DFF_452.D ;
  assign g34034 = \DFF_130.D ;
  assign g34035 = \DFF_160.D ;
  assign g34036 = \DFF_99.D ;
  assign g34037 = \DFF_1199.D ;
  assign g34038 = \DFF_847.D ;
  assign g34039 = \DFF_914.D ;
  assign g34040 = \DFF_892.D ;
  assign g34041 = \DFF_218.D ;
  assign g34052 = \DFF_1111.D ;
  assign g34059 = \DFF_1220.D ;
  assign g3408 = \DFF_1239.Q ;
  assign g341 = \DFF_709.Q ;
  assign g34118 = \DFF_619.D ;
  assign g3412 = \DFF_513.Q ;
  assign g34121 = \DFF_1222.D ;
  assign g34122 = \DFF_761.D ;
  assign g34123 = \DFF_547.D ;
  assign g34126 = \DFF_355.D ;
  assign g34127 = g34425;
  assign g34130 = \DFF_1229.D ;
  assign g34131 = \DFF_790.D ;
  assign g34134 = \DFF_512.D ;
  assign g34142 = \DFF_1229.D ;
  assign g34144 = \DFF_790.D ;
  assign g34145 = \DFF_1222.D ;
  assign g34150 = \DFF_355.D ;
  assign g34151 = \DFF_547.D ;
  assign g34152 = \DFF_619.D ;
  assign g34153 = g34383;
  assign g34159 = \DFF_512.D ;
  assign g3416 = \DFF_1405.Q ;
  assign g34160 = \DFF_761.D ;
  assign g3419 = \DFF_578.Q ;
  assign g34195 = g31521;
  assign g34202 = g34201;
  assign g34208 = g34839;
  assign g34209 = g31656;
  assign g34210 = g31665;
  assign g34222 = g34221;
  assign g3423 = \DFF_801.Q ;
  assign g34232 = 1'b1;
  assign g34233 = 1'b1;
  assign g34234 = 1'b1;
  assign g34235 = 1'b1;
  assign g34236 = 1'b1;
  assign g34237 = 1'b1;
  assign g34238 = 1'b1;
  assign g34239 = 1'b1;
  assign g34240 = 1'b1;
  assign g34241 = \DFF_619.D ;
  assign g34242 = \DFF_1222.D ;
  assign g34243 = \DFF_761.D ;
  assign g34244 = \DFF_547.D ;
  assign g34245 = \DFF_355.D ;
  assign g34246 = \DFF_1229.D ;
  assign g34247 = \DFF_790.D ;
  assign g34248 = \DFF_512.D ;
  assign g34249 = \DFF_555.D ;
  assign g34250 = \DFF_359.D ;
  assign g34251 = \DFF_966.D ;
  assign g34252 = \DFF_50.D ;
  assign g34253 = \DFF_440.D ;
  assign g34254 = \DFF_965.D ;
  assign g34255 = \DFF_549.D ;
  assign g34256 = \DFF_1016.D ;
  assign g34257 = \DFF_1173.D ;
  assign g34258 = \DFF_1374.D ;
  assign g34259 = \DFF_186.D ;
  assign g34260 = \DFF_792.D ;
  assign g34261 = \DFF_1311.D ;
  assign g34262 = \DFF_609.D ;
  assign g34263 = \DFF_207.D ;
  assign g34264 = \DFF_1006.D ;
  assign g34265 = \DFF_935.D ;
  assign g34266 = \DFF_313.D ;
  assign g34267 = \DFF_78.D ;
  assign g34268 = \DFF_684.D ;
  assign g34269 = \DFF_922.D ;
  assign g34272 = g33935;
  assign g34273 = \DFF_673.Q ;
  assign g34274 = \DFF_767.Q ;
  assign g34275 = g33636;
  assign g34276 = g33659;
  assign g34277 = g31521;
  assign g34278 = \DFF_69.Q ;
  assign g34280 = \DFF_236.Q ;
  assign g34282 = \DFF_608.Q ;
  assign g34283 = \DFF_706.Q ;
  assign g34285 = \DFF_1111.D ;
  assign g34286 = \DFF_1357.Q ;
  assign g34288 = \DFF_994.Q ;
  assign g34289 = \DFF_881.Q ;
  assign g34290 = \DFF_1151.Q ;
  assign g34292 = \DFF_1301.Q ;
  assign g34293 = \DFF_1035.Q ;
  assign g34294 = \DFF_311.Q ;
  assign g34296 = \DFF_1220.D ;
  assign g34297 = \DFF_1403.Q ;
  assign g34300 = \DFF_15.Q ;
  assign g34302 = g31656;
  assign g34303 = \DFF_1336.Q ;
  assign g34304 = g31665;
  assign g34305 = \DFF_1289.Q ;
  assign g34306 = \DFF_1282.Q ;
  assign g3431 = \DFF_1168.Q ;
  assign g34314 = \DFF_196.Q ;
  assign g34318 = \DFF_657.Q ;
  assign g34321 = \DFF_144.Q ;
  assign g34331 = \DFF_489.Q ;
  assign g34347 = \DFF_190.Q ;
  assign g34349 = \DFF_80.Q ;
  assign g34350 = \DFF_75.Q ;
  assign g34352 = \DFF_64.Q ;
  assign g34353 = \DFF_498.Q ;
  assign g34358 = g34839;
  assign g3436 = \DFF_437.Q ;
  assign g34366 = \DFF_1340.Q ;
  assign g34368 = \DFF_507.Q ;
  assign g34369 = \DFF_974.Q ;
  assign g34372 = \DFF_941.Q ;
  assign g34373 = \DFF_1067.Q ;
  assign g34374 = \DFF_1041.Q ;
  assign g34376 = \DFF_445.Q ;
  assign g34377 = \DFF_1270.Q ;
  assign g34379 = \DFF_1319.Q ;
  assign g34384 = g34383;
  assign g34387 = g33874;
  assign g34391 = g33894;
  assign g34399 = \DFF_161.Q ;
  assign g344 = \DFF_686.Q ;
  assign g3440 = \DFF_180.Q ;
  assign g34402 = \DFF_177.Q ;
  assign g34403 = \DFF_766.Q ;
  assign g34404 = \DFF_1157.Q ;
  assign g34405 = \DFF_231.Q ;
  assign g34406 = \DFF_677.Q ;
  assign g34407 = \DFF_276.Q ;
  assign g34411 = \DFF_1193.Q ;
  assign g34412 = \DFF_721.Q ;
  assign g34416 = \DFF_855.Q ;
  assign g34417 = \DFF_1242.Q ;
  assign g34421 = \DFF_948.Q ;
  assign g34426 = g34425;
  assign g34427 = \DFF_619.D ;
  assign g34428 = \DFF_1222.D ;
  assign g34429 = \DFF_761.D ;
  assign g3443 = \DFF_830.Q ;
  assign g34430 = \DFF_547.D ;
  assign g34431 = \DFF_355.D ;
  assign g34432 = \DFF_1229.D ;
  assign g34433 = \DFF_790.D ;
  assign g34434 = \DFF_512.D ;
  assign g34435 = g31521;
  assign g34436 = g31656;
  assign g34437 = g31665;
  assign g34438 = \DFF_89.D ;
  assign g34439 = \DFF_789.D ;
  assign g34440 = \DFF_736.D ;
  assign g34441 = \DFF_1.D ;
  assign g34442 = \DFF_319.D ;
  assign g34443 = \DFF_1288.D ;
  assign g34444 = \DFF_931.D ;
  assign g34445 = \DFF_1112.D ;
  assign g34446 = \DFF_302.D ;
  assign g34447 = \DFF_284.D ;
  assign g34448 = \DFF_233.D ;
  assign g34449 = \DFF_1379.D ;
  assign g34450 = \DFF_1084.D ;
  assign g34451 = \DFF_358.D ;
  assign g34452 = \DFF_63.D ;
  assign g34453 = \DFF_718.D ;
  assign g34454 = \DFF_660.D ;
  assign g34455 = \DFF_115.D ;
  assign g34456 = \DFF_807.D ;
  assign g34457 = \DFF_1412.D ;
  assign g34458 = \DFF_674.D ;
  assign g34459 = \DFF_853.D ;
  assign g34460 = \DFF_43.D ;
  assign g34461 = \DFF_1373.D ;
  assign g34462 = \DFF_270.D ;
  assign g34463 = \DFF_461.D ;
  assign g34464 = \DFF_604.D ;
  assign g34465 = \DFF_1029.D ;
  assign g34466 = \DFF_1326.D ;
  assign g34467 = \DFF_985.D ;
  assign g34468 = \DFF_1107.D ;
  assign g3447 = \DFF_1414.Q ;
  assign g34471 = g34221;
  assign g34472 = \DFF_1111.D ;
  assign g34480 = \DFF_1220.D ;
  assign g34494 = \DFF_1125.Q ;
  assign g34501 = \DFF_1229.D ;
  assign g34504 = \DFF_790.D ;
  assign g34505 = \DFF_1222.D ;
  assign g3451 = \DFF_810.Q ;
  assign g34510 = \DFF_355.D ;
  assign g34511 = \DFF_547.D ;
  assign g34512 = \DFF_619.D ;
  assign g34521 = \DFF_512.D ;
  assign g34522 = \DFF_761.D ;
  assign g3454 = \DFF_492.Q ;
  assign g34540 = g34839;
  assign g3457 = \DFF_58.Q ;
  assign g34570 = g34201;
  assign g34579 = g33894;
  assign g34589 = \DFF_619.D ;
  assign g34590 = \DFF_1222.D ;
  assign g34591 = \DFF_761.D ;
  assign g34592 = \DFF_547.D ;
  assign g34593 = \DFF_355.D ;
  assign g34594 = \DFF_1229.D ;
  assign g34595 = \DFF_790.D ;
  assign g34596 = \DFF_512.D ;
  assign g34597 = 1'b0;
  assign g34598 = \DFF_489.D ;
  assign g34599 = \DFF_812.D ;
  assign g34600 = \DFF_896.D ;
  assign g34601 = \DFF_1242.D ;
  assign g34602 = \DFF_948.D ;
  assign g34603 = \DFF_507.D ;
  assign g34604 = \DFF_941.D ;
  assign g34605 = \DFF_445.D ;
  assign g34606 = \DFF_1067.D ;
  assign g34607 = \DFF_1270.D ;
  assign g34608 = \DFF_1319.D ;
  assign g34609 = \DFF_69.D ;
  assign g34610 = \DFF_236.D ;
  assign g34611 = \DFF_608.D ;
  assign g34612 = \DFF_1357.D ;
  assign g34613 = \DFF_994.D ;
  assign g34614 = \DFF_1301.D ;
  assign g34615 = \DFF_881.D ;
  assign g34616 = \DFF_1035.D ;
  assign g34617 = \DFF_15.D ;
  assign g34618 = \DFF_1336.D ;
  assign g34619 = \DFF_1289.D ;
  assign g3462 = \DFF_1134.Q ;
  assign g34620 = \DFF_1282.D ;
  assign g34621 = \DFF_1151.D ;
  assign g34622 = \DFF_311.D ;
  assign g34623 = \DFF_1403.D ;
  assign g34624 = \DFF_706.D ;
  assign g34625 = \DFF_196.D ;
  assign g34626 = \DFF_657.D ;
  assign g34627 = \DFF_144.D ;
  assign g34628 = \DFF_673.D ;
  assign g34629 = \DFF_767.D ;
  assign g34630 = \DFF_1340.D ;
  assign g34631 = \DFF_974.D ;
  assign g34632 = \DFF_1041.D ;
  assign g34633 = \DFF_1157.D ;
  assign g34634 = \DFF_677.D ;
  assign g34635 = \DFF_1193.D ;
  assign g34636 = \DFF_161.D ;
  assign g34637 = \DFF_177.D ;
  assign g34638 = \DFF_276.D ;
  assign g34639 = \DFF_721.D ;
  assign g34640 = \DFF_855.D ;
  assign g34641 = \DFF_766.D ;
  assign g34642 = \DFF_231.D ;
  assign g34643 = \DFF_190.D ;
  assign g34644 = \DFF_80.D ;
  assign g34645 = \DFF_75.D ;
  assign g34646 = \DFF_64.D ;
  assign g34647 = \DFF_498.D ;
  assign g34648 = \DFF_355.D ;
  assign g34649 = \DFF_1424.D ;
  assign g34650 = \DFF_1074.D ;
  assign g34653 = \DFF_547.D ;
  assign g34654 = \DFF_761.D ;
  assign g34656 = \DFF_1222.D ;
  assign g34657 = \DFF_417.D ;
  assign g34659 = \DFF_619.D ;
  assign g3466 = \DFF_688.Q ;
  assign g34660 = g34425;
  assign g34663 = \DFF_304.D ;
  assign g34688 = \DFF_1111.D ;
  assign g34690 = \DFF_1220.D ;
  assign g34699 = g34839;
  assign g347 = \DFF_1014.Q ;
  assign g3470 = \DFF_589.Q ;
  assign g34708 = \DFF_961.D ;
  assign g34711 = g34383;
  assign g34712 = g33894;
  assign g34713 = \DFF_512.D ;
  assign g34714 = \DFF_790.D ;
  assign g34716 = \DFF_1229.D ;
  assign g34717 = \DFF_1111.D ;
  assign g34718 = \DFF_1220.D ;
  assign g34719 = \DFF_593.D ;
  assign g34720 = \DFF_770.D ;
  assign g34721 = \DFF_715.D ;
  assign g34722 = \DFF_1253.D ;
  assign g34723 = \DFF_1391.D ;
  assign g34724 = \DFF_751.D ;
  assign g34725 = \DFF_953.D ;
  assign g34726 = \DFF_453.D ;
  assign g34727 = \DFF_127.D ;
  assign g34728 = \DFF_1314.D ;
  assign g34729 = \DFF_195.D ;
  assign g34730 = \DFF_323.D ;
  assign g34731 = \DFF_932.D ;
  assign g34732 = \DFF_1125.D ;
  assign g34733 = \DFF_25.D ;
  assign g34734 = \DFF_1000.D ;
  assign g34735 = \DFF_1417.D ;
  assign g34736 = \DFF_961.D ;
  assign g34739 = g33894;
  assign g34749 = \DFF_1074.D ;
  assign g34755 = \DFF_1424.D ;
  assign g34759 = \DFF_417.D ;
  assign g3476 = \DFF_341.Q ;
  assign g34760 = \DFF_304.D ;
  assign g34767 = \DFF_619.D ;
  assign g34768 = \DFF_512.D ;
  assign g34769 = \DFF_1222.D ;
  assign g34770 = \DFF_761.D ;
  assign g34772 = \DFF_547.D ;
  assign g34773 = \DFF_1074.D ;
  assign g34775 = \DFF_355.D ;
  assign g34776 = \DFF_1229.D ;
  assign g34777 = \DFF_790.D ;
  assign g34778 = g34839;
  assign g34781 = \DFF_379.D ;
  assign g34783 = \DFF_796.D ;
  assign g34784 = \DFF_1074.D ;
  assign g34785 = \DFF_961.D ;
  assign g34786 = \DFF_1424.D ;
  assign g34787 = \DFF_417.D ;
  assign g34788 = g33894;
  assign g34789 = \DFF_304.D ;
  assign g34790 = \DFF_119.D ;
  assign g34791 = \DFF_1200.D ;
  assign g34792 = \DFF_364.D ;
  assign g34793 = \DFF_1182.D ;
  assign g34794 = \DFF_781.D ;
  assign g34795 = \DFF_223.D ;
  assign g34796 = \DFF_757.D ;
  assign g34797 = \DFF_749.D ;
  assign g34798 = \DFF_242.D ;
  assign g34799 = \DFF_1178.D ;
  assign g3480 = \DFF_778.Q ;
  assign g34800 = \DFF_197.D ;
  assign g34801 = \DFF_531.D ;
  assign g34802 = \DFF_899.D ;
  assign g34803 = \DFF_852.D ;
  assign g34804 = \DFF_399.D ;
  assign g34805 = \DFF_1245.D ;
  assign g34806 = \DFF_155.D ;
  assign g34807 = \DFF_95.D ;
  assign g34808 = \DFF_733.D ;
  assign g34809 = \DFF_743.D ;
  assign g34810 = \DFF_379.D ;
  assign g34812 = \DFF_796.D ;
  assign g34813 = \DFF_619.D ;
  assign g34816 = \DFF_512.D ;
  assign g34820 = \DFF_1222.D ;
  assign g34823 = \DFF_761.D ;
  assign g34827 = \DFF_547.D ;
  assign g34830 = \DFF_355.D ;
  assign g34833 = \DFF_1229.D ;
  assign g34836 = \DFF_790.D ;
  assign g3484 = \DFF_955.Q ;
  assign g34840 = g34839;
  assign g34843 = \DFF_1181.D ;
  assign g34846 = \DFF_1074.D ;
  assign g34847 = \DFF_796.D ;
  assign g34848 = \DFF_379.D ;
  assign g34849 = \DFF_844.D ;
  assign g34850 = \DFF_661.D ;
  assign g34851 = \DFF_1181.D ;
  assign g34852 = \DFF_1074.D ;
  assign g34855 = \DFF_743.D ;
  assign g34877 = \DFF_1074.D ;
  assign g34878 = \DFF_743.D ;
  assign g34879 = \DFF_1181.D ;
  assign g34880 = \DFF_338.D ;
  assign g34881 = \DFF_21.D ;
  assign g34882 = \DFF_26.D ;
  assign g34884 = g34915;
  assign g34887 = g34927;
  assign g34890 = g34925;
  assign g34893 = \DFF_1074.D ;
  assign g34894 = g34923;
  assign g34897 = g34921;
  assign g3490 = \DFF_29.Q ;
  assign g34900 = g34919;
  assign g34903 = g34917;
  assign g34906 = g34913;
  assign g34910 = g34839;
  assign g34911 = \DFF_142.D ;
  assign g34914 = g34913;
  assign g34916 = g34915;
  assign g34918 = g34917;
  assign g34920 = g34919;
  assign g34922 = g34921;
  assign g34924 = g34923;
  assign g34926 = g34925;
  assign g34928 = g34927;
  assign g34929 = \DFF_1074.D ;
  assign g34930 = g34839;
  assign g34935 = \DFF_1074.D ;
  assign g3494 = \DFF_243.Q ;
  assign g34943 = g34839;
  assign g34944 = g34913;
  assign g34945 = g34915;
  assign g34946 = g34917;
  assign g34947 = g34919;
  assign g34949 = g34921;
  assign g34950 = g34923;
  assign g34951 = g34925;
  assign g34952 = g34927;
  assign g34954 = g34839;
  assign g34956 = g34839;
  assign g34957 = g34972;
  assign g34970 = \DFF_514.D ;
  assign g34971 = \DFF_206.D ;
  assign g34973 = g34972;
  assign g34974 = \DFF_477.D ;
  assign g34975 = \DFF_829.D ;
  assign g34976 = \DFF_150.D ;
  assign g34977 = \DFF_1322.D ;
  assign g34978 = \DFF_1012.D ;
  assign g34979 = \DFF_420.D ;
  assign g3498 = \DFF_559.Q ;
  assign g34980 = \DFF_413.D ;
  assign g34982 = \DFF_514.D ;
  assign g34983 = \DFF_206.D ;
  assign g34984 = \DFF_477.D ;
  assign g34985 = \DFF_829.D ;
  assign g34986 = \DFF_150.D ;
  assign g34987 = \DFF_1322.D ;
  assign g34988 = \DFF_1012.D ;
  assign g34989 = \DFF_420.D ;
  assign g34990 = \DFF_514.D ;
  assign g34991 = \DFF_477.D ;
  assign g34992 = \DFF_829.D ;
  assign g34993 = \DFF_150.D ;
  assign g34994 = \DFF_1322.D ;
  assign g34995 = \DFF_1012.D ;
  assign g34996 = \DFF_420.D ;
  assign g34997 = \DFF_206.D ;
  assign g34998 = g34972;
  assign g35000 = \DFF_621.D ;
  assign g35001 = \DFF_621.D ;
  assign g35002 = \DFF_621.D ;
  assign g3502 = \DFF_657.Q ;
  assign g3506 = \DFF_120.Q ;
  assign g351 = \DFF_240.Q ;
  assign g3512 = \DFF_27.Q ;
  assign g3518 = \DFF_245.Q ;
  assign g3522 = \DFF_1408.Q ;
  assign g3530 = \DFF_199.Q ;
  assign g3538 = \DFF_707.Q ;
  assign g3542 = \DFF_12.Q ;
  assign g3546 = \DFF_982.Q ;
  assign g355 = \DFF_294.Q ;
  assign g3550 = \DFF_1259.Q ;
  assign g3554 = \DFF_19.Q ;
  assign g3558 = \DFF_309.Q ;
  assign g3562 = \DFF_738.Q ;
  assign g3566 = \DFF_227.Q ;
  assign g3570 = \DFF_108.Q ;
  assign g3574 = \DFF_321.Q ;
  assign g3578 = \DFF_628.Q ;
  assign g358 = \DFF_798.Q ;
  assign g3582 = \DFF_633.Q ;
  assign g3586 = \DFF_105.Q ;
  assign g3590 = \DFF_1052.Q ;
  assign g3594 = \DFF_1244.Q ;
  assign g3598 = \DFF_72.Q ;
  assign g3602 = \DFF_626.Q ;
  assign g3606 = \DFF_102.Q ;
  assign g3610 = \DFF_1177.Q ;
  assign g3614 = \DFF_1356.Q ;
  assign g3618 = \DFF_220.Q ;
  assign g3625 = \DFF_81.Q ;
  assign g3632 = \DFF_468.Q ;
  assign g3639 = \DFF_536.Q ;
  assign g3649 = \DFF_34.Q ;
  assign g365 = \DFF_269.Q ;
  assign g3654 = \DFF_1420.Q ;
  assign g3661 = \DFF_942.Q ;
  assign g3668 = \DFF_873.Q ;
  assign g3672 = \DFF_369.Q ;
  assign g3676 = \DFF_1300.Q ;
  assign g3680 = \DFF_290.Q ;
  assign g3684 = \DFF_535.Q ;
  assign g3689 = \DFF_664.Q ;
  assign g3694 = \DFF_1214.Q ;
  assign g3698 = \DFF_39.Q ;
  assign g37 = \DFF_994.Q ;
  assign g370 = \DFF_1161.Q ;
  assign g3703 = \DFF_1312.Q ;
  assign g3706 = \DFF_516.Q ;
  assign g3712 = \DFF_405.Q ;
  assign g3719 = \DFF_475.Q ;
  assign g3723 = \DFF_741.Q ;
  assign g3727 = \DFF_1309.Q ;
  assign g3731 = \DFF_1077.Q ;
  assign g3736 = \DFF_335.Q ;
  assign g3742 = \DFF_381.Q ;
  assign g3747 = \DFF_1334.Q ;
  assign g3752 = \DFF_478.Q ;
  assign g3759 = \DFF_548.Q ;
  assign g376 = \DFF_1232.Q ;
  assign g3763 = \DFF_1385.Q ;
  assign g3767 = \DFF_631.Q ;
  assign g3770 = \DFF_495.Q ;
  assign g3774 = \DFF_701.Q ;
  assign g3782 = \DFF_939.Q ;
  assign g3787 = \DFF_523.Q ;
  assign g3791 = \DFF_540.Q ;
  assign g3794 = \DFF_147.Q ;
  assign g3798 = \DFF_460.Q ;
  assign g3802 = \DFF_299.Q ;
  assign g3805 = \DFF_450.Q ;
  assign g3808 = \DFF_546.Q ;
  assign g3813 = \DFF_87.Q ;
  assign g3817 = \DFF_742.Q ;
  assign g3821 = \DFF_1360.Q ;
  assign g3827 = \DFF_693.Q ;
  assign g3831 = \DFF_441.Q ;
  assign g3835 = \DFF_274.Q ;
  assign g3841 = \DFF_1383.Q ;
  assign g3845 = \DFF_1260.Q ;
  assign g3849 = \DFF_1195.Q ;
  assign g385 = \DFF_1393.Q ;
  assign g3853 = \DFF_144.Q ;
  assign g3857 = \DFF_784.Q ;
  assign g3863 = \DFF_776.Q ;
  assign g3869 = \DFF_473.Q ;
  assign g3873 = \DFF_467.Q ;
  assign g3881 = \DFF_587.Q ;
  assign g3889 = \DFF_340.Q ;
  assign g3893 = \DFF_1350.Q ;
  assign g3897 = \DFF_590.Q ;
  assign g3901 = \DFF_312.Q ;
  assign g3905 = \DFF_156.Q ;
  assign g3909 = \DFF_91.Q ;
  assign g391 = \DFF_1099.Q ;
  assign g3913 = \DFF_1264.Q ;
  assign g3917 = \DFF_479.Q ;
  assign g392 = \DFF_1053.Q ;
  assign g3921 = \DFF_1128.Q ;
  assign g3925 = \DFF_986.Q ;
  assign g3929 = \DFF_917.Q ;
  assign g3933 = \DFF_257.Q ;
  assign g3937 = \DFF_868.Q ;
  assign g3941 = \DFF_1160.Q ;
  assign g3945 = \DFF_1013.Q ;
  assign g3949 = \DFF_947.Q ;
  assign g3953 = \DFF_1317.Q ;
  assign g3957 = \DFF_550.Q ;
  assign g3961 = \DFF_414.Q ;
  assign g3965 = \DFF_253.Q ;
  assign g3969 = \DFF_181.Q ;
  assign g3976 = \DFF_785.Q ;
  assign g3983 = \DFF_401.Q ;
  assign g3990 = \DFF_517.Q ;
  assign g4000 = \DFF_642.Q ;
  assign g4005 = \DFF_1001.Q ;
  assign g401 = \DFF_542.Q ;
  assign g4012 = \DFF_305.Q ;
  assign g4019 = \DFF_367.Q ;
  assign g4023 = \DFF_662.Q ;
  assign g4027 = \DFF_1219.Q ;
  assign g4031 = \DFF_995.Q ;
  assign g4035 = \DFF_857.Q ;
  assign g4040 = \DFF_5.Q ;
  assign g4045 = \DFF_423.Q ;
  assign g4049 = \DFF_347.Q ;
  assign g405 = \DFF_601.Q ;
  assign g4054 = \DFF_286.Q ;
  assign g4057 = \DFF_1324.Q ;
  assign g4064 = \DFF_891.Q ;
  assign g4072 = \DFF_685.Q ;
  assign g4076 = \DFF_154.Q ;
  assign g4082 = \DFF_860.Q ;
  assign g4087 = \DFF_411.Q ;
  assign g4093 = \DFF_551.Q ;
  assign g4098 = \DFF_351.Q ;
  assign g4104 = \DFF_201.Q ;
  assign g4108 = \DFF_508.Q ;
  assign g411 = \DFF_1315.Q ;
  assign g4112 = \DFF_1139.Q ;
  assign g4116 = \DFF_689.Q ;
  assign g4119 = \DFF_1187.Q ;
  assign g4122 = \DFF_1083.Q ;
  assign g4125 = \DFF_1204.Q ;
  assign g4129 = \DFF_1152.Q ;
  assign g4132 = \DFF_114.Q ;
  assign g4135 = \DFF_247.Q ;
  assign g4138 = \DFF_330.Q ;
  assign g4141 = \DFF_1361.Q ;
  assign g4145 = \DFF_1230.Q ;
  assign g4146 = \DFF_673.Q ;
  assign g4153 = \DFF_116.Q ;
  assign g4157 = \DFF_767.Q ;
  assign g4164 = \DFF_282.Q ;
  assign g4165 = \DFF_527.Q ;
  assign g4169 = \DFF_434.Q ;
  assign g417 = \DFF_237.Q ;
  assign g4172 = \DFF_25.Q ;
  assign g4176 = \DFF_1000.Q ;
  assign g4180 = \DFF_1389.Q ;
  assign g4185 = \DFF_389.Q ;
  assign g4188 = \DFF_480.Q ;
  assign g4191 = \DFF_1234.Q ;
  assign g4194 = \DFF_909.Q ;
  assign g4197 = \DFF_565.Q ;
  assign g4200 = \DFF_1224.Q ;
  assign g4204 = \DFF_1416.Q ;
  assign g4207 = \DFF_1049.Q ;
  assign g4210 = \DFF_704.Q ;
  assign g4213 = \DFF_1286.Q ;
  assign g4216 = \DFF_485.Q ;
  assign g4219 = \DFF_992.Q ;
  assign g4222 = \DFF_885.Q ;
  assign g4226 = \DFF_418.Q ;
  assign g4229 = \DFF_944.Q ;
  assign g4232 = \DFF_1338.Q ;
  assign g4235 = \DFF_31.Q ;
  assign g4239 = \DFF_1387.Q ;
  assign g424 = \DFF_1108.Q ;
  assign g4242 = \DFF_919.Q ;
  assign g4245 = \DFF_1041.Q ;
  assign g4249 = \DFF_974.Q ;
  assign g4253 = \DFF_1340.Q ;
  assign g4258 = \DFF_1190.Q ;
  assign g4264 = \DFF_73.Q ;
  assign g4269 = \DFF_215.Q ;
  assign g4273 = \DFF_210.Q ;
  assign g4277 = \DFF_831.Q ;
  assign g4281 = \DFF_320.Q ;
  assign g4284 = \DFF_1384.Q ;
  assign g4287 = \DFF_1027.Q ;
  assign g429 = \DFF_972.Q ;
  assign g4291 = \DFF_1043.Q ;
  assign g4294 = \DFF_739.Q ;
  assign g4297 = \DFF_325.Q ;
  assign g43 = \DFF_304.Q ;
  assign g4300 = \DFF_1417.Q ;
  assign g4304 = \DFF_203.Q ;
  assign g4308 = \DFF_509.Q ;
  assign g4311 = \DFF_1379.Q ;
  assign g4322 = \DFF_1084.Q ;
  assign g433 = \DFF_324.Q ;
  assign g4332 = \DFF_115.Q ;
  assign g4340 = \DFF_853.Q ;
  assign g4349 = \DFF_1173.Q ;
  assign g4358 = \DFF_1374.Q ;
  assign g4366 = \DFF_1299.Q ;
  assign g4369 = \DFF_436.Q ;
  assign g437 = \DFF_239.Q ;
  assign g4372 = \DFF_26.Q ;
  assign g4375 = \DFF_159.Q ;
  assign g4382 = \DFF_250.Q ;
  assign g4388 = \DFF_482.Q ;
  assign g4392 = \DFF_980.Q ;
  assign g4401 = \DFF_1146.Q ;
  assign g4405 = \DFF_1002.Q ;
  assign g4408 = \DFF_1073.Q ;
  assign g441 = \DFF_544.Q ;
  assign g4411 = \DFF_613.Q ;
  assign g4414 = \DFF_234.Q ;
  assign g4417 = \DFF_1272.Q ;
  assign g4420 = \DFF_1397.Q ;
  assign g4423 = \DFF_663.Q ;
  assign g4427 = \DFF_1221.Q ;
  assign g4430 = \DFF_490.Q ;
  assign g4434 = \DFF_692.Q ;
  assign g4438 = \DFF_929.Q ;
  assign g4443 = \DFF_687.Q ;
  assign g4446 = \DFF_1225.Q ;
  assign g4449 = \DFF_348.Q ;
  assign g4452 = \DFF_373.Q ;
  assign g4455 = \DFF_530.Q ;
  assign g4456 = \DFF_1305.Q ;
  assign g4459 = \DFF_440.Q ;
  assign g446 = \DFF_1164.Q ;
  assign g4462 = \DFF_965.Q ;
  assign g4467 = \DFF_549.Q ;
  assign g4473 = \DFF_1016.Q ;
  assign g4474 = \DFF_615.Q ;
  assign g4477 = \DFF_184.Q ;
  assign g4480 = \DFF_624.Q ;
  assign g4483 = \DFF_1209.Q ;
  assign g4486 = \DFF_383.Q ;
  assign g4489 = \DFF_911.Q ;
  assign g4492 = \DFF_129.Q ;
  assign g4495 = \DFF_268.Q ;
  assign g4498 = \DFF_352.Q ;
  assign g45 = \DFF_514.Q ;
  assign g4501 = \DFF_744.Q ;
  assign g4504 = \DFF_384.Q ;
  assign g4507 = \DFF_1399.Q ;
  assign g4512 = \DFF_1296.Q ;
  assign g4515 = \DFF_1415.Q ;
  assign g4519 = \DFF_1345.Q ;
  assign g452 = \DFF_10.Q ;
  assign g4520 = \DFF_991.Q ;
  assign g4521 = \DFF_79.Q ;
  assign g4527 = \DFF_813.Q ;
  assign g4531 = \DFF_607.Q ;
  assign g4534 = \DFF_228.Q ;
  assign g4537 = \DFF_1265.Q ;
  assign g4540 = \DFF_1022.Q ;
  assign g4543 = \DFF_226.Q ;
  assign g4546 = \DFF_816.Q ;
  assign g4549 = \DFF_1330.Q ;
  assign g4552 = \DFF_1349.Q ;
  assign g4555 = \DFF_38.Q ;
  assign g4558 = \DFF_121.Q ;
  assign g4561 = \DFF_808.Q ;
  assign g4564 = \DFF_491.Q ;
  assign g4567 = \DFF_56.Q ;
  assign g457 = \DFF_427.Q ;
  assign g4570 = \DFF_1362.Q ;
  assign g4571 = \DFF_528.Q ;
  assign g4572 = \DFF_221.Q ;
  assign g4575 = \DFF_350.Q ;
  assign g4578 = \DFF_439.Q ;
  assign g4581 = \DFF_724.Q ;
  assign g4584 = \DFF_358.Q ;
  assign g4593 = \DFF_63.Q ;
  assign g46 = \DFF_477.Q ;
  assign g460 = \DFF_652.Q ;
  assign g4601 = \DFF_718.Q ;
  assign g4608 = \DFF_660.Q ;
  assign g4616 = \DFF_807.Q ;
  assign g4621 = \DFF_43.Q ;
  assign g4628 = \DFF_1412.Q ;
  assign g4633 = \DFF_674.Q ;
  assign g4639 = \DFF_331.Q ;
  assign g464 = \DFF_11.Q ;
  assign g4643 = \DFF_186.Q ;
  assign g4646 = \DFF_792.Q ;
  assign g4653 = \DFF_270.Q ;
  assign g4659 = \DFF_1373.Q ;
  assign g4664 = \DFF_461.Q ;
  assign g4669 = \DFF_604.Q ;
  assign g4674 = \DFF_107.Q ;
  assign g468 = \DFF_629.Q ;
  assign g4681 = \DFF_699.Q ;
  assign g4688 = \DFF_635.Q ;
  assign g4698 = \DFF_1311.Q ;
  assign g47 = \DFF_829.Q ;
  assign g4704 = \DFF_747.Q ;
  assign g4709 = \DFF_849.Q ;
  assign g471 = \DFF_430.Q ;
  assign g4717 = \DFF_1193.Q ;
  assign g4722 = \DFF_161.Q ;
  assign g4727 = \DFF_1157.Q ;
  assign g4732 = \DFF_677.Q ;
  assign g4737 = \DFF_177.Q ;
  assign g4741 = \DFF_501.Q ;
  assign g4742 = \DFF_200.Q ;
  assign g4743 = \DFF_609.Q ;
  assign g4749 = \DFF_254.Q ;
  assign g475 = \DFF_510.Q ;
  assign g4754 = \DFF_207.Q ;
  assign g4760 = \DFF_647.Q ;
  assign g4765 = \DFF_1006.Q ;
  assign g4771 = \DFF_837.Q ;
  assign g4776 = \DFF_62.Q ;
  assign g4785 = \DFF_894.Q ;
  assign g479 = \DFF_252.Q ;
  assign g4793 = \DFF_452.Q ;
  assign g48 = \DFF_150.Q ;
  assign g4801 = \DFF_412.Q ;
  assign g4809 = \DFF_178.Q ;
  assign g4812 = \DFF_997.Q ;
  assign g4815 = \DFF_1118.Q ;
  assign g4818 = \DFF_1191.Q ;
  assign g482 = \DFF_1145.Q ;
  assign g4821 = \DFF_1205.Q ;
  assign g4826 = \DFF_493.Q ;
  assign g4831 = \DFF_249.Q ;
  assign g4836 = \DFF_935.Q ;
  assign g4843 = \DFF_1326.Q ;
  assign g4849 = \DFF_1029.Q ;
  assign g4854 = \DFF_985.Q ;
  assign g4859 = \DFF_1107.Q ;
  assign g4864 = \DFF_130.Q ;
  assign g4871 = \DFF_160.Q ;
  assign g4878 = \DFF_99.Q ;
  assign g4888 = \DFF_313.Q ;
  assign g4894 = \DFF_782.Q ;
  assign g4899 = \DFF_892.Q ;
  assign g49 = \DFF_1322.Q ;
  assign g490 = \DFF_47.Q ;
  assign g4907 = \DFF_855.Q ;
  assign g4912 = \DFF_766.Q ;
  assign g4917 = \DFF_276.Q ;
  assign g4922 = \DFF_721.Q ;
  assign g4927 = \DFF_231.Q ;
  assign g4931 = \DFF_1402.Q ;
  assign g4932 = \DFF_1165.Q ;
  assign g4933 = \DFF_78.Q ;
  assign g4939 = \DFF_1206.Q ;
  assign g4944 = \DFF_684.Q ;
  assign g4950 = \DFF_574.Q ;
  assign g4955 = \DFF_922.Q ;
  assign g496 = \DFF_143.Q ;
  assign g4961 = \DFF_229.Q ;
  assign g4966 = \DFF_914.Q ;
  assign g4975 = \DFF_1199.Q ;
  assign g4983 = \DFF_218.Q ;
  assign g499 = \DFF_786.Q ;
  assign g4991 = \DFF_847.Q ;
  assign g4999 = \DFF_672.Q ;
  assign g50 = \DFF_1012.Q ;
  assign g5002 = \DFF_981.Q ;
  assign g5005 = \DFF_1100.Q ;
  assign g5008 = \DFF_1176.Q ;
  assign g5011 = \DFF_714.Q ;
  assign g5016 = \DFF_1341.Q ;
  assign g5022 = \DFF_366.Q ;
  assign g5029 = \DFF_432.Q ;
  assign g5033 = \DFF_1192.Q ;
  assign g5037 = \DFF_386.Q ;
  assign g504 = \DFF_622.Q ;
  assign g5041 = \DFF_690.Q ;
  assign g5046 = \DFF_1327.Q ;
  assign g5052 = \DFF_502.Q ;
  assign g5057 = \DFF_0.Q ;
  assign g5062 = \DFF_1065.Q ;
  assign g5069 = \DFF_1124.Q ;
  assign g5073 = \DFF_1116.Q ;
  assign g5077 = \DFF_288.Q ;
  assign g5080 = \DFF_722.Q ;
  assign g5084 = \DFF_883.Q ;
  assign g5092 = \DFF_248.Q ;
  assign g5097 = \DFF_1217.Q ;
  assign g51 = \DFF_420.Q ;
  assign g5101 = \DFF_678.Q ;
  assign g5105 = \DFF_545.Q ;
  assign g5109 = \DFF_458.Q ;
  assign g5112 = \DFF_1228.Q ;
  assign g5115 = \DFF_1346.Q ;
  assign g5120 = \DFF_926.Q ;
  assign g5124 = \DFF_1121.Q ;
  assign g5128 = \DFF_1370.Q ;
  assign g513 = \DFF_447.Q ;
  assign g5134 = \DFF_145.Q ;
  assign g5138 = \DFF_456.Q ;
  assign g5142 = \DFF_1211.Q ;
  assign g5148 = \DFF_1398.Q ;
  assign g5152 = \DFF_1284.Q ;
  assign g5156 = \DFF_826.Q ;
  assign g5160 = \DFF_190.Q ;
  assign g5164 = \DFF_407.Q ;
  assign g5170 = \DFF_1304.Q ;
  assign g5176 = \DFF_1098.Q ;
  assign g518 = \DFF_591.Q ;
  assign g5180 = \DFF_68.Q ;
  assign g5188 = \DFF_598.Q ;
  assign g5196 = \DFF_638.Q ;
  assign g52 = \DFF_206.Q ;
  assign g5200 = \DFF_1325.Q ;
  assign g5204 = \DFF_100.Q ;
  assign g5208 = \DFF_390.Q ;
  assign g5212 = \DFF_1040.Q ;
  assign g5216 = \DFF_602.Q ;
  assign g5220 = \DFF_750.Q ;
  assign g5224 = \DFF_923.Q ;
  assign g5228 = \DFF_1186.Q ;
  assign g5232 = \DFF_13.Q ;
  assign g5236 = \DFF_983.Q ;
  assign g5240 = \DFF_773.Q ;
  assign g5244 = \DFF_950.Q ;
  assign g5248 = \DFF_1212.Q ;
  assign g5252 = \DFF_1095.Q ;
  assign g5256 = \DFF_659.Q ;
  assign g5260 = \DFF_1406.Q ;
  assign g5264 = \DFF_187.Q ;
  assign g5268 = \DFF_497.Q ;
  assign g5272 = \DFF_1363.Q ;
  assign g5276 = \DFF_906.Q ;
  assign g528 = \DFF_353.Q ;
  assign g5283 = \DFF_566.Q ;
  assign g5290 = \DFF_655.Q ;
  assign g5297 = \DFF_449.Q ;
  assign g5308 = \DFF_616.Q ;
  assign g5313 = \DFF_165.Q ;
  assign g5320 = \DFF_927.Q ;
  assign g5327 = \DFF_765.Q ;
  assign g5331 = \DFF_537.Q ;
  assign g5335 = \DFF_360.Q ;
  assign g5339 = \DFF_281.Q ;
  assign g534 = \DFF_1391.Q ;
  assign g5343 = \DFF_141.Q ;
  assign g5348 = \DFF_1400.Q ;
  assign g5352 = \DFF_1285.Q ;
  assign g5357 = \DFF_846.Q ;
  assign g5360 = \DFF_191.Q ;
  assign g5366 = \DFF_1392.Q ;
  assign g5373 = \DFF_557.Q ;
  assign g5377 = \DFF_1132.Q ;
  assign g538 = \DFF_593.Q ;
  assign g5381 = \DFF_665.Q ;
  assign g5385 = \DFF_518.Q ;
  assign g5390 = \DFF_823.Q ;
  assign g5396 = \DFF_639.Q ;
  assign g5401 = \DFF_1238.Q ;
  assign g5406 = \DFF_539.Q ;
  assign g5413 = \DFF_787.Q ;
  assign g5417 = \DFF_1367.Q ;
  assign g542 = \DFF_597.Q ;
  assign g5421 = \DFF_668.Q ;
  assign g5424 = \DFF_285.Q ;
  assign g5428 = \DFF_605.Q ;
  assign g5436 = \DFF_354.Q ;
  assign g5441 = \DFF_691.Q ;
  assign g5445 = \DFF_556.Q ;
  assign g5448 = \DFF_630.Q ;
  assign g5452 = \DFF_503.Q ;
  assign g5456 = \DFF_1396.Q ;
  assign g5459 = \DFF_569.Q ;
  assign g546 = \DFF_1253.Q ;
  assign g5462 = \DFF_1066.Q ;
  assign g5467 = \DFF_651.Q ;
  assign g5471 = \DFF_1021.Q ;
  assign g5475 = \DFF_875.Q ;
  assign g5481 = \DFF_1215.Q ;
  assign g5485 = \DFF_1079.Q ;
  assign g5489 = \DFF_1018.Q ;
  assign g5495 = \DFF_388.Q ;
  assign g5499 = \DFF_310.Q ;
  assign g55 = \DFF_621.Q ;
  assign g550 = \DFF_770.Q ;
  assign g5503 = \DFF_918.Q ;
  assign g5507 = \DFF_80.Q ;
  assign g5511 = \DFF_244.Q ;
  assign g5517 = \DFF_958.Q ;
  assign g5523 = \DFF_289.Q ;
  assign g5527 = \DFF_910.Q ;
  assign g5535 = \DFF_575.Q ;
  assign g554 = \DFF_142.Q ;
  assign g5543 = \DFF_333.Q ;
  assign g5547 = \DFF_938.Q ;
  assign g5551 = \DFF_307.Q ;
  assign g5555 = \DFF_151.Q ;
  assign g5559 = \DFF_84.Q ;
  assign g5563 = \DFF_1007.Q ;
  assign g5567 = \DFF_172.Q ;
  assign g5571 = \DFF_627.Q ;
  assign g5575 = \DFF_476.Q ;
  assign g5579 = \DFF_392.Q ;
  assign g5583 = \DFF_895.Q ;
  assign g5587 = \DFF_51.Q ;
  assign g559 = \DFF_7.Q ;
  assign g5591 = \DFF_71.Q ;
  assign g5595 = \DFF_1355.Q ;
  assign g5599 = \DFF_1297.Q ;
  assign g5603 = \DFF_884.Q ;
  assign g5607 = \DFF_44.Q ;
  assign g5611 = \DFF_219.Q ;
  assign g5615 = \DFF_55.Q ;
  assign g5619 = \DFF_1423.Q ;
  assign g562 = \DFF_88.Q ;
  assign g5623 = \DFF_263.Q ;
  assign g5630 = \DFF_101.Q ;
  assign g5637 = \DFF_1335.Q ;
  assign g5644 = \DFF_1283.Q ;
  assign g5654 = \DFF_1352.Q ;
  assign g5659 = \DFF_46.Q ;
  assign g5666 = \DFF_117.Q ;
  assign g5673 = \DFF_695.Q ;
  assign g5677 = \DFF_1262.Q ;
  assign g568 = \DFF_728.Q ;
  assign g5681 = \DFF_783.Q ;
  assign g5685 = \DFF_666.Q ;
  assign g5689 = \DFF_599.Q ;
  assign g5694 = \DFF_1162.Q ;
  assign g5698 = \DFF_1404.Q ;
  assign g5703 = \DFF_1252.Q ;
  assign g5706 = \DFF_426.Q ;
  assign g5712 = \DFF_329.Q ;
  assign g5719 = \DFF_394.Q ;
  assign g572 = \DFF_506.Q ;
  assign g5723 = \DFF_676.Q ;
  assign g5727 = \DFF_1246.Q ;
  assign g5731 = \DFF_1015.Q ;
  assign g5736 = \DFF_260.Q ;
  assign g5742 = \DFF_308.Q ;
  assign g5747 = \DFF_1271.Q ;
  assign g5752 = \DFF_396.Q ;
  assign g5759 = \DFF_466.Q ;
  assign g5763 = \DFF_1333.Q ;
  assign g5767 = \DFF_572.Q ;
  assign g577 = \DFF_863.Q ;
  assign g5770 = \DFF_415.Q ;
  assign g5774 = \DFF_636.Q ;
  assign g5782 = \DFF_869.Q ;
  assign g5787 = \DFF_438.Q ;
  assign g5791 = \DFF_459.Q ;
  assign g5794 = \DFF_85.Q ;
  assign g5798 = \DFF_376.Q ;
  assign g5802 = \DFF_235.Q ;
  assign g5805 = \DFF_365.Q ;
  assign g5808 = \DFF_463.Q ;
  assign g5813 = \DFF_14.Q ;
  assign g5817 = \DFF_679.Q ;
  assign g582 = \DFF_1235.Q ;
  assign g5821 = \DFF_1306.Q ;
  assign g5827 = \DFF_632.Q ;
  assign g5831 = \DFF_361.Q ;
  assign g5835 = \DFF_213.Q ;
  assign g5841 = \DFF_1332.Q ;
  assign g5845 = \DFF_1198.Q ;
  assign g5849 = \DFF_1138.Q ;
  assign g5853 = \DFF_75.Q ;
  assign g5857 = \DFF_734.Q ;
  assign g586 = \DFF_560.Q ;
  assign g5863 = \DFF_723.Q ;
  assign g5869 = \DFF_393.Q ;
  assign g5873 = \DFF_385.Q ;
  assign g5881 = \DFF_519.Q ;
  assign g5889 = \DFF_267.Q ;
  assign g5893 = \DFF_1291.Q ;
  assign g5897 = \DFF_526.Q ;
  assign g59 = \DFF_1425.Q ;
  assign g590 = \DFF_162.Q ;
  assign g5901 = \DFF_241.Q ;
  assign g5905 = \DFF_93.Q ;
  assign g5909 = \DFF_17.Q ;
  assign g5913 = \DFF_1201.Q ;
  assign g5917 = \DFF_398.Q ;
  assign g5921 = \DFF_1058.Q ;
  assign g5925 = \DFF_920.Q ;
  assign g5929 = \DFF_854.Q ;
  assign g5933 = \DFF_192.Q ;
  assign g5937 = \DFF_815.Q ;
  assign g5941 = \DFF_1085.Q ;
  assign g5945 = \DFF_949.Q ;
  assign g5949 = \DFF_877.Q ;
  assign g595 = \DFF_1090.Q ;
  assign g5953 = \DFF_1255.Q ;
  assign g5957 = \DFF_471.Q ;
  assign g5961 = \DFF_336.Q ;
  assign g5965 = \DFF_183.Q ;
  assign g5969 = \DFF_110.Q ;
  assign g5976 = \DFF_737.Q ;
  assign g5983 = \DFF_326.Q ;
  assign g599 = \DFF_874.Q ;
  assign g5990 = \DFF_429.Q ;
  assign g6 = \DFF_619.Q ;
  assign g6000 = \DFF_1087.Q ;
  assign g6005 = \DFF_30.Q ;
  assign g6012 = \DFF_797.Q ;
  assign g6019 = \DFF_848.Q ;
  assign g6023 = \DFF_1102.Q ;
  assign g6027 = \DFF_279.Q ;
  assign g6031 = \DFF_22.Q ;
  assign g6035 = \DFF_1320.Q ;
  assign g604 = \DFF_966.Q ;
  assign g6040 = \DFF_543.Q ;
  assign g6044 = \DFF_731.Q ;
  assign g6049 = \DFF_833.Q ;
  assign g6052 = \DFF_851.Q ;
  assign g6058 = \DFF_1048.Q ;
  assign g6065 = \DFF_122.Q ;
  assign g6069 = \DFF_49.Q ;
  assign g6073 = \DFF_40.Q ;
  assign g6077 = \DFF_712.Q ;
  assign g608 = \DFF_89.Q ;
  assign g6082 = \DFF_1321.Q ;
  assign g6088 = \DFF_97.Q ;
  assign g6093 = \DFF_998.Q ;
  assign g6098 = \DFF_838.Q ;
  assign g6105 = \DFF_879.Q ;
  assign g6109 = \DFF_821.Q ;
  assign g6113 = \DFF_596.Q ;
  assign g6116 = \DFF_1142.Q ;
  assign g6120 = \DFF_1287.Q ;
  assign g6128 = \DFF_344.Q ;
  assign g613 = \DFF_812.Q ;
  assign g6133 = \DFF_978.Q ;
  assign g6137 = \DFF_138.Q ;
  assign g6140 = \DFF_1316.Q ;
  assign g6144 = \DFF_86.Q ;
  assign g6148 = \DFF_377.Q ;
  assign g6151 = \DFF_553.Q ;
  assign g6154 = \DFF_170.Q ;
  assign g6159 = \DFF_300.Q ;
  assign g6163 = \DFF_1203.Q ;
  assign g6167 = \DFF_400.Q ;
  assign g617 = \DFF_751.Q ;
  assign g6173 = \DFF_897.Q ;
  assign g6177 = \DFF_52.Q ;
  assign g6181 = \DFF_1004.Q ;
  assign g6187 = \DFF_275.Q ;
  assign g6191 = \DFF_287.Q ;
  assign g6195 = \DFF_136.Q ;
  assign g6199 = \DFF_64.Q ;
  assign g6203 = \DFF_925.Q ;
  assign g6209 = \DFF_653.Q ;
  assign g6215 = \DFF_104.Q ;
  assign g6219 = \DFF_20.Q ;
  assign g622 = \DFF_119.Q ;
  assign g6227 = \DFF_916.Q ;
  assign g6235 = \DFF_579.Q ;
  assign g6239 = \DFF_494.Q ;
  assign g6243 = \DFF_337.Q ;
  assign g6247 = \DFF_945.Q ;
  assign g6251 = \DFF_314.Q ;
  assign g6255 = \DFF_158.Q ;
  assign g6259 = \DFF_92.Q ;
  assign g626 = \DFF_844.Q ;
  assign g6263 = \DFF_1011.Q ;
  assign g6267 = \DFF_179.Q ;
  assign g6271 = \DFF_634.Q ;
  assign g6275 = \DFF_483.Q ;
  assign g6279 = \DFF_397.Q ;
  assign g6283 = \DFF_904.Q ;
  assign g6287 = \DFF_59.Q ;
  assign g6291 = \DFF_82.Q ;
  assign g6295 = \DFF_1366.Q ;
  assign g6299 = \DFF_1307.Q ;
  assign g63 = \DFF_796.Q ;
  assign g6303 = \DFF_1123.Q ;
  assign g6307 = \DFF_298.Q ;
  assign g6311 = \DFF_484.Q ;
  assign g6315 = \DFF_315.Q ;
  assign g632 = \DFF_338.Q ;
  assign g6322 = \DFF_123.Q ;
  assign g6329 = \DFF_188.Q ;
  assign g6336 = \DFF_118.Q ;
  assign g6346 = \DFF_1119.Q ;
  assign g6351 = \DFF_554.Q ;
  assign g6358 = \DFF_474.Q ;
  assign g6365 = \DFF_970.Q ;
  assign g6369 = \DFF_905.Q ;
  assign g637 = \DFF_752.Q ;
  assign g6373 = \DFF_898.Q ;
  assign g6377 = \DFF_53.Q ;
  assign g6381 = \DFF_1005.Q ;
  assign g6386 = \DFF_251.Q ;
  assign g6390 = \DFF_1188.Q ;
  assign g6395 = \DFF_139.Q ;
  assign g6398 = \DFF_230.Q ;
  assign g640 = \DFF_109.Q ;
  assign g6404 = \DFF_1279.Q ;
  assign g6411 = \DFF_1056.Q ;
  assign g6415 = \DFF_915.Q ;
  assign g6419 = \DFF_850.Q ;
  assign g6423 = \DFF_1105.Q ;
  assign g6428 = \DFF_940.Q ;
  assign g6434 = \DFF_1147.Q ;
  assign g6439 = \DFF_1257.Q ;
  assign g6444 = \DFF_732.Q ;
  assign g645 = \DFF_1042.Q ;
  assign g6451 = \DFF_1113.Q ;
  assign g6455 = \DFF_975.Q ;
  assign g6459 = \DFF_907.Q ;
  assign g6462 = \DFF_3.Q ;
  assign g6466 = \DFF_969.Q ;
  assign g6474 = \DFF_1062.Q ;
  assign g6479 = \DFF_1183.Q ;
  assign g6483 = \DFF_266.Q ;
  assign g6486 = \DFF_861.Q ;
  assign g6490 = \DFF_371.Q ;
  assign g6494 = \DFF_603.Q ;
  assign g6497 = \DFF_168.Q ;
  assign g65 = \DFF_961.Q ;
  assign g650 = \DFF_1126.Q ;
  assign g6500 = \DFF_694.Q ;
  assign g6505 = \DFF_1055.Q ;
  assign g6509 = \DFF_987.Q ;
  assign g6513 = \DFF_755.Q ;
  assign g6519 = \DFF_433.Q ;
  assign g6523 = \DFF_716.Q ;
  assign g6527 = \DFF_1278.Q ;
  assign g6533 = \DFF_1154.Q ;
  assign g6537 = \DFF_332.Q ;
  assign g6541 = \DFF_644.Q ;
  assign g6545 = \DFF_498.Q ;
  assign g6549 = \DFF_410.Q ;
  assign g655 = \DFF_656.Q ;
  assign g6555 = \DFF_584.Q ;
  assign g6561 = \DFF_1273.Q ;
  assign g6565 = \DFF_1150.Q ;
  assign g6573 = \DFF_1068.Q ;
  assign g6581 = \DFF_1174.Q ;
  assign g6585 = \DFF_1032.Q ;
  assign g6589 = \DFF_967.Q ;
  assign g6593 = \DFF_610.Q ;
  assign g6597 = \DFF_1175.Q ;
  assign g66 = \DFF_934.Q ;
  assign g6601 = \DFF_1169.Q ;
  assign g6605 = \DFF_1024.Q ;
  assign g6609 = \DFF_957.Q ;
  assign g661 = \DFF_573.Q ;
  assign g6613 = \DFF_730.Q ;
  assign g6617 = \DFF_1294.Q ;
  assign g6621 = \DFF_588.Q ;
  assign g6625 = \DFF_419.Q ;
  assign g6629 = \DFF_345.Q ;
  assign g6633 = \DFF_1120.Q ;
  assign g6637 = \DFF_291.Q ;
  assign g6641 = \DFF_617.Q ;
  assign g6645 = \DFF_464.Q ;
  assign g6649 = \DFF_378.Q ;
  assign g6653 = \DFF_779.Q ;
  assign g6657 = \DFF_1348.Q ;
  assign g6661 = \DFF_1248.Q ;
  assign g6668 = \DFF_1185.Q ;
  assign g667 = \DFF_866.Q ;
  assign g6675 = \DFF_806.Q ;
  assign g6682 = \DFF_878.Q ;
  assign g6692 = \DFF_163.Q ;
  assign g6697 = \DFF_1158.Q ;
  assign g6704 = \DFF_1196.Q ;
  assign g671 = \DFF_902.Q ;
  assign g6711 = \DFF_971.Q ;
  assign g6715 = \DFF_836.Q ;
  assign g6719 = \DFF_780.Q ;
  assign g6723 = \DFF_1023.Q ;
  assign g6727 = \DFF_198.Q ;
  assign g6732 = \DFF_1130.Q ;
  assign g6736 = \DFF_683.Q ;
  assign g6741 = \DFF_952.Q ;
  assign g6754 = \DFF_1411.Q ;
  assign g6755 = \DFF_1411.Q ;
  assign g6756 = \DFF_790.Q ;
  assign g676 = \DFF_112.Q ;
  assign g6767 = \DFF_512.Q ;
  assign g6772 = \DFF_1229.Q ;
  assign g6782 = \DFF_355.Q ;
  assign g6789 = \DFF_547.Q ;
  assign g681 = \DFF_238.Q ;
  assign g6821 = \DFF_343.Q ;
  assign g6832 = \DFF_395.Q ;
  assign g6856 = \DFF_428.Q ;
  assign g686 = \DFF_900.Q ;
  assign g6867 = \DFF_125.Q ;
  assign g6868 = \DFF_650.Q ;
  assign g6869 = g36;
  assign g6875 = \DFF_1347.Q ;
  assign g6888 = \DFF_282.Q ;
  assign g6905 = \DFF_1312.Q ;
  assign g691 = \DFF_1390.Q ;
  assign g6928 = \DFF_286.Q ;
  assign g6946 = \DFF_1230.Q ;
  assign g6955 = \DFF_210.Q ;
  assign g6961 = \DFF_1016.Q ;
  assign g6971 = \DFF_549.Q ;
  assign g6972 = \DFF_1345.Q ;
  assign g6973 = \DFF_491.Q ;
  assign g6974 = \DFF_1362.Q ;
  assign g6976 = \DFF_615.Q ;
  assign g6977 = \DFF_129.Q ;
  assign g699 = \DFF_1250.Q ;
  assign g7 = \DFF_1222.Q ;
  assign g70 = \DFF_650.Q ;
  assign g7004 = \DFF_846.Q ;
  assign g7028 = \DFF_1252.Q ;
  assign g703 = \DFF_667.Q ;
  assign g7051 = \DFF_833.Q ;
  assign g7074 = \DFF_139.Q ;
  assign g7097 = \DFF_952.Q ;
  assign g71 = \DFF_1424.Q ;
  assign g7117 = \DFF_743.Q ;
  assign g7121 = \DFF_473.Q ;
  assign g714 = \DFF_1019.Q ;
  assign g7148 = \DFF_417.Q ;
  assign g7161 = \DFF_1220.Q ;
  assign g718 = \DFF_135.Q ;
  assign g7196 = \DFF_304.Q ;
  assign g723 = \DFF_1251.Q ;
  assign g7231 = g12833;
  assign g7243 = \DFF_1073.Q ;
  assign g7245 = \DFF_1225.Q ;
  assign g7257 = \DFF_234.Q ;
  assign g7260 = \DFF_348.Q ;
  assign g728 = \DFF_1365.Q ;
  assign g732 = \DFF_988.Q ;
  assign g736 = \DFF_256.Q ;
  assign g739 = \DFF_876.Q ;
  assign g74 = \DFF_654.Q ;
  assign g744 = \DFF_175.Q ;
  assign g7474 = \DFF_934.Q ;
  assign g749 = \DFF_28.Q ;
  assign g7502 = \DFF_157.Q ;
  assign g7515 = \DFF_1235.Q ;
  assign g7516 = \DFF_74.Q ;
  assign g7526 = \DFF_162.Q ;
  assign g7527 = \DFF_50.Q ;
  assign g753 = \DFF_194.Q ;
  assign g7540 = \DFF_686.Q ;
  assign g7542 = \DFF_1090.Q ;
  assign g7543 = \DFF_789.Q ;
  assign g7558 = \DFF_1080.Q ;
  assign g7565 = \DFF_812.Q ;
  assign g7566 = \DFF_896.Q ;
  assign g758 = \DFF_328.Q ;
  assign g7586 = \DFF_1020.Q ;
  assign g7593 = \DFF_88.Q ;
  assign g7594 = \DFF_751.Q ;
  assign g7595 = \DFF_876.Q ;
  assign g7596 = \DFF_953.Q ;
  assign g7615 = \DFF_728.Q ;
  assign g7616 = \DFF_119.Q ;
  assign g7617 = \DFF_175.Q ;
  assign g7618 = \DFF_1200.Q ;
  assign g7623 = \DFF_506.Q ;
  assign g7624 = \DFF_844.Q ;
  assign g7625 = \DFF_28.Q ;
  assign g7626 = \DFF_661.Q ;
  assign g763 = \DFF_157.Q ;
  assign g7632 = \DFF_560.Q ;
  assign g7633 = \DFF_338.Q ;
  assign g7634 = \DFF_328.Q ;
  assign g7640 = \DFF_1340.Q ;
  assign g7647 = \DFF_863.Q ;
  assign g7648 = \DFF_21.Q ;
  assign g7659 = \DFF_874.Q ;
  assign g7660 = \DFF_142.Q ;
  assign g767 = \DFF_74.Q ;
  assign g7674 = \DFF_966.Q ;
  assign g7689 = \DFF_89.Q ;
  assign g7704 = \DFF_1098.Q ;
  assign g7717 = \DFF_962.Q ;
  assign g772 = \DFF_50.Q ;
  assign g7738 = \DFF_289.Q ;
  assign g7753 = \DFF_893.Q ;
  assign g776 = \DFF_789.Q ;
  assign g7766 = \DFF_393.Q ;
  assign g7791 = \DFF_104.Q ;
  assign g781 = \DFF_896.Q ;
  assign g7812 = \DFF_1273.Q ;
  assign g7831 = \DFF_1074.Q ;
  assign g785 = \DFF_953.Q ;
  assign g79 = \DFF_1044.Q ;
  assign g790 = \DFF_1200.Q ;
  assign g7916 = \DFF_675.Q ;
  assign g794 = \DFF_661.Q ;
  assign g7946 = \DFF_60.Q ;
  assign g799 = \DFF_515.Q ;
  assign g7993 = \DFF_514.Q ;
  assign g7994 = \DFF_206.Q ;
  assign g8 = \DFF_761.Q ;
  assign g802 = \DFF_1081.Q ;
  assign g8032 = \DFF_477.Q ;
  assign g8038 = \DFF_353.Q ;
  assign g807 = \DFF_21.Q ;
  assign g8085 = \DFF_829.Q ;
  assign g812 = \DFF_524.Q ;
  assign g8132 = \DFF_178.Q ;
  assign g8134 = \DFF_150.Q ;
  assign g8135 = \DFF_621.Q ;
  assign g817 = \DFF_870.Q ;
  assign g8178 = \DFF_672.Q ;
  assign g8215 = \DFF_317.Q ;
  assign g822 = \DFF_278.Q ;
  assign g8235 = \DFF_997.Q ;
  assign g827 = \DFF_710.Q ;
  assign g8277 = \DFF_1256.Q ;
  assign g8279 = \DFF_830.Q ;
  assign g8283 = \DFF_981.Q ;
  assign g8285 = \DFF_1322.Q ;
  assign g8291 = \DFF_612.Q ;
  assign g832 = \DFF_525.Q ;
  assign g8342 = \DFF_1414.Q ;
  assign g8344 = \DFF_147.Q ;
  assign g8353 = \DFF_1118.Q ;
  assign g8355 = \DFF_1012.Q ;
  assign g8358 = \DFF_824.Q ;
  assign g837 = \DFF_872.Q ;
  assign g8398 = \DFF_460.Q ;
  assign g8403 = \DFF_1100.Q ;
  assign g8405 = \DFF_420.Q ;
  assign g8411 = \DFF_339.Q ;
  assign g8416 = \DFF_1308.Q ;
  assign g843 = \DFF_113.Q ;
  assign g847 = \DFF_23.Q ;
  assign g8470 = \DFF_1275.Q ;
  assign g8475 = \DFF_334.Q ;
  assign g8481 = \DFF_538.Q ;
  assign g85 = \DFF_1111.Q ;
  assign g8515 = \DFF_828.Q ;
  assign g854 = \DFF_719.Q ;
  assign g8542 = \DFF_664.Q ;
  assign g8572 = \DFF_481.Q ;
  assign g859 = \DFF_585.Q ;
  assign g8595 = \DFF_5.Q ;
  assign g86 = \DFF_1078.Q ;
  assign g8607 = g23002;
  assign g862 = \DFF_669.Q ;
  assign g869 = \DFF_561.Q ;
  assign g8703 = \DFF_1384.Q ;
  assign g8712 = \DFF_1425.Q ;
  assign g8719 = \DFF_269.Q ;
  assign g872 = \DFF_1003.Q ;
  assign g8740 = \DFF_221.Q ;
  assign g875 = \DFF_1106.Q ;
  assign g8757 = \DFF_411.Q ;
  assign g8763 = \DFF_350.Q ;
  assign g8778 = \DFF_551.Q ;
  assign g878 = \DFF_152.Q ;
  assign g8783 = \DFF_480.Q ;
  assign g8784 = \DFF_909.Q ;
  assign g8785 = \DFF_565.Q ;
  assign g8786 = \DFF_1224.Q ;
  assign g8787 = \DFF_1416.Q ;
  assign g8788 = \DFF_1049.Q ;
  assign g8789 = \DFF_704.Q ;
  assign g8791 = \DFF_1379.Q ;
  assign g8792 = \DFF_853.Q ;
  assign g8795 = \DFF_439.Q ;
  assign g8805 = \DFF_1425.Q ;
  assign g881 = \DFF_404.Q ;
  assign g8812 = \DFF_351.Q ;
  assign g8818 = \DFF_1084.Q ;
  assign g8821 = \DFF_853.Q ;
  assign g8839 = \DFF_831.Q ;
  assign g884 = \DFF_380.Q ;
  assign g8841 = \DFF_1379.Q ;
  assign g8844 = \DFF_1173.Q ;
  assign g887 = \DFF_764.Q ;
  assign g8870 = \DFF_885.Q ;
  assign g8876 = \DFF_1379.Q ;
  assign g8879 = \DFF_853.Q ;
  assign g8880 = \DFF_26.Q ;
  assign g890 = \DFF_736.Q ;
  assign g8915 = \DFF_1286.Q ;
  assign g8916 = \DFF_485.Q ;
  assign g8917 = \DFF_992.Q ;
  assign g8918 = \DFF_418.Q ;
  assign g8919 = \DFF_944.Q ;
  assign g8920 = \DFF_1338.Q ;
  assign g8922 = \DFF_1084.Q ;
  assign g8925 = \DFF_853.Q ;
  assign g896 = \DFF_799.Q ;
  assign g8971 = \DFF_115.Q ;
  assign g8974 = \DFF_1173.Q ;
  assign g8989 = g6753;
  assign g9 = \DFF_547.Q ;
  assign g901 = \DFF_908.Q ;
  assign g9019 = \DFF_1027.Q ;
  assign g9021 = \DFF_1374.Q ;
  assign g904 = \DFF_880.Q ;
  assign g9048 = \DFF_109.Q ;
  assign g907 = \DFF_1241.Q ;
  assign g9071 = g23759;
  assign g911 = \DFF_303.Q ;
  assign g914 = \DFF_280.Q ;
  assign g9152 = g23652;
  assign g9153 = g6752;
  assign g9154 = g6748;
  assign g9155 = \DFF_240.Q ;
  assign g918 = \DFF_859.Q ;
  assign g9185 = \DFF_961.Q ;
  assign g9186 = g6749;
  assign g921 = \DFF_94.Q ;
  assign g9213 = g6750;
  assign g9245 = g6747;
  assign g925 = \DFF_149.Q ;
  assign g9251 = \DFF_203.Q ;
  assign g9280 = g6744;
  assign g9281 = \DFF_1181.Q ;
  assign g929 = \DFF_1353.Q ;
  assign g93 = \DFF_743.Q ;
  assign g930 = \DFF_867.Q ;
  assign g933 = \DFF_758.Q ;
  assign g9340 = \DFF_746.Q ;
  assign g936 = \DFF_963.Q ;
  assign g939 = \DFF_127.Q ;
  assign g94 = \DFF_1301.Q ;
  assign g9417 = \DFF_845.Q ;
  assign g943 = \DFF_1314.Q ;
  assign g947 = \DFF_1242.Q ;
  assign g9477 = g6745;
  assign g9478 = g6746;
  assign g9497 = \DFF_678.Q ;
  assign g952 = \DFF_453.Q ;
  assign g9553 = \DFF_545.Q ;
  assign g9555 = \DFF_630.Q ;
  assign g956 = \DFF_1136.Q ;
  assign g9615 = \DFF_503.Q ;
  assign g9617 = \DFF_85.Q ;
  assign g962 = \DFF_416.Q ;
  assign g9637 = g6751;
  assign g967 = \DFF_800.Q ;
  assign g968 = \DFF_999.Q ;
  assign g9680 = \DFF_376.Q ;
  assign g9682 = \DFF_1316.Q ;
  assign g9687 = \DFF_379.Q ;
  assign g969 = \DFF_283.Q ;
  assign g9741 = \DFF_86.Q ;
  assign g9743 = \DFF_861.Q ;
  assign g9746 = \DFF_934.Q ;
  assign g9747 = \DFF_1078.Q ;
  assign g976 = \DFF_24.Q ;
  assign g9772 = \DFF_673.Q ;
  assign g9780 = \DFF_141.Q ;
  assign g979 = \DFF_698.Q ;
  assign g9817 = \DFF_371.Q ;
  assign g9864 = \DFF_599.Q ;
  assign g990 = \DFF_511.Q ;
  assign g9917 = \DFF_767.Q ;
  assign g9935 = \DFF_1320.Q ;
  assign g996 = \DFF_606.Q ;
endmodule
