
module c499(N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  input N1;
  input N101;
  input N105;
  input N109;
  input N113;
  input N117;
  input N121;
  input N125;
  input N129;
  input N13;
  input N130;
  input N131;
  input N132;
  input N133;
  input N134;
  input N135;
  input N136;
  input N137;
  input N17;
  input N21;
  input N25;
  input N29;
  input N33;
  input N37;
  input N41;
  input N45;
  input N49;
  input N5;
  input N53;
  input N57;
  input N61;
  input N65;
  input N69;
  output N724;
  output N725;
  output N726;
  output N727;
  output N728;
  output N729;
  input N73;
  output N730;
  output N731;
  output N732;
  output N733;
  output N734;
  output N735;
  output N736;
  output N737;
  output N738;
  output N739;
  output N740;
  output N741;
  output N742;
  output N743;
  output N744;
  output N745;
  output N746;
  output N747;
  output N748;
  output N749;
  output N750;
  output N751;
  output N752;
  output N753;
  output N754;
  output N755;
  input N77;
  input N81;
  input N85;
  input N89;
  input N9;
  input N93;
  input N97;
  al_inv _332_ (
    .a(N1),
    .y(_306_)
  );
  al_nand2 _333_ (
    .a(N33),
    .b(N49),
    .y(_307_)
  );
  al_nor2 _334_ (
    .a(N33),
    .b(N49),
    .y(_308_)
  );
  al_nand2ft _335_ (
    .a(_308_),
    .b(_307_),
    .y(_309_)
  );
  al_nand2 _336_ (
    .a(N129),
    .b(N137),
    .y(_310_)
  );
  al_nand2 _337_ (
    .a(N1),
    .b(N17),
    .y(_311_)
  );
  al_or2 _338_ (
    .a(N1),
    .b(N17),
    .y(_312_)
  );
  al_ao21 _339_ (
    .a(_312_),
    .b(_311_),
    .c(_310_),
    .y(_313_)
  );
  al_nand3 _340_ (
    .a(_312_),
    .b(_310_),
    .c(_311_),
    .y(_314_)
  );
  al_nand3 _341_ (
    .a(_313_),
    .b(_309_),
    .c(_314_),
    .y(_315_)
  );
  al_aoi21 _342_ (
    .a(_313_),
    .b(_314_),
    .c(_309_),
    .y(_316_)
  );
  al_nand2ft _343_ (
    .a(_316_),
    .b(_315_),
    .y(_317_)
  );
  al_and2ft _344_ (
    .a(N73),
    .b(N77),
    .y(_318_)
  );
  al_nand2ft _345_ (
    .a(N77),
    .b(N73),
    .y(_319_)
  );
  al_and2ft _346_ (
    .a(N69),
    .b(N65),
    .y(_320_)
  );
  al_nand2ft _347_ (
    .a(N65),
    .b(N69),
    .y(_321_)
  );
  al_nand2ft _348_ (
    .a(_320_),
    .b(_321_),
    .y(_322_)
  );
  al_and3fft _349_ (
    .a(_318_),
    .b(_322_),
    .c(_319_),
    .y(_323_)
  );
  al_aoi21ftf _350_ (
    .a(_318_),
    .b(_319_),
    .c(_322_),
    .y(_324_)
  );
  al_or2 _351_ (
    .a(_324_),
    .b(_323_),
    .y(_325_)
  );
  al_and2ft _352_ (
    .a(N89),
    .b(N93),
    .y(_326_)
  );
  al_nand2ft _353_ (
    .a(N93),
    .b(N89),
    .y(_327_)
  );
  al_and2ft _354_ (
    .a(N85),
    .b(N81),
    .y(_328_)
  );
  al_nand2ft _355_ (
    .a(N81),
    .b(N85),
    .y(_329_)
  );
  al_nand2ft _356_ (
    .a(_328_),
    .b(_329_),
    .y(_330_)
  );
  al_or3ftt _357_ (
    .a(_327_),
    .b(_326_),
    .c(_330_),
    .y(_331_)
  );
  al_ao21ftf _358_ (
    .a(_326_),
    .b(_327_),
    .c(_330_),
    .y(_000_)
  );
  al_or3fft _359_ (
    .a(_331_),
    .b(_000_),
    .c(_325_),
    .y(_001_)
  );
  al_nand3ftt _360_ (
    .a(_326_),
    .b(_327_),
    .c(_330_),
    .y(_002_)
  );
  al_ao21ftt _361_ (
    .a(_326_),
    .b(_327_),
    .c(_330_),
    .y(_003_)
  );
  al_nand3 _362_ (
    .a(_002_),
    .b(_003_),
    .c(_325_),
    .y(_004_)
  );
  al_and3 _363_ (
    .a(_317_),
    .b(_004_),
    .c(_001_),
    .y(_005_)
  );
  al_nand3 _364_ (
    .a(_331_),
    .b(_000_),
    .c(_325_),
    .y(_006_)
  );
  al_or3fft _365_ (
    .a(_002_),
    .b(_003_),
    .c(_325_),
    .y(_007_)
  );
  al_nand3ftt _366_ (
    .a(_317_),
    .b(_006_),
    .c(_007_),
    .y(_008_)
  );
  al_nand2ft _367_ (
    .a(_005_),
    .b(_008_),
    .y(_009_)
  );
  al_nand2 _368_ (
    .a(N137),
    .b(N133),
    .y(_010_)
  );
  al_nand2 _369_ (
    .a(N97),
    .b(N113),
    .y(_011_)
  );
  al_nor2 _370_ (
    .a(N97),
    .b(N113),
    .y(_012_)
  );
  al_nand2ft _371_ (
    .a(_012_),
    .b(_011_),
    .y(_013_)
  );
  al_nand2 _372_ (
    .a(N65),
    .b(N81),
    .y(_014_)
  );
  al_or2 _373_ (
    .a(N65),
    .b(N81),
    .y(_015_)
  );
  al_nand3 _374_ (
    .a(_014_),
    .b(_015_),
    .c(_013_),
    .y(_016_)
  );
  al_ao21 _375_ (
    .a(_014_),
    .b(_015_),
    .c(_013_),
    .y(_017_)
  );
  al_ao21 _376_ (
    .a(_016_),
    .b(_017_),
    .c(_010_),
    .y(_018_)
  );
  al_and3 _377_ (
    .a(_010_),
    .b(_016_),
    .c(_017_),
    .y(_019_)
  );
  al_and2ft _378_ (
    .a(_019_),
    .b(_018_),
    .y(_020_)
  );
  al_and2ft _379_ (
    .a(N9),
    .b(N13),
    .y(_021_)
  );
  al_nand2ft _380_ (
    .a(N13),
    .b(N9),
    .y(_022_)
  );
  al_nand2 _381_ (
    .a(N1),
    .b(N5),
    .y(_023_)
  );
  al_nor2 _382_ (
    .a(N1),
    .b(N5),
    .y(_024_)
  );
  al_nand2ft _383_ (
    .a(_024_),
    .b(_023_),
    .y(_025_)
  );
  al_and3ftt _384_ (
    .a(_021_),
    .b(_022_),
    .c(_025_),
    .y(_026_)
  );
  al_aoi21ftt _385_ (
    .a(_021_),
    .b(_022_),
    .c(_025_),
    .y(_027_)
  );
  al_or2 _386_ (
    .a(_026_),
    .b(_027_),
    .y(_028_)
  );
  al_and2ft _387_ (
    .a(N25),
    .b(N29),
    .y(_029_)
  );
  al_nand2ft _388_ (
    .a(N29),
    .b(N25),
    .y(_030_)
  );
  al_and2ft _389_ (
    .a(N21),
    .b(N17),
    .y(_031_)
  );
  al_nand2ft _390_ (
    .a(N17),
    .b(N21),
    .y(_032_)
  );
  al_nand2ft _391_ (
    .a(_031_),
    .b(_032_),
    .y(_033_)
  );
  al_and3ftt _392_ (
    .a(_029_),
    .b(_030_),
    .c(_033_),
    .y(_034_)
  );
  al_aoi21ftt _393_ (
    .a(_029_),
    .b(_030_),
    .c(_033_),
    .y(_035_)
  );
  al_or3 _394_ (
    .a(_034_),
    .b(_035_),
    .c(_028_),
    .y(_036_)
  );
  al_or3ftt _395_ (
    .a(_030_),
    .b(_029_),
    .c(_033_),
    .y(_037_)
  );
  al_aoi21ftf _396_ (
    .a(_029_),
    .b(_030_),
    .c(_033_),
    .y(_038_)
  );
  al_and3ftt _397_ (
    .a(_038_),
    .b(_037_),
    .c(_028_),
    .y(_039_)
  );
  al_oa21ftf _398_ (
    .a(_036_),
    .b(_039_),
    .c(_020_),
    .y(_040_)
  );
  al_nand3ftt _399_ (
    .a(_039_),
    .b(_020_),
    .c(_036_),
    .y(_041_)
  );
  al_nand2 _400_ (
    .a(N101),
    .b(N117),
    .y(_042_)
  );
  al_nor2 _401_ (
    .a(N101),
    .b(N117),
    .y(_043_)
  );
  al_nand2ft _402_ (
    .a(_043_),
    .b(_042_),
    .y(_044_)
  );
  al_nand2 _403_ (
    .a(N137),
    .b(N134),
    .y(_045_)
  );
  al_nand2 _404_ (
    .a(N69),
    .b(N85),
    .y(_046_)
  );
  al_or2 _405_ (
    .a(N69),
    .b(N85),
    .y(_047_)
  );
  al_ao21 _406_ (
    .a(_047_),
    .b(_046_),
    .c(_045_),
    .y(_048_)
  );
  al_nand3 _407_ (
    .a(_047_),
    .b(_045_),
    .c(_046_),
    .y(_049_)
  );
  al_nand3 _408_ (
    .a(_048_),
    .b(_044_),
    .c(_049_),
    .y(_050_)
  );
  al_aoi21 _409_ (
    .a(_048_),
    .b(_049_),
    .c(_044_),
    .y(_051_)
  );
  al_nand2ft _410_ (
    .a(_051_),
    .b(_050_),
    .y(_052_)
  );
  al_and2ft _411_ (
    .a(N41),
    .b(N45),
    .y(_053_)
  );
  al_nand2ft _412_ (
    .a(N45),
    .b(N41),
    .y(_054_)
  );
  al_nand2ft _413_ (
    .a(_053_),
    .b(_054_),
    .y(_055_)
  );
  al_nand2ft _414_ (
    .a(N37),
    .b(N33),
    .y(_056_)
  );
  al_nand2ft _415_ (
    .a(N33),
    .b(N37),
    .y(_057_)
  );
  al_aoi21 _416_ (
    .a(_056_),
    .b(_057_),
    .c(_055_),
    .y(_058_)
  );
  al_nand3 _417_ (
    .a(_056_),
    .b(_057_),
    .c(_055_),
    .y(_059_)
  );
  al_or2ft _418_ (
    .a(_059_),
    .b(_058_),
    .y(_060_)
  );
  al_nand2ft _419_ (
    .a(N57),
    .b(N61),
    .y(_061_)
  );
  al_nand2ft _420_ (
    .a(N61),
    .b(N57),
    .y(_062_)
  );
  al_and2ft _421_ (
    .a(N53),
    .b(N49),
    .y(_063_)
  );
  al_nand2ft _422_ (
    .a(N49),
    .b(N53),
    .y(_064_)
  );
  al_nand2ft _423_ (
    .a(_063_),
    .b(_064_),
    .y(_065_)
  );
  al_and3 _424_ (
    .a(_061_),
    .b(_062_),
    .c(_065_),
    .y(_066_)
  );
  al_and2ft _425_ (
    .a(N57),
    .b(N61),
    .y(_067_)
  );
  al_nand2ft _426_ (
    .a(_067_),
    .b(_062_),
    .y(_068_)
  );
  al_nand3ftt _427_ (
    .a(_063_),
    .b(_064_),
    .c(_068_),
    .y(_069_)
  );
  al_nand3ftt _428_ (
    .a(_066_),
    .b(_069_),
    .c(_060_),
    .y(_070_)
  );
  al_nand2ft _429_ (
    .a(_066_),
    .b(_069_),
    .y(_071_)
  );
  al_nand3ftt _430_ (
    .a(_058_),
    .b(_059_),
    .c(_071_),
    .y(_072_)
  );
  al_aoi21 _431_ (
    .a(_072_),
    .b(_070_),
    .c(_052_),
    .y(_073_)
  );
  al_nand3 _432_ (
    .a(_052_),
    .b(_072_),
    .c(_070_),
    .y(_074_)
  );
  al_or2ft _433_ (
    .a(_074_),
    .b(_073_),
    .y(_075_)
  );
  al_aoi21ftf _434_ (
    .a(_040_),
    .b(_041_),
    .c(_075_),
    .y(_076_)
  );
  al_and2 _435_ (
    .a(N137),
    .b(N135),
    .y(_077_)
  );
  al_nand2 _436_ (
    .a(N105),
    .b(N121),
    .y(_078_)
  );
  al_nor2 _437_ (
    .a(N105),
    .b(N121),
    .y(_079_)
  );
  al_nand2ft _438_ (
    .a(_079_),
    .b(_078_),
    .y(_080_)
  );
  al_nand2 _439_ (
    .a(N73),
    .b(N89),
    .y(_081_)
  );
  al_or2 _440_ (
    .a(N73),
    .b(N89),
    .y(_082_)
  );
  al_nand3 _441_ (
    .a(_081_),
    .b(_082_),
    .c(_080_),
    .y(_083_)
  );
  al_ao21 _442_ (
    .a(_081_),
    .b(_082_),
    .c(_080_),
    .y(_084_)
  );
  al_ao21 _443_ (
    .a(_083_),
    .b(_084_),
    .c(_077_),
    .y(_085_)
  );
  al_and3 _444_ (
    .a(_077_),
    .b(_083_),
    .c(_084_),
    .y(_086_)
  );
  al_nand2ft _445_ (
    .a(_086_),
    .b(_085_),
    .y(_087_)
  );
  al_ao21ftf _446_ (
    .a(_058_),
    .b(_059_),
    .c(_028_),
    .y(_088_)
  );
  al_or3 _447_ (
    .a(_026_),
    .b(_027_),
    .c(_060_),
    .y(_089_)
  );
  al_or3fft _448_ (
    .a(_088_),
    .b(_089_),
    .c(_087_),
    .y(_090_)
  );
  al_ao21ttf _449_ (
    .a(_088_),
    .b(_089_),
    .c(_087_),
    .y(_091_)
  );
  al_nand2 _450_ (
    .a(N109),
    .b(N125),
    .y(_092_)
  );
  al_nor2 _451_ (
    .a(N109),
    .b(N125),
    .y(_093_)
  );
  al_nand2ft _452_ (
    .a(_093_),
    .b(_092_),
    .y(_094_)
  );
  al_nand2 _453_ (
    .a(N137),
    .b(N136),
    .y(_095_)
  );
  al_nand2 _454_ (
    .a(N77),
    .b(N93),
    .y(_096_)
  );
  al_or2 _455_ (
    .a(N77),
    .b(N93),
    .y(_097_)
  );
  al_ao21 _456_ (
    .a(_097_),
    .b(_096_),
    .c(_095_),
    .y(_098_)
  );
  al_nand3 _457_ (
    .a(_097_),
    .b(_095_),
    .c(_096_),
    .y(_099_)
  );
  al_nand3 _458_ (
    .a(_098_),
    .b(_094_),
    .c(_099_),
    .y(_100_)
  );
  al_aoi21 _459_ (
    .a(_098_),
    .b(_099_),
    .c(_094_),
    .y(_101_)
  );
  al_nand2ft _460_ (
    .a(_101_),
    .b(_100_),
    .y(_102_)
  );
  al_nand3fft _461_ (
    .a(_034_),
    .b(_035_),
    .c(_071_),
    .y(_103_)
  );
  al_or3fft _462_ (
    .a(_061_),
    .b(_062_),
    .c(_065_),
    .y(_104_)
  );
  al_aoi21ftf _463_ (
    .a(_067_),
    .b(_062_),
    .c(_065_),
    .y(_105_)
  );
  al_nand2ft _464_ (
    .a(_105_),
    .b(_104_),
    .y(_106_)
  );
  al_and3ftt _465_ (
    .a(_038_),
    .b(_037_),
    .c(_106_),
    .y(_107_)
  );
  al_nor3fft _466_ (
    .a(_102_),
    .b(_103_),
    .c(_107_),
    .y(_108_)
  );
  al_oai21ftf _467_ (
    .a(_103_),
    .b(_107_),
    .c(_102_),
    .y(_109_)
  );
  al_nand2ft _468_ (
    .a(_108_),
    .b(_109_),
    .y(_110_)
  );
  al_and3 _469_ (
    .a(_090_),
    .b(_091_),
    .c(_110_),
    .y(_111_)
  );
  al_ao21ftf _470_ (
    .a(_318_),
    .b(_319_),
    .c(_322_),
    .y(_112_)
  );
  al_and2 _471_ (
    .a(N137),
    .b(N131),
    .y(_113_)
  );
  al_nor3fft _472_ (
    .a(_113_),
    .b(_112_),
    .c(_323_),
    .y(_114_)
  );
  al_oai21ftf _473_ (
    .a(_112_),
    .b(_323_),
    .c(_113_),
    .y(_115_)
  );
  al_and2ft _474_ (
    .a(_114_),
    .b(_115_),
    .y(_116_)
  );
  al_and2ft _475_ (
    .a(N105),
    .b(N109),
    .y(_117_)
  );
  al_nand2ft _476_ (
    .a(N109),
    .b(N105),
    .y(_118_)
  );
  al_and2ft _477_ (
    .a(N101),
    .b(N97),
    .y(_119_)
  );
  al_nand2ft _478_ (
    .a(N97),
    .b(N101),
    .y(_120_)
  );
  al_nand2ft _479_ (
    .a(_119_),
    .b(_120_),
    .y(_121_)
  );
  al_and3ftt _480_ (
    .a(_117_),
    .b(_118_),
    .c(_121_),
    .y(_122_)
  );
  al_ao21ftt _481_ (
    .a(_117_),
    .b(_118_),
    .c(_121_),
    .y(_123_)
  );
  al_nand2ft _482_ (
    .a(_122_),
    .b(_123_),
    .y(_124_)
  );
  al_and2ft _483_ (
    .a(N41),
    .b(N57),
    .y(_125_)
  );
  al_nand2ft _484_ (
    .a(N57),
    .b(N41),
    .y(_126_)
  );
  al_nand2ft _485_ (
    .a(_125_),
    .b(_126_),
    .y(_127_)
  );
  al_and2ft _486_ (
    .a(N25),
    .b(N9),
    .y(_128_)
  );
  al_nand2ft _487_ (
    .a(N9),
    .b(N25),
    .y(_129_)
  );
  al_aoi21ftt _488_ (
    .a(_128_),
    .b(_129_),
    .c(_127_),
    .y(_130_)
  );
  al_nand3ftt _489_ (
    .a(_128_),
    .b(_129_),
    .c(_127_),
    .y(_131_)
  );
  al_aoi21ftt _490_ (
    .a(_130_),
    .b(_131_),
    .c(_124_),
    .y(_132_)
  );
  al_nand3ftt _491_ (
    .a(_130_),
    .b(_131_),
    .c(_124_),
    .y(_133_)
  );
  al_nor3fft _492_ (
    .a(_133_),
    .b(_116_),
    .c(_132_),
    .y(_134_)
  );
  al_oa21ftf _493_ (
    .a(_133_),
    .b(_132_),
    .c(_116_),
    .y(_135_)
  );
  al_or2 _494_ (
    .a(_135_),
    .b(_134_),
    .y(_136_)
  );
  al_nand2 _495_ (
    .a(N37),
    .b(N53),
    .y(_137_)
  );
  al_nor2 _496_ (
    .a(N37),
    .b(N53),
    .y(_138_)
  );
  al_nand2ft _497_ (
    .a(_138_),
    .b(_137_),
    .y(_139_)
  );
  al_nand2 _498_ (
    .a(N137),
    .b(N130),
    .y(_140_)
  );
  al_nand2 _499_ (
    .a(N5),
    .b(N21),
    .y(_141_)
  );
  al_or2 _500_ (
    .a(N5),
    .b(N21),
    .y(_142_)
  );
  al_ao21 _501_ (
    .a(_142_),
    .b(_141_),
    .c(_140_),
    .y(_143_)
  );
  al_nand3 _502_ (
    .a(_142_),
    .b(_140_),
    .c(_141_),
    .y(_144_)
  );
  al_nand3 _503_ (
    .a(_143_),
    .b(_139_),
    .c(_144_),
    .y(_145_)
  );
  al_aoi21 _504_ (
    .a(_143_),
    .b(_144_),
    .c(_139_),
    .y(_146_)
  );
  al_nand2ft _505_ (
    .a(_146_),
    .b(_145_),
    .y(_147_)
  );
  al_and2ft _506_ (
    .a(N121),
    .b(N125),
    .y(_148_)
  );
  al_nand2ft _507_ (
    .a(N125),
    .b(N121),
    .y(_149_)
  );
  al_nand2 _508_ (
    .a(N113),
    .b(N117),
    .y(_150_)
  );
  al_nor2 _509_ (
    .a(N113),
    .b(N117),
    .y(_151_)
  );
  al_nand2ft _510_ (
    .a(_151_),
    .b(_150_),
    .y(_152_)
  );
  al_and3ftt _511_ (
    .a(_148_),
    .b(_149_),
    .c(_152_),
    .y(_153_)
  );
  al_aoi21ftt _512_ (
    .a(_148_),
    .b(_149_),
    .c(_152_),
    .y(_154_)
  );
  al_nand3fft _513_ (
    .a(_153_),
    .b(_154_),
    .c(_124_),
    .y(_155_)
  );
  al_or2 _514_ (
    .a(_153_),
    .b(_154_),
    .y(_156_)
  );
  al_and3ftt _515_ (
    .a(_122_),
    .b(_123_),
    .c(_156_),
    .y(_157_)
  );
  al_and3fft _516_ (
    .a(_147_),
    .b(_157_),
    .c(_155_),
    .y(_158_)
  );
  al_oai21ftt _517_ (
    .a(_155_),
    .b(_157_),
    .c(_147_),
    .y(_159_)
  );
  al_nand2ft _518_ (
    .a(_158_),
    .b(_159_),
    .y(_160_)
  );
  al_or3 _519_ (
    .a(_160_),
    .b(_009_),
    .c(_136_),
    .y(_161_)
  );
  al_aoi21ftf _520_ (
    .a(_005_),
    .b(_008_),
    .c(_160_),
    .y(_162_)
  );
  al_ao21ftf _521_ (
    .a(_136_),
    .b(_162_),
    .c(_161_),
    .y(_163_)
  );
  al_and2 _522_ (
    .a(N137),
    .b(N132),
    .y(_164_)
  );
  al_nand3ftt _523_ (
    .a(_164_),
    .b(_000_),
    .c(_331_),
    .y(_165_)
  );
  al_and3 _524_ (
    .a(_164_),
    .b(_002_),
    .c(_003_),
    .y(_166_)
  );
  al_nand2ft _525_ (
    .a(_166_),
    .b(_165_),
    .y(_167_)
  );
  al_and2ft _526_ (
    .a(N45),
    .b(N61),
    .y(_168_)
  );
  al_nand2ft _527_ (
    .a(N61),
    .b(N45),
    .y(_169_)
  );
  al_nand2 _528_ (
    .a(N13),
    .b(N29),
    .y(_170_)
  );
  al_nor2 _529_ (
    .a(N13),
    .b(N29),
    .y(_171_)
  );
  al_and2ft _530_ (
    .a(_171_),
    .b(_170_),
    .y(_172_)
  );
  al_or3ftt _531_ (
    .a(_169_),
    .b(_168_),
    .c(_172_),
    .y(_173_)
  );
  al_ao21ftf _532_ (
    .a(_168_),
    .b(_169_),
    .c(_172_),
    .y(_174_)
  );
  al_nand3 _533_ (
    .a(_173_),
    .b(_174_),
    .c(_156_),
    .y(_175_)
  );
  al_ao21 _534_ (
    .a(_173_),
    .b(_174_),
    .c(_156_),
    .y(_176_)
  );
  al_nand3 _535_ (
    .a(_175_),
    .b(_167_),
    .c(_176_),
    .y(_177_)
  );
  al_aoi21 _536_ (
    .a(_175_),
    .b(_176_),
    .c(_167_),
    .y(_178_)
  );
  al_nand2ft _537_ (
    .a(_178_),
    .b(_177_),
    .y(_179_)
  );
  al_and3ftt _538_ (
    .a(_178_),
    .b(_177_),
    .c(_136_),
    .y(_180_)
  );
  al_nand3fft _539_ (
    .a(_134_),
    .b(_135_),
    .c(_179_),
    .y(_181_)
  );
  al_nand3ftt _540_ (
    .a(_005_),
    .b(_008_),
    .c(_160_),
    .y(_182_)
  );
  al_oai21ftf _541_ (
    .a(_181_),
    .b(_180_),
    .c(_182_),
    .y(_183_)
  );
  al_ao21ftf _542_ (
    .a(_179_),
    .b(_163_),
    .c(_183_),
    .y(_184_)
  );
  al_and3 _543_ (
    .a(_076_),
    .b(_111_),
    .c(_184_),
    .y(_185_)
  );
  al_ao21 _544_ (
    .a(_009_),
    .b(_185_),
    .c(_306_),
    .y(_186_)
  );
  al_and3 _545_ (
    .a(_306_),
    .b(_009_),
    .c(_185_),
    .y(_187_)
  );
  al_nand2ft _546_ (
    .a(_187_),
    .b(_186_),
    .y(N724)
  );
  al_inv _547_ (
    .a(N5),
    .y(_188_)
  );
  al_inv _548_ (
    .a(_160_),
    .y(_189_)
  );
  al_ao21 _549_ (
    .a(_189_),
    .b(_185_),
    .c(_188_),
    .y(_190_)
  );
  al_and3 _550_ (
    .a(_188_),
    .b(_189_),
    .c(_185_),
    .y(_191_)
  );
  al_nand2ft _551_ (
    .a(_191_),
    .b(_190_),
    .y(N725)
  );
  al_inv _552_ (
    .a(N9),
    .y(_192_)
  );
  al_and3 _553_ (
    .a(_192_),
    .b(_136_),
    .c(_185_),
    .y(_193_)
  );
  al_ao21 _554_ (
    .a(_136_),
    .b(_185_),
    .c(_192_),
    .y(_194_)
  );
  al_nand2ft _555_ (
    .a(_193_),
    .b(_194_),
    .y(N726)
  );
  al_inv _556_ (
    .a(N13),
    .y(_195_)
  );
  al_and3 _557_ (
    .a(_195_),
    .b(_179_),
    .c(_185_),
    .y(_196_)
  );
  al_ao21 _558_ (
    .a(_179_),
    .b(_185_),
    .c(_195_),
    .y(_197_)
  );
  al_nand2ft _559_ (
    .a(_196_),
    .b(_197_),
    .y(N727)
  );
  al_inv _560_ (
    .a(N17),
    .y(_198_)
  );
  al_aoi21 _561_ (
    .a(_088_),
    .b(_089_),
    .c(_087_),
    .y(_199_)
  );
  al_nand3 _562_ (
    .a(_088_),
    .b(_087_),
    .c(_089_),
    .y(_200_)
  );
  al_and2ft _563_ (
    .a(_108_),
    .b(_109_),
    .y(_201_)
  );
  al_nand3ftt _564_ (
    .a(_199_),
    .b(_200_),
    .c(_201_),
    .y(_202_)
  );
  al_inv _565_ (
    .a(_202_),
    .y(_203_)
  );
  al_and3 _566_ (
    .a(_076_),
    .b(_203_),
    .c(_184_),
    .y(_204_)
  );
  al_ao21 _567_ (
    .a(_009_),
    .b(_204_),
    .c(_198_),
    .y(_205_)
  );
  al_and3 _568_ (
    .a(_198_),
    .b(_009_),
    .c(_204_),
    .y(_206_)
  );
  al_nand2ft _569_ (
    .a(_206_),
    .b(_205_),
    .y(N728)
  );
  al_inv _570_ (
    .a(N21),
    .y(_207_)
  );
  al_ao21 _571_ (
    .a(_189_),
    .b(_204_),
    .c(_207_),
    .y(_208_)
  );
  al_and3 _572_ (
    .a(_207_),
    .b(_189_),
    .c(_204_),
    .y(_209_)
  );
  al_nand2ft _573_ (
    .a(_209_),
    .b(_208_),
    .y(N729)
  );
  al_inv _574_ (
    .a(N25),
    .y(_210_)
  );
  al_and3 _575_ (
    .a(_210_),
    .b(_136_),
    .c(_204_),
    .y(_211_)
  );
  al_ao21 _576_ (
    .a(_136_),
    .b(_204_),
    .c(_210_),
    .y(_212_)
  );
  al_nand2ft _577_ (
    .a(_211_),
    .b(_212_),
    .y(N730)
  );
  al_inv _578_ (
    .a(N29),
    .y(_213_)
  );
  al_and3 _579_ (
    .a(_213_),
    .b(_179_),
    .c(_204_),
    .y(_214_)
  );
  al_ao21 _580_ (
    .a(_179_),
    .b(_204_),
    .c(_213_),
    .y(_215_)
  );
  al_nand2ft _581_ (
    .a(_214_),
    .b(_215_),
    .y(N731)
  );
  al_inv _582_ (
    .a(N33),
    .y(_216_)
  );
  al_nor2ft _583_ (
    .a(_074_),
    .b(_073_),
    .y(_217_)
  );
  al_and3ftt _584_ (
    .a(_040_),
    .b(_041_),
    .c(_217_),
    .y(_218_)
  );
  al_and3 _585_ (
    .a(_111_),
    .b(_218_),
    .c(_184_),
    .y(_219_)
  );
  al_ao21 _586_ (
    .a(_009_),
    .b(_219_),
    .c(_216_),
    .y(_220_)
  );
  al_and3 _587_ (
    .a(_216_),
    .b(_009_),
    .c(_219_),
    .y(_221_)
  );
  al_nand2ft _588_ (
    .a(_221_),
    .b(_220_),
    .y(N732)
  );
  al_inv _589_ (
    .a(N37),
    .y(_222_)
  );
  al_ao21 _590_ (
    .a(_189_),
    .b(_219_),
    .c(_222_),
    .y(_223_)
  );
  al_and3 _591_ (
    .a(_222_),
    .b(_189_),
    .c(_219_),
    .y(_224_)
  );
  al_nand2ft _592_ (
    .a(_224_),
    .b(_223_),
    .y(N733)
  );
  al_inv _593_ (
    .a(N41),
    .y(_225_)
  );
  al_and3 _594_ (
    .a(_225_),
    .b(_136_),
    .c(_219_),
    .y(_226_)
  );
  al_ao21 _595_ (
    .a(_136_),
    .b(_219_),
    .c(_225_),
    .y(_227_)
  );
  al_nand2ft _596_ (
    .a(_226_),
    .b(_227_),
    .y(N734)
  );
  al_inv _597_ (
    .a(N45),
    .y(_228_)
  );
  al_and3 _598_ (
    .a(_228_),
    .b(_179_),
    .c(_219_),
    .y(_229_)
  );
  al_ao21 _599_ (
    .a(_179_),
    .b(_219_),
    .c(_228_),
    .y(_230_)
  );
  al_nand2ft _600_ (
    .a(_229_),
    .b(_230_),
    .y(N735)
  );
  al_inv _601_ (
    .a(N49),
    .y(_231_)
  );
  al_and3 _602_ (
    .a(_203_),
    .b(_218_),
    .c(_184_),
    .y(_232_)
  );
  al_ao21 _603_ (
    .a(_009_),
    .b(_232_),
    .c(_231_),
    .y(_233_)
  );
  al_and3 _604_ (
    .a(_231_),
    .b(_009_),
    .c(_232_),
    .y(_234_)
  );
  al_nand2ft _605_ (
    .a(_234_),
    .b(_233_),
    .y(N736)
  );
  al_inv _606_ (
    .a(N53),
    .y(_235_)
  );
  al_ao21 _607_ (
    .a(_189_),
    .b(_232_),
    .c(_235_),
    .y(_236_)
  );
  al_and3 _608_ (
    .a(_235_),
    .b(_189_),
    .c(_232_),
    .y(_237_)
  );
  al_nand2ft _609_ (
    .a(_237_),
    .b(_236_),
    .y(N737)
  );
  al_inv _610_ (
    .a(N57),
    .y(_238_)
  );
  al_and3 _611_ (
    .a(_238_),
    .b(_136_),
    .c(_232_),
    .y(_239_)
  );
  al_ao21 _612_ (
    .a(_136_),
    .b(_232_),
    .c(_238_),
    .y(_240_)
  );
  al_nand2ft _613_ (
    .a(_239_),
    .b(_240_),
    .y(N738)
  );
  al_inv _614_ (
    .a(N61),
    .y(_241_)
  );
  al_ao21 _615_ (
    .a(_179_),
    .b(_232_),
    .c(_241_),
    .y(_242_)
  );
  al_and3 _616_ (
    .a(_241_),
    .b(_179_),
    .c(_232_),
    .y(_243_)
  );
  al_nand2ft _617_ (
    .a(_243_),
    .b(_242_),
    .y(N739)
  );
  al_inv _618_ (
    .a(N65),
    .y(_244_)
  );
  al_or2ft _619_ (
    .a(_041_),
    .b(_040_),
    .y(_245_)
  );
  al_nand3ftt _620_ (
    .a(_199_),
    .b(_200_),
    .c(_110_),
    .y(_246_)
  );
  al_oai21ttf _621_ (
    .a(_076_),
    .b(_218_),
    .c(_246_),
    .y(_247_)
  );
  al_nand2ft _622_ (
    .a(_111_),
    .b(_202_),
    .y(_248_)
  );
  al_and3ftt _623_ (
    .a(_040_),
    .b(_041_),
    .c(_075_),
    .y(_249_)
  );
  al_ao21ttf _624_ (
    .a(_249_),
    .b(_248_),
    .c(_247_),
    .y(_250_)
  );
  al_and3 _625_ (
    .a(_162_),
    .b(_180_),
    .c(_250_),
    .y(_251_)
  );
  al_ao21 _626_ (
    .a(_245_),
    .b(_251_),
    .c(_244_),
    .y(_252_)
  );
  al_and3 _627_ (
    .a(_244_),
    .b(_245_),
    .c(_251_),
    .y(_253_)
  );
  al_nand2ft _628_ (
    .a(_253_),
    .b(_252_),
    .y(N740)
  );
  al_inv _629_ (
    .a(N69),
    .y(_254_)
  );
  al_ao21 _630_ (
    .a(_217_),
    .b(_251_),
    .c(_254_),
    .y(_255_)
  );
  al_and3 _631_ (
    .a(_254_),
    .b(_217_),
    .c(_251_),
    .y(_256_)
  );
  al_nand2ft _632_ (
    .a(_256_),
    .b(_255_),
    .y(N741)
  );
  al_inv _633_ (
    .a(N73),
    .y(_257_)
  );
  al_nand2ft _634_ (
    .a(_199_),
    .b(_200_),
    .y(_258_)
  );
  al_and3 _635_ (
    .a(_257_),
    .b(_258_),
    .c(_251_),
    .y(_259_)
  );
  al_ao21 _636_ (
    .a(_258_),
    .b(_251_),
    .c(_257_),
    .y(_260_)
  );
  al_nand2ft _637_ (
    .a(_259_),
    .b(_260_),
    .y(N742)
  );
  al_inv _638_ (
    .a(N77),
    .y(_261_)
  );
  al_ao21 _639_ (
    .a(_201_),
    .b(_251_),
    .c(_261_),
    .y(_262_)
  );
  al_and3 _640_ (
    .a(_261_),
    .b(_201_),
    .c(_251_),
    .y(_263_)
  );
  al_nand2ft _641_ (
    .a(_263_),
    .b(_262_),
    .y(N743)
  );
  al_inv _642_ (
    .a(N81),
    .y(_264_)
  );
  al_nor3fft _643_ (
    .a(_160_),
    .b(_009_),
    .c(_136_),
    .y(_265_)
  );
  al_and3 _644_ (
    .a(_265_),
    .b(_179_),
    .c(_250_),
    .y(_266_)
  );
  al_ao21 _645_ (
    .a(_245_),
    .b(_266_),
    .c(_264_),
    .y(_267_)
  );
  al_and3 _646_ (
    .a(_264_),
    .b(_245_),
    .c(_266_),
    .y(_268_)
  );
  al_nand2ft _647_ (
    .a(_268_),
    .b(_267_),
    .y(N744)
  );
  al_inv _648_ (
    .a(N85),
    .y(_269_)
  );
  al_ao21 _649_ (
    .a(_217_),
    .b(_266_),
    .c(_269_),
    .y(_270_)
  );
  al_and3 _650_ (
    .a(_269_),
    .b(_217_),
    .c(_266_),
    .y(_271_)
  );
  al_nand2ft _651_ (
    .a(_271_),
    .b(_270_),
    .y(N745)
  );
  al_inv _652_ (
    .a(N89),
    .y(_272_)
  );
  al_ao21 _653_ (
    .a(_258_),
    .b(_266_),
    .c(_272_),
    .y(_273_)
  );
  al_and3 _654_ (
    .a(_272_),
    .b(_258_),
    .c(_266_),
    .y(_274_)
  );
  al_nand2ft _655_ (
    .a(_274_),
    .b(_273_),
    .y(N746)
  );
  al_inv _656_ (
    .a(N93),
    .y(_275_)
  );
  al_ao21 _657_ (
    .a(_201_),
    .b(_266_),
    .c(_275_),
    .y(_276_)
  );
  al_and3 _658_ (
    .a(_275_),
    .b(_201_),
    .c(_266_),
    .y(_277_)
  );
  al_nand2ft _659_ (
    .a(_277_),
    .b(_276_),
    .y(N747)
  );
  al_inv _660_ (
    .a(N97),
    .y(_278_)
  );
  al_and3fft _661_ (
    .a(_005_),
    .b(_160_),
    .c(_008_),
    .y(_279_)
  );
  al_and3 _662_ (
    .a(_279_),
    .b(_180_),
    .c(_250_),
    .y(_280_)
  );
  al_ao21 _663_ (
    .a(_245_),
    .b(_280_),
    .c(_278_),
    .y(_281_)
  );
  al_and3 _664_ (
    .a(_278_),
    .b(_245_),
    .c(_280_),
    .y(_282_)
  );
  al_nand2ft _665_ (
    .a(_282_),
    .b(_281_),
    .y(N748)
  );
  al_inv _666_ (
    .a(N101),
    .y(_283_)
  );
  al_ao21 _667_ (
    .a(_217_),
    .b(_280_),
    .c(_283_),
    .y(_284_)
  );
  al_and3 _668_ (
    .a(_283_),
    .b(_217_),
    .c(_280_),
    .y(_285_)
  );
  al_nand2ft _669_ (
    .a(_285_),
    .b(_284_),
    .y(N749)
  );
  al_inv _670_ (
    .a(N105),
    .y(_286_)
  );
  al_and3 _671_ (
    .a(_286_),
    .b(_258_),
    .c(_280_),
    .y(_287_)
  );
  al_ao21 _672_ (
    .a(_258_),
    .b(_280_),
    .c(_286_),
    .y(_288_)
  );
  al_nand2ft _673_ (
    .a(_287_),
    .b(_288_),
    .y(N750)
  );
  al_inv _674_ (
    .a(N109),
    .y(_289_)
  );
  al_ao21 _675_ (
    .a(_201_),
    .b(_280_),
    .c(_289_),
    .y(_290_)
  );
  al_and3 _676_ (
    .a(_289_),
    .b(_201_),
    .c(_280_),
    .y(_291_)
  );
  al_nand2ft _677_ (
    .a(_291_),
    .b(_290_),
    .y(N751)
  );
  al_inv _678_ (
    .a(N113),
    .y(_292_)
  );
  al_inv _679_ (
    .a(_161_),
    .y(_293_)
  );
  al_and3 _680_ (
    .a(_293_),
    .b(_179_),
    .c(_250_),
    .y(_294_)
  );
  al_ao21 _681_ (
    .a(_245_),
    .b(_294_),
    .c(_292_),
    .y(_295_)
  );
  al_and3 _682_ (
    .a(_292_),
    .b(_245_),
    .c(_294_),
    .y(_296_)
  );
  al_nand2ft _683_ (
    .a(_296_),
    .b(_295_),
    .y(N752)
  );
  al_inv _684_ (
    .a(N117),
    .y(_297_)
  );
  al_ao21 _685_ (
    .a(_217_),
    .b(_294_),
    .c(_297_),
    .y(_298_)
  );
  al_and3 _686_ (
    .a(_297_),
    .b(_217_),
    .c(_294_),
    .y(_299_)
  );
  al_nand2ft _687_ (
    .a(_299_),
    .b(_298_),
    .y(N753)
  );
  al_inv _688_ (
    .a(N121),
    .y(_300_)
  );
  al_ao21 _689_ (
    .a(_258_),
    .b(_294_),
    .c(_300_),
    .y(_301_)
  );
  al_and3 _690_ (
    .a(_300_),
    .b(_258_),
    .c(_294_),
    .y(_302_)
  );
  al_nand2ft _691_ (
    .a(_302_),
    .b(_301_),
    .y(N754)
  );
  al_inv _692_ (
    .a(N125),
    .y(_303_)
  );
  al_ao21 _693_ (
    .a(_201_),
    .b(_294_),
    .c(_303_),
    .y(_304_)
  );
  al_and3 _694_ (
    .a(_303_),
    .b(_201_),
    .c(_294_),
    .y(_305_)
  );
  al_nand2ft _695_ (
    .a(_305_),
    .b(_304_),
    .y(N755)
  );
endmodule
