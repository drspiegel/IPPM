
module c3540(N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97, N107, N116, N124, N125, N128, N132, N137, N143, N150, N159, N169, N179, N190, N200, N213, N222, N223, N226, N232, N238, N244, N250, N257, N264, N270, N274, N283, N294, N303, N311, N317, N322, N326, N329, N330, N343, N349, N350, N1713, N1947, N3195, N3833, N3987, N4028, N4145, N4589, N4667, N4815, N4944, N5002, N5045, N5047, N5078, N5102, N5120, N5121, N5192, N5231, N5360, N5361);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  input N1;
  input N107;
  input N116;
  input N124;
  input N125;
  wire N1279;
  input N128;
  input N13;
  input N132;
  wire N1334;
  wire N1345;
  wire N1346;
  wire N1347;
  wire N1348;
  wire N1349;
  wire N1350;
  wire N1351;
  wire N1352;
  wire N1369;
  input N137;
  input N143;
  wire N1493;
  wire N1496;
  wire N1499;
  input N150;
  wire N1502;
  input N159;
  input N169;
  output N1713;
  wire N1726;
  wire N1735;
  wire N1736;
  wire N1737;
  input N179;
  wire N1849;
  wire N1851;
  wire N1853;
  wire N1855;
  wire N1857;
  wire N1859;
  wire N1861;
  wire N1863;
  input N190;
  wire N1939;
  wire N1941;
  wire N1942;
  wire N1943;
  wire N1944;
  wire N1945;
  wire N1946;
  output N1947;
  input N20;
  input N200;
  input N213;
  input N222;
  input N223;
  input N226;
  input N232;
  input N238;
  input N244;
  input N250;
  input N257;
  input N264;
  input N270;
  input N274;
  input N283;
  input N294;
  input N303;
  input N311;
  input N317;
  output N3195;
  input N322;
  input N326;
  input N329;
  input N33;
  input N330;
  input N343;
  input N349;
  input N350;
  output N3833;
  output N3987;
  output N4028;
  input N41;
  output N4145;
  input N45;
  output N4589;
  output N4667;
  output N4815;
  output N4944;
  input N50;
  output N5002;
  output N5045;
  output N5047;
  output N5078;
  output N5102;
  output N5120;
  output N5121;
  output N5192;
  output N5231;
  output N5360;
  output N5361;
  input N58;
  wire N655;
  wire N670;
  input N68;
  wire N683;
  wire N690;
  wire N699;
  wire N706;
  wire N715;
  wire N727;
  wire N740;
  wire N753;
  input N77;
  wire N772;
  wire N782;
  wire N798;
  wire N821;
  wire N836;
  wire N845;
  wire N851;
  wire N858;
  wire N864;
  input N87;
  wire N874;
  wire N877;
  wire N880;
  wire N886;
  wire N917;
  wire N923;
  wire N926;
  wire N929;
  wire N932;
  wire N935;
  wire N938;
  wire N941;
  wire N944;
  wire N947;
  wire N950;
  wire N953;
  wire N956;
  wire N959;
  wire N962;
  wire N965;
  input N97;
  al_oai21 _0646_ (
    .a(N97),
    .b(N107),
    .c(N87),
    .y(N1947)
  );
  al_and2 _0647_ (
    .a(N20),
    .b(N1),
    .y(_0621_)
  );
  al_oa21 _0648_ (
    .a(N257),
    .b(N264),
    .c(N250),
    .y(_0622_)
  );
  al_oa21 _0649_ (
    .a(N58),
    .b(N68),
    .c(N50),
    .y(_0623_)
  );
  al_mux2l _0650_ (
    .a(_0623_),
    .b(_0622_),
    .s(N13),
    .y(_0624_)
  );
  al_nand2 _0651_ (
    .a(N238),
    .b(N68),
    .y(_0625_)
  );
  al_aoi21ttf _0652_ (
    .a(N264),
    .b(N107),
    .c(_0625_),
    .y(_0626_)
  );
  al_nand2 _0653_ (
    .a(N87),
    .b(N250),
    .y(_0627_)
  );
  al_aoi21ttf _0654_ (
    .a(N226),
    .b(N50),
    .c(_0627_),
    .y(_0628_)
  );
  al_nand2 _0655_ (
    .a(N77),
    .b(N244),
    .y(_0629_)
  );
  al_nand2 _0656_ (
    .a(N97),
    .b(N257),
    .y(_0630_)
  );
  al_nand2 _0657_ (
    .a(N232),
    .b(N58),
    .y(_0631_)
  );
  al_nand2 _0658_ (
    .a(N116),
    .b(N270),
    .y(_0632_)
  );
  al_and3 _0659_ (
    .a(_0630_),
    .b(_0631_),
    .c(_0632_),
    .y(_0633_)
  );
  al_and3 _0660_ (
    .a(_0629_),
    .b(_0628_),
    .c(_0633_),
    .y(_0634_)
  );
  al_nand3ftt _0661_ (
    .a(_0621_),
    .b(_0626_),
    .c(_0634_),
    .y(_0635_)
  );
  al_ao21ftf _0662_ (
    .a(_0624_),
    .b(_0621_),
    .c(_0635_),
    .y(N3195)
  );
  al_and2ft _0663_ (
    .a(N264),
    .b(N270),
    .y(_0636_)
  );
  al_nand2ft _0664_ (
    .a(N270),
    .b(N264),
    .y(_0637_)
  );
  al_nand2 _0665_ (
    .a(N250),
    .b(N257),
    .y(_0638_)
  );
  al_nor2 _0666_ (
    .a(N250),
    .b(N257),
    .y(_0639_)
  );
  al_nand2ft _0667_ (
    .a(_0639_),
    .b(_0638_),
    .y(_0640_)
  );
  al_and3ftt _0668_ (
    .a(_0636_),
    .b(_0637_),
    .c(_0640_),
    .y(_0641_)
  );
  al_aoi21ftt _0669_ (
    .a(_0636_),
    .b(_0637_),
    .c(_0640_),
    .y(_0642_)
  );
  al_or2 _0670_ (
    .a(_0641_),
    .b(_0642_),
    .y(_0643_)
  );
  al_and2ft _0671_ (
    .a(N238),
    .b(N244),
    .y(_0644_)
  );
  al_nand2ft _0672_ (
    .a(N244),
    .b(N238),
    .y(_0645_)
  );
  al_and2ft _0673_ (
    .a(N232),
    .b(N226),
    .y(_0000_)
  );
  al_nand2ft _0674_ (
    .a(N226),
    .b(N232),
    .y(_0001_)
  );
  al_nand2ft _0675_ (
    .a(_0000_),
    .b(_0001_),
    .y(_0002_)
  );
  al_and3ftt _0676_ (
    .a(_0644_),
    .b(_0645_),
    .c(_0002_),
    .y(_0003_)
  );
  al_ao21ftt _0677_ (
    .a(_0644_),
    .b(_0645_),
    .c(_0002_),
    .y(_0004_)
  );
  al_ao21ftt _0678_ (
    .a(_0003_),
    .b(_0004_),
    .c(_0643_),
    .y(_0005_)
  );
  al_and3ftt _0679_ (
    .a(_0003_),
    .b(_0004_),
    .c(_0643_),
    .y(_0006_)
  );
  al_nand2ft _0680_ (
    .a(_0006_),
    .b(_0005_),
    .y(N3833)
  );
  al_nor2 _0681_ (
    .a(N58),
    .b(N50),
    .y(_0007_)
  );
  al_nand2 _0682_ (
    .a(N58),
    .b(N50),
    .y(_0008_)
  );
  al_nand2ft _0683_ (
    .a(_0007_),
    .b(_0008_),
    .y(_0009_)
  );
  al_nand2 _0684_ (
    .a(N77),
    .b(N68),
    .y(_0010_)
  );
  al_or2 _0685_ (
    .a(N77),
    .b(N68),
    .y(_0011_)
  );
  al_ao21 _0686_ (
    .a(_0010_),
    .b(_0011_),
    .c(_0009_),
    .y(_0012_)
  );
  al_and3 _0687_ (
    .a(_0010_),
    .b(_0011_),
    .c(_0009_),
    .y(_0013_)
  );
  al_nor2 _0688_ (
    .a(N97),
    .b(N107),
    .y(_0014_)
  );
  al_nand2 _0689_ (
    .a(N97),
    .b(N107),
    .y(_0015_)
  );
  al_nand2ft _0690_ (
    .a(_0014_),
    .b(_0015_),
    .y(_0016_)
  );
  al_and2ft _0691_ (
    .a(N116),
    .b(N87),
    .y(_0017_)
  );
  al_nand2ft _0692_ (
    .a(N87),
    .b(N116),
    .y(_0018_)
  );
  al_aoi21ftt _0693_ (
    .a(_0017_),
    .b(_0018_),
    .c(_0016_),
    .y(_0019_)
  );
  al_nand3ftt _0694_ (
    .a(_0017_),
    .b(_0018_),
    .c(_0016_),
    .y(_0020_)
  );
  al_or2ft _0695_ (
    .a(_0020_),
    .b(_0019_),
    .y(_0021_)
  );
  al_ao21ftt _0696_ (
    .a(_0013_),
    .b(_0012_),
    .c(_0021_),
    .y(_0022_)
  );
  al_and3ftt _0697_ (
    .a(_0013_),
    .b(_0012_),
    .c(_0021_),
    .y(_0023_)
  );
  al_nand2ft _0698_ (
    .a(_0023_),
    .b(_0022_),
    .y(N3987)
  );
  al_nand3ftt _0699_ (
    .a(N1),
    .b(N13),
    .c(N20),
    .y(_0024_)
  );
  al_nand2ft _0700_ (
    .a(N1),
    .b(N20),
    .y(_0025_)
  );
  al_and2 _0701_ (
    .a(N13),
    .b(N1),
    .y(_0026_)
  );
  al_nand3 _0702_ (
    .a(N20),
    .b(N1),
    .c(N33),
    .y(_0027_)
  );
  al_or3fft _0703_ (
    .a(_0025_),
    .b(_0027_),
    .c(_0026_),
    .y(_0028_)
  );
  al_mux2h _0704_ (
    .a(_0024_),
    .b(_0028_),
    .s(N50),
    .y(_0029_)
  );
  al_aoi21ttf _0705_ (
    .a(N13),
    .b(N1),
    .c(_0027_),
    .y(_0030_)
  );
  al_nand3fft _0706_ (
    .a(N20),
    .b(N33),
    .c(N150),
    .y(_0031_)
  );
  al_or3 _0707_ (
    .a(N58),
    .b(N50),
    .c(N68),
    .y(_0032_)
  );
  al_and3ftt _0708_ (
    .a(N20),
    .b(N58),
    .c(N33),
    .y(_0033_)
  );
  al_aoi21 _0709_ (
    .a(N20),
    .b(_0032_),
    .c(_0033_),
    .y(_0034_)
  );
  al_ao21 _0710_ (
    .a(_0031_),
    .b(_0034_),
    .c(_0030_),
    .y(_0035_)
  );
  al_and2 _0711_ (
    .a(_0035_),
    .b(_0029_),
    .y(_0036_)
  );
  al_nand2 _0712_ (
    .a(N41),
    .b(N33),
    .y(_0037_)
  );
  al_nand3 _0713_ (
    .a(N13),
    .b(N1),
    .c(_0037_),
    .y(_0038_)
  );
  al_nand3ftt _0714_ (
    .a(N33),
    .b(N349),
    .c(N223),
    .y(_0039_)
  );
  al_nand3fft _0715_ (
    .a(N33),
    .b(N349),
    .c(N222),
    .y(_0040_)
  );
  al_aoi21ttf _0716_ (
    .a(N77),
    .b(N33),
    .c(_0040_),
    .y(_0041_)
  );
  al_ao21 _0717_ (
    .a(_0039_),
    .b(_0041_),
    .c(_0038_),
    .y(_0042_)
  );
  al_oai21ttf _0718_ (
    .a(N41),
    .b(N45),
    .c(N1),
    .y(_0043_)
  );
  al_and3ftt _0719_ (
    .a(_0043_),
    .b(N274),
    .c(_0038_),
    .y(_0044_)
  );
  al_nand3 _0720_ (
    .a(N226),
    .b(_0043_),
    .c(_0038_),
    .y(_0045_)
  );
  al_nand3ftt _0721_ (
    .a(_0044_),
    .b(_0042_),
    .c(_0045_),
    .y(_0046_)
  );
  al_mux2l _0722_ (
    .a(N200),
    .b(N190),
    .s(_0046_),
    .y(_0047_)
  );
  al_inv _0723_ (
    .a(N179),
    .y(_0048_)
  );
  al_inv _0724_ (
    .a(N169),
    .y(_0049_)
  );
  al_mux2l _0725_ (
    .a(_0049_),
    .b(_0048_),
    .s(_0046_),
    .y(_0050_)
  );
  al_mux2l _0726_ (
    .a(_0047_),
    .b(_0050_),
    .s(_0036_),
    .y(_0051_)
  );
  al_nand3ftt _0727_ (
    .a(N33),
    .b(N226),
    .c(N349),
    .y(_0052_)
  );
  al_nand3fft _0728_ (
    .a(N33),
    .b(N349),
    .c(N223),
    .y(_0053_)
  );
  al_aoi21ttf _0729_ (
    .a(N87),
    .b(N33),
    .c(_0053_),
    .y(_0054_)
  );
  al_ao21 _0730_ (
    .a(_0052_),
    .b(_0054_),
    .c(_0038_),
    .y(_0055_)
  );
  al_aoi21ttf _0731_ (
    .a(_0037_),
    .b(_0026_),
    .c(_0043_),
    .y(_0056_)
  );
  al_aoi21 _0732_ (
    .a(N232),
    .b(_0056_),
    .c(_0044_),
    .y(_0057_)
  );
  al_nand3 _0733_ (
    .a(_0048_),
    .b(_0055_),
    .c(_0057_),
    .y(_0058_)
  );
  al_ao21 _0734_ (
    .a(_0055_),
    .b(_0057_),
    .c(N169),
    .y(_0059_)
  );
  al_nand3fft _0735_ (
    .a(N20),
    .b(N33),
    .c(N159),
    .y(_0060_)
  );
  al_inv _0736_ (
    .a(N20),
    .y(_0061_)
  );
  al_or2 _0737_ (
    .a(N58),
    .b(N68),
    .y(_0062_)
  );
  al_nand2 _0738_ (
    .a(N58),
    .b(N68),
    .y(_0063_)
  );
  al_ao21 _0739_ (
    .a(_0062_),
    .b(_0063_),
    .c(_0061_),
    .y(_0064_)
  );
  al_nand3ftt _0740_ (
    .a(N20),
    .b(N68),
    .c(N33),
    .y(_0065_)
  );
  al_nand3 _0741_ (
    .a(_0060_),
    .b(_0065_),
    .c(_0064_),
    .y(_0066_)
  );
  al_mux2h _0742_ (
    .a(_0024_),
    .b(_0028_),
    .s(N58),
    .y(_0067_)
  );
  al_ao21ftf _0743_ (
    .a(_0030_),
    .b(_0066_),
    .c(_0067_),
    .y(_0068_)
  );
  al_nand3 _0744_ (
    .a(_0068_),
    .b(_0058_),
    .c(_0059_),
    .y(_0069_)
  );
  al_nand3 _0745_ (
    .a(N190),
    .b(_0055_),
    .c(_0057_),
    .y(_0070_)
  );
  al_inv _0746_ (
    .a(N200),
    .y(_0071_)
  );
  al_ao21 _0747_ (
    .a(_0055_),
    .b(_0057_),
    .c(_0071_),
    .y(_0072_)
  );
  al_nand3ftt _0748_ (
    .a(_0068_),
    .b(_0070_),
    .c(_0072_),
    .y(_0073_)
  );
  al_and3 _0749_ (
    .a(_0069_),
    .b(_0073_),
    .c(_0051_),
    .y(_0074_)
  );
  al_nand3ftt _0750_ (
    .a(N20),
    .b(N13),
    .c(N1),
    .y(_0075_)
  );
  al_mux2l _0751_ (
    .a(N87),
    .b(N58),
    .s(N33),
    .y(_0076_)
  );
  al_and3ftt _0752_ (
    .a(N1),
    .b(N13),
    .c(N20),
    .y(_0077_)
  );
  al_nand3 _0753_ (
    .a(N77),
    .b(_0075_),
    .c(_0025_),
    .y(_0078_)
  );
  al_aoi21ftf _0754_ (
    .a(N77),
    .b(_0077_),
    .c(_0078_),
    .y(_0079_)
  );
  al_ao21ftf _0755_ (
    .a(_0075_),
    .b(_0076_),
    .c(_0079_),
    .y(_0080_)
  );
  al_nand3ftt _0756_ (
    .a(N33),
    .b(N238),
    .c(N349),
    .y(_0081_)
  );
  al_and3fft _0757_ (
    .a(N33),
    .b(N349),
    .c(N232),
    .y(_0082_)
  );
  al_aoi21 _0758_ (
    .a(N107),
    .b(N33),
    .c(_0082_),
    .y(_0083_)
  );
  al_ao21 _0759_ (
    .a(_0081_),
    .b(_0083_),
    .c(_0038_),
    .y(_0084_)
  );
  al_aoi21 _0760_ (
    .a(N244),
    .b(_0056_),
    .c(_0044_),
    .y(_0085_)
  );
  al_ao21 _0761_ (
    .a(_0084_),
    .b(_0085_),
    .c(N169),
    .y(_0086_)
  );
  al_nand3 _0762_ (
    .a(_0048_),
    .b(_0084_),
    .c(_0085_),
    .y(_0087_)
  );
  al_nand3 _0763_ (
    .a(_0080_),
    .b(_0087_),
    .c(_0086_),
    .y(_0088_)
  );
  al_ao21 _0764_ (
    .a(_0084_),
    .b(_0085_),
    .c(_0071_),
    .y(_0089_)
  );
  al_nand3 _0765_ (
    .a(N190),
    .b(_0084_),
    .c(_0085_),
    .y(_0090_)
  );
  al_nand3ftt _0766_ (
    .a(_0080_),
    .b(_0090_),
    .c(_0089_),
    .y(_0091_)
  );
  al_and2 _0767_ (
    .a(_0088_),
    .b(_0091_),
    .y(_0092_)
  );
  al_and2ft _0768_ (
    .a(N20),
    .b(N13),
    .y(_0093_)
  );
  al_mux2l _0769_ (
    .a(N77),
    .b(N50),
    .s(N33),
    .y(_0094_)
  );
  al_nand3 _0770_ (
    .a(N1),
    .b(_0094_),
    .c(_0093_),
    .y(_0095_)
  );
  al_ao21ttf _0771_ (
    .a(N13),
    .b(N20),
    .c(_0027_),
    .y(_0096_)
  );
  al_aoi21ftf _0772_ (
    .a(N68),
    .b(_0096_),
    .c(_0095_),
    .y(_0097_)
  );
  al_ao21ftf _0773_ (
    .a(_0028_),
    .b(N68),
    .c(_0097_),
    .y(_0098_)
  );
  al_nand3ftt _0774_ (
    .a(N33),
    .b(N232),
    .c(N349),
    .y(_0099_)
  );
  al_and3fft _0775_ (
    .a(N33),
    .b(N349),
    .c(N226),
    .y(_0100_)
  );
  al_aoi21 _0776_ (
    .a(N97),
    .b(N33),
    .c(_0100_),
    .y(_0101_)
  );
  al_ao21 _0777_ (
    .a(_0099_),
    .b(_0101_),
    .c(_0038_),
    .y(_0102_)
  );
  al_aoi21 _0778_ (
    .a(N238),
    .b(_0056_),
    .c(_0044_),
    .y(_0103_)
  );
  al_ao21 _0779_ (
    .a(_0102_),
    .b(_0103_),
    .c(N169),
    .y(_0104_)
  );
  al_nand3 _0780_ (
    .a(_0048_),
    .b(_0102_),
    .c(_0103_),
    .y(_0105_)
  );
  al_and3 _0781_ (
    .a(_0098_),
    .b(_0105_),
    .c(_0104_),
    .y(_0106_)
  );
  al_nand3 _0782_ (
    .a(N190),
    .b(_0102_),
    .c(_0103_),
    .y(_0107_)
  );
  al_ao21 _0783_ (
    .a(_0102_),
    .b(_0103_),
    .c(_0071_),
    .y(_0108_)
  );
  al_nand3ftt _0784_ (
    .a(_0098_),
    .b(_0107_),
    .c(_0108_),
    .y(_0109_)
  );
  al_nand2ft _0785_ (
    .a(_0106_),
    .b(_0109_),
    .y(_0110_)
  );
  al_and3ftt _0786_ (
    .a(_0110_),
    .b(_0092_),
    .c(_0074_),
    .y(_0111_)
  );
  al_nand2ft _0787_ (
    .a(N87),
    .b(_0024_),
    .y(_0112_)
  );
  al_aoi21ftf _0788_ (
    .a(N1),
    .b(N33),
    .c(_0024_),
    .y(_0113_)
  );
  al_ao21ttf _0789_ (
    .a(_0113_),
    .b(_0030_),
    .c(N87),
    .y(_0114_)
  );
  al_or3ftt _0790_ (
    .a(N68),
    .b(N20),
    .c(N33),
    .y(_0115_)
  );
  al_or3 _0791_ (
    .a(N87),
    .b(N97),
    .c(N107),
    .y(_0116_)
  );
  al_aoi21 _0792_ (
    .a(N97),
    .b(N33),
    .c(N20),
    .y(_0117_)
  );
  al_oai21ftf _0793_ (
    .a(N20),
    .b(_0116_),
    .c(_0117_),
    .y(_0118_)
  );
  al_ao21 _0794_ (
    .a(_0115_),
    .b(_0118_),
    .c(_0030_),
    .y(_0119_)
  );
  al_aoi21ttf _0795_ (
    .a(_0112_),
    .b(_0114_),
    .c(_0119_),
    .y(_0120_)
  );
  al_nand2ft _0796_ (
    .a(N1),
    .b(N45),
    .y(_0121_)
  );
  al_mux2l _0797_ (
    .a(N250),
    .b(N274),
    .s(_0121_),
    .y(_0122_)
  );
  al_and3ftt _0798_ (
    .a(N33),
    .b(N244),
    .c(N349),
    .y(_0123_)
  );
  al_and3fft _0799_ (
    .a(N33),
    .b(N349),
    .c(N238),
    .y(_0124_)
  );
  al_nand2 _0800_ (
    .a(N116),
    .b(N33),
    .y(_0125_)
  );
  al_nand3fft _0801_ (
    .a(_0123_),
    .b(_0124_),
    .c(_0125_),
    .y(_0126_)
  );
  al_mux2l _0802_ (
    .a(_0122_),
    .b(_0126_),
    .s(_0038_),
    .y(_0127_)
  );
  al_mux2l _0803_ (
    .a(N200),
    .b(N190),
    .s(_0127_),
    .y(_0128_)
  );
  al_mux2l _0804_ (
    .a(_0049_),
    .b(_0048_),
    .s(_0127_),
    .y(_0129_)
  );
  al_mux2l _0805_ (
    .a(_0128_),
    .b(_0129_),
    .s(_0120_),
    .y(_0130_)
  );
  al_or3fft _0806_ (
    .a(N20),
    .b(_0015_),
    .c(_0014_),
    .y(_0131_)
  );
  al_mux2l _0807_ (
    .a(N107),
    .b(N77),
    .s(N33),
    .y(_0132_)
  );
  al_or2 _0808_ (
    .a(N20),
    .b(_0132_),
    .y(_0133_)
  );
  al_nand3ftt _0809_ (
    .a(_0030_),
    .b(_0131_),
    .c(_0133_),
    .y(_0134_)
  );
  al_nand2ft _0810_ (
    .a(N97),
    .b(_0077_),
    .y(_0135_)
  );
  al_nand3 _0811_ (
    .a(N97),
    .b(_0113_),
    .c(_0030_),
    .y(_0136_)
  );
  al_nand3 _0812_ (
    .a(_0135_),
    .b(_0136_),
    .c(_0134_),
    .y(_0137_)
  );
  al_or3ftt _0813_ (
    .a(N45),
    .b(N41),
    .c(N1),
    .y(_0138_)
  );
  al_nand3ftt _0814_ (
    .a(_0138_),
    .b(N274),
    .c(_0038_),
    .y(_0139_)
  );
  al_nand3ftt _0815_ (
    .a(N33),
    .b(N250),
    .c(N349),
    .y(_0140_)
  );
  al_nand2 _0816_ (
    .a(N33),
    .b(N283),
    .y(_0141_)
  );
  al_and3fft _0817_ (
    .a(N33),
    .b(N349),
    .c(N244),
    .y(_0142_)
  );
  al_and3ftt _0818_ (
    .a(_0142_),
    .b(_0140_),
    .c(_0141_),
    .y(_0143_)
  );
  al_nand2 _0819_ (
    .a(N257),
    .b(_0138_),
    .y(_0144_)
  );
  al_mux2l _0820_ (
    .a(_0144_),
    .b(_0143_),
    .s(_0038_),
    .y(_0145_)
  );
  al_aoi21 _0821_ (
    .a(_0139_),
    .b(_0145_),
    .c(N169),
    .y(_0146_)
  );
  al_and3ftt _0822_ (
    .a(_0138_),
    .b(N274),
    .c(_0038_),
    .y(_0147_)
  );
  al_nand3fft _0823_ (
    .a(N179),
    .b(_0147_),
    .c(_0145_),
    .y(_0148_)
  );
  al_or3fft _0824_ (
    .a(_0137_),
    .b(_0148_),
    .c(_0146_),
    .y(_0149_)
  );
  al_inv _0825_ (
    .a(N190),
    .y(_0150_)
  );
  al_nand3fft _0826_ (
    .a(_0150_),
    .b(_0147_),
    .c(_0145_),
    .y(_0151_)
  );
  al_ao21 _0827_ (
    .a(_0139_),
    .b(_0145_),
    .c(_0071_),
    .y(_0152_)
  );
  al_and3ftt _0828_ (
    .a(_0137_),
    .b(_0151_),
    .c(_0152_),
    .y(_0153_)
  );
  al_and3ftt _0829_ (
    .a(_0153_),
    .b(_0149_),
    .c(_0130_),
    .y(_0154_)
  );
  al_nand3ftt _0830_ (
    .a(N33),
    .b(N257),
    .c(N349),
    .y(_0155_)
  );
  al_and3fft _0831_ (
    .a(N33),
    .b(N349),
    .c(N250),
    .y(_0156_)
  );
  al_aoi21 _0832_ (
    .a(N33),
    .b(N294),
    .c(_0156_),
    .y(_0157_)
  );
  al_ao21 _0833_ (
    .a(_0155_),
    .b(_0157_),
    .c(_0038_),
    .y(_0158_)
  );
  al_ao21ttf _0834_ (
    .a(_0037_),
    .b(_0026_),
    .c(N274),
    .y(_0159_)
  );
  al_inv _0835_ (
    .a(N264),
    .y(_0160_)
  );
  al_ao21 _0836_ (
    .a(_0037_),
    .b(_0026_),
    .c(_0160_),
    .y(_0161_)
  );
  al_mux2l _0837_ (
    .a(_0161_),
    .b(_0159_),
    .s(_0138_),
    .y(_0162_)
  );
  al_nand3 _0838_ (
    .a(_0048_),
    .b(_0158_),
    .c(_0162_),
    .y(_0163_)
  );
  al_ao21 _0839_ (
    .a(_0158_),
    .b(_0162_),
    .c(N169),
    .y(_0164_)
  );
  al_mux2l _0840_ (
    .a(N116),
    .b(N87),
    .s(N33),
    .y(_0165_)
  );
  al_nand3 _0841_ (
    .a(N1),
    .b(_0165_),
    .c(_0093_),
    .y(_0166_)
  );
  al_inv _0842_ (
    .a(N107),
    .y(_0167_)
  );
  al_nand2 _0843_ (
    .a(_0167_),
    .b(_0096_),
    .y(_0168_)
  );
  al_nand3 _0844_ (
    .a(N107),
    .b(_0113_),
    .c(_0030_),
    .y(_0169_)
  );
  al_nand3 _0845_ (
    .a(_0166_),
    .b(_0168_),
    .c(_0169_),
    .y(_0170_)
  );
  al_nand3 _0846_ (
    .a(_0170_),
    .b(_0163_),
    .c(_0164_),
    .y(_0171_)
  );
  al_nand3 _0847_ (
    .a(N116),
    .b(_0113_),
    .c(_0030_),
    .y(_0172_)
  );
  al_nand2 _0848_ (
    .a(N116),
    .b(N20),
    .y(_0173_)
  );
  al_oai21ftf _0849_ (
    .a(_0027_),
    .b(_0026_),
    .c(_0173_),
    .y(_0174_)
  );
  al_mux2l _0850_ (
    .a(N283),
    .b(N97),
    .s(N33),
    .y(_0175_)
  );
  al_nand2ft _0851_ (
    .a(N116),
    .b(_0077_),
    .y(_0176_)
  );
  al_aoi21ftf _0852_ (
    .a(_0075_),
    .b(_0175_),
    .c(_0176_),
    .y(_0177_)
  );
  al_nand3 _0853_ (
    .a(_0174_),
    .b(_0177_),
    .c(_0172_),
    .y(_0178_)
  );
  al_nand3ftt _0854_ (
    .a(N33),
    .b(N264),
    .c(N349),
    .y(_0179_)
  );
  al_and3fft _0855_ (
    .a(N33),
    .b(N349),
    .c(N257),
    .y(_0180_)
  );
  al_aoi21 _0856_ (
    .a(N33),
    .b(N303),
    .c(_0180_),
    .y(_0181_)
  );
  al_ao21 _0857_ (
    .a(_0179_),
    .b(_0181_),
    .c(_0038_),
    .y(_0182_)
  );
  al_ao21ttf _0858_ (
    .a(_0037_),
    .b(_0026_),
    .c(N270),
    .y(_0183_)
  );
  al_mux2l _0859_ (
    .a(_0183_),
    .b(_0159_),
    .s(_0138_),
    .y(_0184_)
  );
  al_ao21 _0860_ (
    .a(_0182_),
    .b(_0184_),
    .c(N169),
    .y(_0185_)
  );
  al_nand3 _0861_ (
    .a(_0048_),
    .b(_0182_),
    .c(_0184_),
    .y(_0186_)
  );
  al_nand3 _0862_ (
    .a(_0178_),
    .b(_0186_),
    .c(_0185_),
    .y(_0187_)
  );
  al_ao21 _0863_ (
    .a(_0158_),
    .b(_0162_),
    .c(_0071_),
    .y(_0188_)
  );
  al_nand3 _0864_ (
    .a(N190),
    .b(_0158_),
    .c(_0162_),
    .y(_0189_)
  );
  al_nand3ftt _0865_ (
    .a(_0170_),
    .b(_0189_),
    .c(_0188_),
    .y(_0190_)
  );
  al_oa21ftt _0866_ (
    .a(_0190_),
    .b(_0187_),
    .c(_0171_),
    .y(_0191_)
  );
  al_ao21ttf _0867_ (
    .a(_0112_),
    .b(_0114_),
    .c(_0119_),
    .y(_0192_)
  );
  al_or2 _0868_ (
    .a(_0192_),
    .b(_0128_),
    .y(_0193_)
  );
  al_nor2 _0869_ (
    .a(_0120_),
    .b(_0129_),
    .y(_0194_)
  );
  al_nor3fft _0870_ (
    .a(_0137_),
    .b(_0148_),
    .c(_0146_),
    .y(_0195_)
  );
  al_ao21 _0871_ (
    .a(_0193_),
    .b(_0195_),
    .c(_0194_),
    .y(_0196_)
  );
  al_oai21ftf _0872_ (
    .a(_0154_),
    .b(_0191_),
    .c(_0196_),
    .y(_0197_)
  );
  al_oai21ftf _0873_ (
    .a(_0109_),
    .b(_0088_),
    .c(_0106_),
    .y(_0198_)
  );
  al_or3fft _0874_ (
    .a(_0029_),
    .b(_0035_),
    .c(_0047_),
    .y(_0199_)
  );
  al_or2 _0875_ (
    .a(_0036_),
    .b(_0050_),
    .y(_0200_)
  );
  al_ao21ftf _0876_ (
    .a(_0069_),
    .b(_0199_),
    .c(_0200_),
    .y(_0201_)
  );
  al_aoi21 _0877_ (
    .a(_0198_),
    .b(_0074_),
    .c(_0201_),
    .y(_0202_)
  );
  al_ao21ttf _0878_ (
    .a(_0197_),
    .b(_0111_),
    .c(_0202_),
    .y(N4145)
  );
  al_nand3ftt _0879_ (
    .a(N1),
    .b(N213),
    .c(_0093_),
    .y(_0203_)
  );
  al_and2ft _0880_ (
    .a(_0203_),
    .b(_0068_),
    .y(_0204_)
  );
  al_and3ftt _0881_ (
    .a(_0204_),
    .b(_0069_),
    .c(_0073_),
    .y(_0205_)
  );
  al_ao21ttf _0882_ (
    .a(_0069_),
    .b(_0073_),
    .c(_0204_),
    .y(_0206_)
  );
  al_nand2ft _0883_ (
    .a(_0205_),
    .b(_0206_),
    .y(_0207_)
  );
  al_nand3 _0884_ (
    .a(_0098_),
    .b(_0105_),
    .c(_0104_),
    .y(_0208_)
  );
  al_inv _0885_ (
    .a(N343),
    .y(_0209_)
  );
  al_nor2 _0886_ (
    .a(_0209_),
    .b(_0203_),
    .y(_0210_)
  );
  al_and2 _0887_ (
    .a(_0210_),
    .b(_0098_),
    .y(_0211_)
  );
  al_ao21 _0888_ (
    .a(_0208_),
    .b(_0109_),
    .c(_0211_),
    .y(_0212_)
  );
  al_and3 _0889_ (
    .a(_0211_),
    .b(_0208_),
    .c(_0109_),
    .y(_0213_)
  );
  al_nand2 _0890_ (
    .a(_0210_),
    .b(_0080_),
    .y(_0214_)
  );
  al_and3 _0891_ (
    .a(_0214_),
    .b(_0088_),
    .c(_0091_),
    .y(_0215_)
  );
  al_ao21 _0892_ (
    .a(_0088_),
    .b(_0091_),
    .c(_0214_),
    .y(_0216_)
  );
  al_nand2ft _0893_ (
    .a(_0215_),
    .b(_0216_),
    .y(_0217_)
  );
  al_and3ftt _0894_ (
    .a(_0213_),
    .b(_0212_),
    .c(_0217_),
    .y(_0218_)
  );
  al_inv _0895_ (
    .a(_0210_),
    .y(_0219_)
  );
  al_and2 _0896_ (
    .a(_0219_),
    .b(_0197_),
    .y(_0220_)
  );
  al_and2 _0897_ (
    .a(_0219_),
    .b(_0198_),
    .y(_0221_)
  );
  al_aoi21 _0898_ (
    .a(_0220_),
    .b(_0218_),
    .c(_0221_),
    .y(_0222_)
  );
  al_and3 _0899_ (
    .a(N264),
    .b(_0138_),
    .c(_0038_),
    .y(_0223_)
  );
  al_nand3ftt _0900_ (
    .a(_0223_),
    .b(_0139_),
    .c(_0158_),
    .y(_0224_)
  );
  al_mux2l _0901_ (
    .a(_0071_),
    .b(_0150_),
    .s(_0224_),
    .y(_0225_)
  );
  al_ao21ftf _0902_ (
    .a(_0170_),
    .b(_0225_),
    .c(_0171_),
    .y(_0226_)
  );
  al_and3 _0903_ (
    .a(N190),
    .b(_0182_),
    .c(_0184_),
    .y(_0227_)
  );
  al_and3 _0904_ (
    .a(N270),
    .b(_0138_),
    .c(_0038_),
    .y(_0228_)
  );
  al_nand3ftt _0905_ (
    .a(_0228_),
    .b(_0139_),
    .c(_0182_),
    .y(_0229_)
  );
  al_aoi21 _0906_ (
    .a(N200),
    .b(_0229_),
    .c(_0178_),
    .y(_0230_)
  );
  al_aoi21ftf _0907_ (
    .a(_0227_),
    .b(_0230_),
    .c(_0187_),
    .y(_0231_)
  );
  al_nand3ftt _0908_ (
    .a(_0226_),
    .b(_0231_),
    .c(_0154_),
    .y(_0232_)
  );
  al_or2 _0909_ (
    .a(_0048_),
    .b(_0127_),
    .y(_0233_)
  );
  al_and3fft _0910_ (
    .a(_0147_),
    .b(_0224_),
    .c(_0145_),
    .y(_0234_)
  );
  al_nand3fft _0911_ (
    .a(_0233_),
    .b(_0229_),
    .c(_0234_),
    .y(_0235_)
  );
  al_aoi21ftf _0912_ (
    .a(_0147_),
    .b(_0145_),
    .c(_0224_),
    .y(_0236_)
  );
  al_and3 _0913_ (
    .a(_0048_),
    .b(_0127_),
    .c(_0229_),
    .y(_0237_)
  );
  al_aoi21 _0914_ (
    .a(_0237_),
    .b(_0236_),
    .c(_0219_),
    .y(_0238_)
  );
  al_ao21ttf _0915_ (
    .a(_0235_),
    .b(_0238_),
    .c(N330),
    .y(_0239_)
  );
  al_aoi21 _0916_ (
    .a(_0219_),
    .b(_0232_),
    .c(_0239_),
    .y(_0240_)
  );
  al_ao21 _0917_ (
    .a(_0240_),
    .b(_0218_),
    .c(_0207_),
    .y(_0241_)
  );
  al_nand3 _0918_ (
    .a(_0207_),
    .b(_0240_),
    .c(_0218_),
    .y(_0242_)
  );
  al_ao21ttf _0919_ (
    .a(_0242_),
    .b(_0241_),
    .c(_0222_),
    .y(_0243_)
  );
  al_ao21ftf _0920_ (
    .a(_0222_),
    .b(_0207_),
    .c(_0243_),
    .y(_0244_)
  );
  al_inv _0921_ (
    .a(N1),
    .y(_0245_)
  );
  al_ao21 _0922_ (
    .a(N45),
    .b(_0093_),
    .c(_0245_),
    .y(_0246_)
  );
  al_and3ftt _0923_ (
    .a(N13),
    .b(N20),
    .c(N1),
    .y(_0247_)
  );
  al_and2ft _0924_ (
    .a(N41),
    .b(_0247_),
    .y(_0248_)
  );
  al_and2ft _0925_ (
    .a(_0213_),
    .b(_0212_),
    .y(_0249_)
  );
  al_and3 _0926_ (
    .a(_0249_),
    .b(_0217_),
    .c(_0240_),
    .y(_0250_)
  );
  al_nand3 _0927_ (
    .a(_0092_),
    .b(_0219_),
    .c(_0197_),
    .y(_0251_)
  );
  al_aoi21ftf _0928_ (
    .a(_0088_),
    .b(_0219_),
    .c(_0251_),
    .y(_0252_)
  );
  al_ao21 _0929_ (
    .a(_0217_),
    .b(_0240_),
    .c(_0249_),
    .y(_0253_)
  );
  al_ao21ftf _0930_ (
    .a(_0250_),
    .b(_0253_),
    .c(_0252_),
    .y(_0254_)
  );
  al_nand3fft _0931_ (
    .a(_0250_),
    .b(_0252_),
    .c(_0253_),
    .y(_0255_)
  );
  al_nand2 _0932_ (
    .a(_0111_),
    .b(_0240_),
    .y(_0256_)
  );
  al_nand3 _0933_ (
    .a(_0219_),
    .b(_0197_),
    .c(_0111_),
    .y(_0257_)
  );
  al_and3 _0934_ (
    .a(_0202_),
    .b(_0257_),
    .c(_0256_),
    .y(_0258_)
  );
  al_nand3 _0935_ (
    .a(_0258_),
    .b(_0255_),
    .c(_0254_),
    .y(_0259_)
  );
  al_ao21 _0936_ (
    .a(_0248_),
    .b(_0259_),
    .c(_0246_),
    .y(_0260_)
  );
  al_nand3 _0937_ (
    .a(_0242_),
    .b(_0241_),
    .c(_0222_),
    .y(_0261_)
  );
  al_aoi21 _0938_ (
    .a(_0242_),
    .b(_0241_),
    .c(_0222_),
    .y(_0262_)
  );
  al_nor3fft _0939_ (
    .a(_0248_),
    .b(_0261_),
    .c(_0262_),
    .y(_0263_)
  );
  al_nor2 _0940_ (
    .a(N13),
    .b(N33),
    .y(_0264_)
  );
  al_aoi21ftf _0941_ (
    .a(N169),
    .b(N20),
    .c(_0026_),
    .y(_0265_)
  );
  al_and3ftt _0942_ (
    .a(N179),
    .b(N200),
    .c(N20),
    .y(_0266_)
  );
  al_nand3ftt _0943_ (
    .a(N190),
    .b(N68),
    .c(_0266_),
    .y(_0267_)
  );
  al_and3ftt _0944_ (
    .a(N200),
    .b(N20),
    .c(N179),
    .y(_0268_)
  );
  al_and2ft _0945_ (
    .a(N190),
    .b(_0268_),
    .y(_0269_)
  );
  al_aoi21ttf _0946_ (
    .a(N97),
    .b(_0269_),
    .c(_0267_),
    .y(_0270_)
  );
  al_oai21 _0947_ (
    .a(N200),
    .b(N179),
    .c(N20),
    .y(_0271_)
  );
  al_aoi21ftf _0948_ (
    .a(N190),
    .b(N20),
    .c(_0271_),
    .y(_0272_)
  );
  al_nand2 _0949_ (
    .a(N77),
    .b(_0272_),
    .y(_0273_)
  );
  al_and3 _0950_ (
    .a(N200),
    .b(N20),
    .c(N179),
    .y(_0274_)
  );
  al_nand3 _0951_ (
    .a(N190),
    .b(N283),
    .c(_0274_),
    .y(_0275_)
  );
  al_nand3 _0952_ (
    .a(N116),
    .b(N190),
    .c(_0268_),
    .y(_0276_)
  );
  al_and3 _0953_ (
    .a(_0275_),
    .b(_0276_),
    .c(_0273_),
    .y(_0277_)
  );
  al_inv _0954_ (
    .a(N33),
    .y(_0278_)
  );
  al_and3ftt _0955_ (
    .a(N190),
    .b(N20),
    .c(_0271_),
    .y(_0279_)
  );
  al_aoi21 _0956_ (
    .a(N294),
    .b(_0279_),
    .c(_0278_),
    .y(_0280_)
  );
  al_and3ftt _0957_ (
    .a(N190),
    .b(N107),
    .c(_0274_),
    .y(_0281_)
  );
  al_and2 _0958_ (
    .a(N190),
    .b(_0266_),
    .y(_0282_)
  );
  al_aoi21 _0959_ (
    .a(N87),
    .b(_0282_),
    .c(_0281_),
    .y(_0283_)
  );
  al_nand3 _0960_ (
    .a(_0280_),
    .b(_0283_),
    .c(_0277_),
    .y(_0284_)
  );
  al_and3 _0961_ (
    .a(N190),
    .b(N150),
    .c(_0266_),
    .y(_0285_)
  );
  al_aoi21 _0962_ (
    .a(N125),
    .b(_0279_),
    .c(_0285_),
    .y(_0286_)
  );
  al_aoi21ttf _0963_ (
    .a(N143),
    .b(_0269_),
    .c(_0286_),
    .y(_0287_)
  );
  al_inv _0964_ (
    .a(N137),
    .y(_0288_)
  );
  al_and2ft _0965_ (
    .a(N190),
    .b(_0274_),
    .y(_0289_)
  );
  al_and2 _0966_ (
    .a(N190),
    .b(_0268_),
    .y(_0290_)
  );
  al_and3ftt _0967_ (
    .a(N190),
    .b(N50),
    .c(_0266_),
    .y(_0291_)
  );
  al_aoi21 _0968_ (
    .a(N132),
    .b(_0290_),
    .c(_0291_),
    .y(_0292_)
  );
  al_aoi21ftf _0969_ (
    .a(_0288_),
    .b(_0289_),
    .c(_0292_),
    .y(_0293_)
  );
  al_nand3 _0970_ (
    .a(N190),
    .b(N128),
    .c(_0274_),
    .y(_0294_)
  );
  al_nand2 _0971_ (
    .a(N159),
    .b(_0272_),
    .y(_0295_)
  );
  al_and3 _0972_ (
    .a(_0278_),
    .b(_0294_),
    .c(_0295_),
    .y(_0296_)
  );
  al_nand3 _0973_ (
    .a(_0296_),
    .b(_0293_),
    .c(_0287_),
    .y(_0297_)
  );
  al_ao21ftf _0974_ (
    .a(_0284_),
    .b(_0270_),
    .c(_0297_),
    .y(_0298_)
  );
  al_inv _0975_ (
    .a(N58),
    .y(_0299_)
  );
  al_aoi21ftt _0976_ (
    .a(N41),
    .b(_0247_),
    .c(_0246_),
    .y(_0300_)
  );
  al_nor2 _0977_ (
    .a(_0264_),
    .b(_0265_),
    .y(_0301_)
  );
  al_ao21ttf _0978_ (
    .a(_0299_),
    .b(_0301_),
    .c(_0300_),
    .y(_0302_)
  );
  al_aoi21 _0979_ (
    .a(_0265_),
    .b(_0298_),
    .c(_0302_),
    .y(_0303_)
  );
  al_oai21ftt _0980_ (
    .a(_0264_),
    .b(_0207_),
    .c(_0303_),
    .y(_0304_)
  );
  al_aoi21ftf _0981_ (
    .a(_0259_),
    .b(_0263_),
    .c(_0304_),
    .y(_0305_)
  );
  al_ao21ftf _0982_ (
    .a(_0244_),
    .b(_0260_),
    .c(_0305_),
    .y(N5102)
  );
  al_or3fft _0983_ (
    .a(_0254_),
    .b(_0255_),
    .c(_0244_),
    .y(_0306_)
  );
  al_and2 _0984_ (
    .a(_0202_),
    .b(_0257_),
    .y(_0307_)
  );
  al_and3ftt _0985_ (
    .a(_0246_),
    .b(_0256_),
    .c(_0307_),
    .y(_0308_)
  );
  al_inv _0986_ (
    .a(_0300_),
    .y(_0309_)
  );
  al_and3 _0987_ (
    .a(_0217_),
    .b(_0249_),
    .c(_0207_),
    .y(_0310_)
  );
  al_or2ft _0988_ (
    .a(_0203_),
    .b(_0069_),
    .y(_0311_)
  );
  al_ao21ttf _0989_ (
    .a(_0221_),
    .b(_0207_),
    .c(_0311_),
    .y(_0312_)
  );
  al_aoi21 _0990_ (
    .a(_0220_),
    .b(_0310_),
    .c(_0312_),
    .y(_0313_)
  );
  al_ao21 _0991_ (
    .a(_0035_),
    .b(_0029_),
    .c(_0203_),
    .y(_0314_)
  );
  al_nand3 _0992_ (
    .a(_0314_),
    .b(_0199_),
    .c(_0200_),
    .y(_0315_)
  );
  al_or3 _0993_ (
    .a(_0036_),
    .b(_0203_),
    .c(_0051_),
    .y(_0316_)
  );
  al_and2 _0994_ (
    .a(_0315_),
    .b(_0316_),
    .y(_0317_)
  );
  al_ao21 _0995_ (
    .a(_0240_),
    .b(_0310_),
    .c(_0317_),
    .y(_0318_)
  );
  al_and3 _0996_ (
    .a(_0240_),
    .b(_0317_),
    .c(_0310_),
    .y(_0319_)
  );
  al_ao21ftt _0997_ (
    .a(_0319_),
    .b(_0318_),
    .c(_0313_),
    .y(_0320_)
  );
  al_nand3ftt _0998_ (
    .a(_0319_),
    .b(_0318_),
    .c(_0313_),
    .y(_0321_)
  );
  al_and3 _0999_ (
    .a(_0309_),
    .b(_0321_),
    .c(_0320_),
    .y(_0322_)
  );
  al_ao21ttf _1000_ (
    .a(_0308_),
    .b(_0306_),
    .c(_0322_),
    .y(_0323_)
  );
  al_inv _1001_ (
    .a(N150),
    .y(_0324_)
  );
  al_and3ftt _1002_ (
    .a(N190),
    .b(N132),
    .c(_0274_),
    .y(_0325_)
  );
  al_aoi21 _1003_ (
    .a(N124),
    .b(_0279_),
    .c(_0325_),
    .y(_0326_)
  );
  al_ao21ftf _1004_ (
    .a(_0324_),
    .b(_0272_),
    .c(_0326_),
    .y(_0327_)
  );
  al_and3ftt _1005_ (
    .a(N190),
    .b(N159),
    .c(_0266_),
    .y(_0328_)
  );
  al_aoi21 _1006_ (
    .a(N128),
    .b(_0290_),
    .c(_0328_),
    .y(_0329_)
  );
  al_ao21ftf _1007_ (
    .a(_0288_),
    .b(_0269_),
    .c(_0329_),
    .y(_0330_)
  );
  al_nand3 _1008_ (
    .a(N190),
    .b(N125),
    .c(_0274_),
    .y(_0331_)
  );
  al_nand3 _1009_ (
    .a(N190),
    .b(N143),
    .c(_0266_),
    .y(_0332_)
  );
  al_and3 _1010_ (
    .a(_0278_),
    .b(_0332_),
    .c(_0331_),
    .y(_0333_)
  );
  al_or3ftt _1011_ (
    .a(_0333_),
    .b(_0330_),
    .c(_0327_),
    .y(_0334_)
  );
  al_nand3ftt _1012_ (
    .a(N190),
    .b(N58),
    .c(_0266_),
    .y(_0335_)
  );
  al_and3ftt _1013_ (
    .a(N190),
    .b(N97),
    .c(_0274_),
    .y(_0336_)
  );
  al_aoi21 _1014_ (
    .a(N107),
    .b(_0290_),
    .c(_0336_),
    .y(_0337_)
  );
  al_nand3 _1015_ (
    .a(N33),
    .b(_0335_),
    .c(_0337_),
    .y(_0338_)
  );
  al_inv _1016_ (
    .a(N283),
    .y(_0339_)
  );
  al_and3ftt _1017_ (
    .a(N190),
    .b(N87),
    .c(_0268_),
    .y(_0340_)
  );
  al_aoi21 _1018_ (
    .a(N77),
    .b(_0282_),
    .c(_0340_),
    .y(_0341_)
  );
  al_ao21ftf _1019_ (
    .a(_0339_),
    .b(_0279_),
    .c(_0341_),
    .y(_0342_)
  );
  al_inv _1020_ (
    .a(N116),
    .y(_0343_)
  );
  al_and2 _1021_ (
    .a(N190),
    .b(_0274_),
    .y(_0344_)
  );
  al_nand2 _1022_ (
    .a(N68),
    .b(_0272_),
    .y(_0345_)
  );
  al_ao21ftf _1023_ (
    .a(_0343_),
    .b(_0344_),
    .c(_0345_),
    .y(_0346_)
  );
  al_or3 _1024_ (
    .a(_0346_),
    .b(_0338_),
    .c(_0342_),
    .y(_0347_)
  );
  al_nand3ftt _1025_ (
    .a(N41),
    .b(_0347_),
    .c(_0334_),
    .y(_0348_)
  );
  al_nand2 _1026_ (
    .a(N41),
    .b(N50),
    .y(_0349_)
  );
  al_nand3 _1027_ (
    .a(_0265_),
    .b(_0349_),
    .c(_0348_),
    .y(_0350_)
  );
  al_or3 _1028_ (
    .a(N50),
    .b(_0264_),
    .c(_0265_),
    .y(_0351_)
  );
  al_and3 _1029_ (
    .a(_0300_),
    .b(_0351_),
    .c(_0350_),
    .y(_0352_)
  );
  al_aoi21ttf _1030_ (
    .a(_0264_),
    .b(_0317_),
    .c(_0352_),
    .y(_0353_)
  );
  al_and3fft _1031_ (
    .a(_0353_),
    .b(N5102),
    .c(_0323_),
    .y(_0354_)
  );
  al_or3fft _1032_ (
    .a(_0264_),
    .b(_0216_),
    .c(_0215_),
    .y(_0355_)
  );
  al_and3 _1033_ (
    .a(N190),
    .b(N137),
    .c(_0274_),
    .y(_0356_)
  );
  al_aoi21 _1034_ (
    .a(N58),
    .b(_0272_),
    .c(_0356_),
    .y(_0357_)
  );
  al_aoi21ttf _1035_ (
    .a(N132),
    .b(_0279_),
    .c(_0357_),
    .y(_0358_)
  );
  al_and3 _1036_ (
    .a(N50),
    .b(N190),
    .c(_0266_),
    .y(_0359_)
  );
  al_aoi21 _1037_ (
    .a(N143),
    .b(_0290_),
    .c(_0359_),
    .y(_0360_)
  );
  al_aoi21ttf _1038_ (
    .a(N159),
    .b(_0269_),
    .c(_0360_),
    .y(_0361_)
  );
  al_nand3ftt _1039_ (
    .a(N190),
    .b(N150),
    .c(_0274_),
    .y(_0362_)
  );
  al_and3 _1040_ (
    .a(_0278_),
    .b(_0267_),
    .c(_0362_),
    .y(_0363_)
  );
  al_nand3 _1041_ (
    .a(_0363_),
    .b(_0361_),
    .c(_0358_),
    .y(_0364_)
  );
  al_inv _1042_ (
    .a(N303),
    .y(_0365_)
  );
  al_and3ftt _1043_ (
    .a(N190),
    .b(N283),
    .c(_0274_),
    .y(_0366_)
  );
  al_aoi21 _1044_ (
    .a(N116),
    .b(_0269_),
    .c(_0366_),
    .y(_0367_)
  );
  al_aoi21ftf _1045_ (
    .a(_0365_),
    .b(_0344_),
    .c(_0367_),
    .y(_0368_)
  );
  al_aoi21 _1046_ (
    .a(N311),
    .b(_0279_),
    .c(_0278_),
    .y(_0369_)
  );
  al_nand3 _1047_ (
    .a(N190),
    .b(N294),
    .c(_0268_),
    .y(_0370_)
  );
  al_aoi21ttf _1048_ (
    .a(N107),
    .b(_0282_),
    .c(_0370_),
    .y(_0371_)
  );
  al_nand2 _1049_ (
    .a(N97),
    .b(_0272_),
    .y(_0372_)
  );
  al_nand3ftt _1050_ (
    .a(N190),
    .b(N87),
    .c(_0266_),
    .y(_0373_)
  );
  al_and3 _1051_ (
    .a(_0373_),
    .b(_0372_),
    .c(_0371_),
    .y(_0374_)
  );
  al_nand3 _1052_ (
    .a(_0369_),
    .b(_0374_),
    .c(_0368_),
    .y(_0375_)
  );
  al_ao21ttf _1053_ (
    .a(_0375_),
    .b(_0364_),
    .c(_0265_),
    .y(_0376_)
  );
  al_aoi21ftf _1054_ (
    .a(N77),
    .b(_0301_),
    .c(_0300_),
    .y(_0377_)
  );
  al_nand3 _1055_ (
    .a(_0376_),
    .b(_0377_),
    .c(_0355_),
    .y(_0378_)
  );
  al_and2 _1056_ (
    .a(_0217_),
    .b(_0240_),
    .y(_0379_)
  );
  al_ao21 _1057_ (
    .a(_0219_),
    .b(_0197_),
    .c(_0217_),
    .y(_0380_)
  );
  al_ao21 _1058_ (
    .a(_0251_),
    .b(_0380_),
    .c(_0240_),
    .y(_0381_)
  );
  al_nand3fft _1059_ (
    .a(_0379_),
    .b(_0300_),
    .c(_0381_),
    .y(_0382_)
  );
  al_and2 _1060_ (
    .a(_0378_),
    .b(_0382_),
    .y(_0383_)
  );
  al_and2 _1061_ (
    .a(_0255_),
    .b(_0254_),
    .y(_0384_)
  );
  al_nand2 _1062_ (
    .a(_0384_),
    .b(_0260_),
    .y(_0385_)
  );
  al_ao21ftf _1063_ (
    .a(_0213_),
    .b(_0212_),
    .c(_0264_),
    .y(_0386_)
  );
  al_and3 _1064_ (
    .a(N190),
    .b(N159),
    .c(_0266_),
    .y(_0387_)
  );
  al_aoi21 _1065_ (
    .a(N137),
    .b(_0290_),
    .c(_0387_),
    .y(_0388_)
  );
  al_aoi21ttf _1066_ (
    .a(N128),
    .b(_0279_),
    .c(_0388_),
    .y(_0389_)
  );
  al_inv _1067_ (
    .a(N50),
    .y(_0390_)
  );
  al_and3ftt _1068_ (
    .a(N190),
    .b(N143),
    .c(_0274_),
    .y(_0391_)
  );
  al_ao21 _1069_ (
    .a(N150),
    .b(_0269_),
    .c(_0391_),
    .y(_0392_)
  );
  al_ao21ftt _1070_ (
    .a(_0390_),
    .b(_0272_),
    .c(_0392_),
    .y(_0393_)
  );
  al_nand3 _1071_ (
    .a(N190),
    .b(N132),
    .c(_0274_),
    .y(_0394_)
  );
  al_and3 _1072_ (
    .a(_0278_),
    .b(_0335_),
    .c(_0394_),
    .y(_0395_)
  );
  al_or3fft _1073_ (
    .a(_0395_),
    .b(_0389_),
    .c(_0393_),
    .y(_0396_)
  );
  al_and3 _1074_ (
    .a(N97),
    .b(N190),
    .c(_0266_),
    .y(_0397_)
  );
  al_aoi21 _1075_ (
    .a(N303),
    .b(_0279_),
    .c(_0397_),
    .y(_0398_)
  );
  al_ao21ftf _1076_ (
    .a(_0339_),
    .b(_0290_),
    .c(_0398_),
    .y(_0399_)
  );
  al_and2 _1077_ (
    .a(N87),
    .b(_0272_),
    .y(_0400_)
  );
  al_and3ftt _1078_ (
    .a(N190),
    .b(N77),
    .c(_0266_),
    .y(_0401_)
  );
  al_nand3 _1079_ (
    .a(N190),
    .b(N294),
    .c(_0274_),
    .y(_0402_)
  );
  al_or3ftt _1080_ (
    .a(_0402_),
    .b(_0401_),
    .c(_0400_),
    .y(_0403_)
  );
  al_aoi21 _1081_ (
    .a(N107),
    .b(_0269_),
    .c(_0278_),
    .y(_0404_)
  );
  al_ao21ftf _1082_ (
    .a(_0343_),
    .b(_0289_),
    .c(_0404_),
    .y(_0405_)
  );
  al_or3 _1083_ (
    .a(_0403_),
    .b(_0405_),
    .c(_0399_),
    .y(_0406_)
  );
  al_ao21ttf _1084_ (
    .a(_0406_),
    .b(_0396_),
    .c(_0265_),
    .y(_0407_)
  );
  al_aoi21ftf _1085_ (
    .a(N68),
    .b(_0301_),
    .c(_0300_),
    .y(_0408_)
  );
  al_nand3 _1086_ (
    .a(_0407_),
    .b(_0408_),
    .c(_0386_),
    .y(_0409_)
  );
  al_inv _1087_ (
    .a(_0248_),
    .y(_0410_)
  );
  al_nand3 _1088_ (
    .a(_0202_),
    .b(_0257_),
    .c(_0256_),
    .y(_0411_)
  );
  al_nand3fft _1089_ (
    .a(_0410_),
    .b(_0411_),
    .c(_0259_),
    .y(_0412_)
  );
  al_and2 _1090_ (
    .a(_0409_),
    .b(_0412_),
    .y(_0413_)
  );
  al_and3 _1091_ (
    .a(_0383_),
    .b(_0413_),
    .c(_0385_),
    .y(_0414_)
  );
  al_ao21ftt _1092_ (
    .a(_0219_),
    .b(_0178_),
    .c(_0231_),
    .y(_0415_)
  );
  al_nand3 _1093_ (
    .a(_0178_),
    .b(_0210_),
    .c(_0231_),
    .y(_0416_)
  );
  al_or3 _1094_ (
    .a(N13),
    .b(N20),
    .c(N33),
    .y(_0417_)
  );
  al_aoi21 _1095_ (
    .a(_0416_),
    .b(_0415_),
    .c(_0417_),
    .y(_0418_)
  );
  al_and3ftt _1096_ (
    .a(N190),
    .b(N283),
    .c(_0266_),
    .y(_0419_)
  );
  al_aoi21 _1097_ (
    .a(N329),
    .b(_0279_),
    .c(_0419_),
    .y(_0420_)
  );
  al_ao21ttf _1098_ (
    .a(N294),
    .b(_0272_),
    .c(_0420_),
    .y(_0421_)
  );
  al_and3 _1099_ (
    .a(N190),
    .b(N326),
    .c(_0274_),
    .y(_0422_)
  );
  al_aoi21 _1100_ (
    .a(N303),
    .b(_0282_),
    .c(_0422_),
    .y(_0423_)
  );
  al_ao21ttf _1101_ (
    .a(N322),
    .b(_0290_),
    .c(_0423_),
    .y(_0424_)
  );
  al_nand3ftt _1102_ (
    .a(N190),
    .b(N311),
    .c(_0268_),
    .y(_0425_)
  );
  al_nand3ftt _1103_ (
    .a(N190),
    .b(N317),
    .c(_0274_),
    .y(_0426_)
  );
  al_and3 _1104_ (
    .a(N33),
    .b(_0425_),
    .c(_0426_),
    .y(_0427_)
  );
  al_or3ftt _1105_ (
    .a(_0427_),
    .b(_0424_),
    .c(_0421_),
    .y(_0428_)
  );
  al_nand3ftt _1106_ (
    .a(N190),
    .b(N107),
    .c(_0266_),
    .y(_0429_)
  );
  al_ao21ttf _1107_ (
    .a(N50),
    .b(_0344_),
    .c(_0429_),
    .y(_0430_)
  );
  al_and3ftt _1108_ (
    .a(N190),
    .b(N77),
    .c(_0268_),
    .y(_0431_)
  );
  al_aoi21 _1109_ (
    .a(N58),
    .b(_0290_),
    .c(_0431_),
    .y(_0432_)
  );
  al_ao21ttf _1110_ (
    .a(N68),
    .b(_0289_),
    .c(_0432_),
    .y(_0433_)
  );
  al_and2 _1111_ (
    .a(N159),
    .b(_0279_),
    .y(_0434_)
  );
  al_aoi21 _1112_ (
    .a(N87),
    .b(_0282_),
    .c(N33),
    .y(_0435_)
  );
  al_and3ftt _1113_ (
    .a(_0434_),
    .b(_0372_),
    .c(_0435_),
    .y(_0436_)
  );
  al_nand3fft _1114_ (
    .a(_0430_),
    .b(_0433_),
    .c(_0436_),
    .y(_0437_)
  );
  al_ao21ttf _1115_ (
    .a(_0437_),
    .b(_0428_),
    .c(_0265_),
    .y(_0438_)
  );
  al_nor2ft _1116_ (
    .a(_0417_),
    .b(_0265_),
    .y(_0439_)
  );
  al_or3fft _1117_ (
    .a(N45),
    .b(_0012_),
    .c(_0013_),
    .y(_0440_)
  );
  al_and2 _1118_ (
    .a(N33),
    .b(_0247_),
    .y(_0441_)
  );
  al_nand3ftt _1119_ (
    .a(N45),
    .b(N50),
    .c(_0062_),
    .y(_0442_)
  );
  al_nand3 _1120_ (
    .a(_0441_),
    .b(_0442_),
    .c(_0440_),
    .y(_0443_)
  );
  al_nand3ftt _1121_ (
    .a(N33),
    .b(_0247_),
    .c(N1947),
    .y(_0444_)
  );
  al_aoi21ftf _1122_ (
    .a(_0247_),
    .b(_0343_),
    .c(_0444_),
    .y(_0445_)
  );
  al_ao21ttf _1123_ (
    .a(_0445_),
    .b(_0443_),
    .c(_0439_),
    .y(_0446_)
  );
  al_and3 _1124_ (
    .a(_0300_),
    .b(_0446_),
    .c(_0438_),
    .y(_0447_)
  );
  al_ao21 _1125_ (
    .a(_0416_),
    .b(_0415_),
    .c(N330),
    .y(_0448_)
  );
  al_nand3 _1126_ (
    .a(N330),
    .b(_0416_),
    .c(_0415_),
    .y(_0449_)
  );
  al_nand3 _1127_ (
    .a(_0309_),
    .b(_0449_),
    .c(_0448_),
    .y(_0450_)
  );
  al_aoi21ftf _1128_ (
    .a(_0418_),
    .b(_0447_),
    .c(_0450_),
    .y(_0451_)
  );
  al_nand2 _1129_ (
    .a(_0210_),
    .b(_0170_),
    .y(_0452_)
  );
  al_ao21ttf _1130_ (
    .a(_0171_),
    .b(_0190_),
    .c(_0452_),
    .y(_0453_)
  );
  al_nand3ftt _1131_ (
    .a(_0452_),
    .b(_0171_),
    .c(_0190_),
    .y(_0454_)
  );
  al_and2 _1132_ (
    .a(_0454_),
    .b(_0453_),
    .y(_0455_)
  );
  al_nor2 _1133_ (
    .a(N107),
    .b(_0247_),
    .y(_0456_)
  );
  al_nand3fft _1134_ (
    .a(N116),
    .b(N87),
    .c(_0014_),
    .y(_0457_)
  );
  al_and3 _1135_ (
    .a(_0278_),
    .b(_0247_),
    .c(_0457_),
    .y(_0458_)
  );
  al_or3fft _1136_ (
    .a(N45),
    .b(_0004_),
    .c(_0003_),
    .y(_0459_)
  );
  al_ao21 _1137_ (
    .a(_0441_),
    .b(_0459_),
    .c(_0458_),
    .y(_0460_)
  );
  al_and3fft _1138_ (
    .a(N45),
    .b(N50),
    .c(N58),
    .y(_0461_)
  );
  al_or3fft _1139_ (
    .a(_0010_),
    .b(_0461_),
    .c(_0457_),
    .y(_0462_)
  );
  al_aoi21 _1140_ (
    .a(_0462_),
    .b(_0460_),
    .c(_0456_),
    .y(_0463_)
  );
  al_and3 _1141_ (
    .a(N190),
    .b(N317),
    .c(_0268_),
    .y(_0464_)
  );
  al_aoi21 _1142_ (
    .a(N283),
    .b(_0272_),
    .c(_0464_),
    .y(_0465_)
  );
  al_ao21ttf _1143_ (
    .a(N326),
    .b(_0279_),
    .c(_0465_),
    .y(_0466_)
  );
  al_and3ftt _1144_ (
    .a(N190),
    .b(N311),
    .c(_0274_),
    .y(_0467_)
  );
  al_aoi21 _1145_ (
    .a(N294),
    .b(_0282_),
    .c(_0467_),
    .y(_0468_)
  );
  al_ao21ftf _1146_ (
    .a(_0365_),
    .b(_0269_),
    .c(_0468_),
    .y(_0469_)
  );
  al_nand3ftt _1147_ (
    .a(N190),
    .b(N116),
    .c(_0266_),
    .y(_0470_)
  );
  al_nand3 _1148_ (
    .a(N190),
    .b(N322),
    .c(_0274_),
    .y(_0471_)
  );
  al_and3 _1149_ (
    .a(N33),
    .b(_0470_),
    .c(_0471_),
    .y(_0472_)
  );
  al_or3ftt _1150_ (
    .a(_0472_),
    .b(_0469_),
    .c(_0466_),
    .y(_0473_)
  );
  al_and3ftt _1151_ (
    .a(N190),
    .b(N68),
    .c(_0268_),
    .y(_0474_)
  );
  al_aoi21 _1152_ (
    .a(N50),
    .b(_0290_),
    .c(_0474_),
    .y(_0475_)
  );
  al_ao21ftf _1153_ (
    .a(_0299_),
    .b(_0289_),
    .c(_0475_),
    .y(_0476_)
  );
  al_and3ftt _1154_ (
    .a(N190),
    .b(N97),
    .c(_0266_),
    .y(_0477_)
  );
  al_aoi21 _1155_ (
    .a(N159),
    .b(_0344_),
    .c(_0477_),
    .y(_0478_)
  );
  al_aoi21 _1156_ (
    .a(N77),
    .b(_0282_),
    .c(N33),
    .y(_0479_)
  );
  al_aoi21ftt _1157_ (
    .a(_0324_),
    .b(_0279_),
    .c(_0400_),
    .y(_0480_)
  );
  al_and3 _1158_ (
    .a(_0478_),
    .b(_0479_),
    .c(_0480_),
    .y(_0481_)
  );
  al_ao21ftf _1159_ (
    .a(_0476_),
    .b(_0481_),
    .c(_0473_),
    .y(_0482_)
  );
  al_aoi21 _1160_ (
    .a(_0265_),
    .b(_0482_),
    .c(_0309_),
    .y(_0483_)
  );
  al_aoi21ftf _1161_ (
    .a(_0463_),
    .b(_0439_),
    .c(_0483_),
    .y(_0484_)
  );
  al_oai21 _1162_ (
    .a(_0417_),
    .b(_0455_),
    .c(_0484_),
    .y(_0485_)
  );
  al_and3 _1163_ (
    .a(N330),
    .b(_0416_),
    .c(_0415_),
    .y(_0486_)
  );
  al_nand3 _1164_ (
    .a(_0453_),
    .b(_0454_),
    .c(_0486_),
    .y(_0487_)
  );
  al_nor2 _1165_ (
    .a(_0210_),
    .b(_0187_),
    .y(_0488_)
  );
  al_nand3ftt _1166_ (
    .a(_0488_),
    .b(_0454_),
    .c(_0453_),
    .y(_0489_)
  );
  al_nand3ftt _1167_ (
    .a(_0187_),
    .b(_0219_),
    .c(_0226_),
    .y(_0490_)
  );
  al_nand3 _1168_ (
    .a(_0489_),
    .b(_0490_),
    .c(_0449_),
    .y(_0491_)
  );
  al_nand3 _1169_ (
    .a(_0246_),
    .b(_0491_),
    .c(_0487_),
    .y(_0492_)
  );
  al_and2 _1170_ (
    .a(_0485_),
    .b(_0492_),
    .y(_0493_)
  );
  al_ao21ftt _1171_ (
    .a(_0210_),
    .b(_0197_),
    .c(_0240_),
    .y(_0494_)
  );
  al_ao21ttf _1172_ (
    .a(_0487_),
    .b(_0491_),
    .c(_0494_),
    .y(_0495_)
  );
  al_or3fft _1173_ (
    .a(_0487_),
    .b(_0491_),
    .c(_0494_),
    .y(_0496_)
  );
  al_nand3 _1174_ (
    .a(_0248_),
    .b(_0495_),
    .c(_0496_),
    .y(_0497_)
  );
  al_and3 _1175_ (
    .a(_0451_),
    .b(_0493_),
    .c(_0497_),
    .y(_0498_)
  );
  al_nor2 _1176_ (
    .a(_0210_),
    .b(_0191_),
    .y(_0499_)
  );
  al_nand3ftt _1177_ (
    .a(_0137_),
    .b(_0151_),
    .c(_0152_),
    .y(_0500_)
  );
  al_nand2 _1178_ (
    .a(_0210_),
    .b(_0137_),
    .y(_0501_)
  );
  al_and3 _1179_ (
    .a(_0501_),
    .b(_0500_),
    .c(_0149_),
    .y(_0502_)
  );
  al_ao21 _1180_ (
    .a(_0500_),
    .b(_0149_),
    .c(_0501_),
    .y(_0503_)
  );
  al_nand2ft _1181_ (
    .a(_0502_),
    .b(_0503_),
    .y(_0504_)
  );
  al_nand3 _1182_ (
    .a(_0504_),
    .b(_0455_),
    .c(_0486_),
    .y(_0505_)
  );
  al_ao21 _1183_ (
    .a(_0455_),
    .b(_0486_),
    .c(_0504_),
    .y(_0506_)
  );
  al_nand3 _1184_ (
    .a(_0499_),
    .b(_0505_),
    .c(_0506_),
    .y(_0507_)
  );
  al_ao21 _1185_ (
    .a(_0505_),
    .b(_0506_),
    .c(_0499_),
    .y(_0508_)
  );
  al_or3fft _1186_ (
    .a(_0507_),
    .b(_0508_),
    .c(_0496_),
    .y(_0509_)
  );
  al_nor2 _1187_ (
    .a(_0246_),
    .b(_0494_),
    .y(_0510_)
  );
  al_oai21ftf _1188_ (
    .a(_0500_),
    .b(_0171_),
    .c(_0195_),
    .y(_0511_)
  );
  al_nand2 _1189_ (
    .a(_0219_),
    .b(_0511_),
    .y(_0512_)
  );
  al_and3 _1190_ (
    .a(_0149_),
    .b(_0500_),
    .c(_0488_),
    .y(_0513_)
  );
  al_nand3 _1191_ (
    .a(_0453_),
    .b(_0454_),
    .c(_0513_),
    .y(_0514_)
  );
  al_aoi21ftf _1192_ (
    .a(_0120_),
    .b(_0210_),
    .c(_0130_),
    .y(_0515_)
  );
  al_or3fft _1193_ (
    .a(_0192_),
    .b(_0210_),
    .c(_0130_),
    .y(_0516_)
  );
  al_and2ft _1194_ (
    .a(_0515_),
    .b(_0516_),
    .y(_0517_)
  );
  al_and3 _1195_ (
    .a(_0512_),
    .b(_0517_),
    .c(_0514_),
    .y(_0518_)
  );
  al_ao21 _1196_ (
    .a(_0512_),
    .b(_0514_),
    .c(_0517_),
    .y(_0519_)
  );
  al_nand3fft _1197_ (
    .a(_0518_),
    .b(_0505_),
    .c(_0519_),
    .y(_0520_)
  );
  al_ao21ftf _1198_ (
    .a(_0518_),
    .b(_0519_),
    .c(_0505_),
    .y(_0521_)
  );
  al_nand3 _1199_ (
    .a(_0309_),
    .b(_0520_),
    .c(_0521_),
    .y(_0522_)
  );
  al_ao21 _1200_ (
    .a(_0510_),
    .b(_0509_),
    .c(_0522_),
    .y(_0523_)
  );
  al_nand3fft _1201_ (
    .a(_0417_),
    .b(_0515_),
    .c(_0516_),
    .y(_0524_)
  );
  al_and3 _1202_ (
    .a(N190),
    .b(N143),
    .c(_0274_),
    .y(_0525_)
  );
  al_aoi21 _1203_ (
    .a(N58),
    .b(_0282_),
    .c(_0525_),
    .y(_0526_)
  );
  al_and3ftt _1204_ (
    .a(N190),
    .b(N50),
    .c(_0268_),
    .y(_0527_)
  );
  al_aoi21 _1205_ (
    .a(N137),
    .b(_0279_),
    .c(_0527_),
    .y(_0528_)
  );
  al_aoi21 _1206_ (
    .a(N159),
    .b(_0289_),
    .c(_0401_),
    .y(_0529_)
  );
  al_aoi21ftf _1207_ (
    .a(_0324_),
    .b(_0290_),
    .c(_0345_),
    .y(_0530_)
  );
  al_and3 _1208_ (
    .a(_0528_),
    .b(_0529_),
    .c(_0530_),
    .y(_0531_)
  );
  al_ao21 _1209_ (
    .a(_0526_),
    .b(_0531_),
    .c(N33),
    .y(_0532_)
  );
  al_nand3 _1210_ (
    .a(N190),
    .b(N311),
    .c(_0274_),
    .y(_0533_)
  );
  al_aoi21ttf _1211_ (
    .a(N107),
    .b(_0272_),
    .c(_0533_),
    .y(_0534_)
  );
  al_nand3ftt _1212_ (
    .a(N190),
    .b(N283),
    .c(_0268_),
    .y(_0535_)
  );
  al_aoi21ttf _1213_ (
    .a(N317),
    .b(_0279_),
    .c(_0535_),
    .y(_0536_)
  );
  al_aoi21 _1214_ (
    .a(N303),
    .b(_0290_),
    .c(_0477_),
    .y(_0537_)
  );
  al_nand3ftt _1215_ (
    .a(N190),
    .b(N294),
    .c(_0274_),
    .y(_0538_)
  );
  al_ao21ttf _1216_ (
    .a(N116),
    .b(_0282_),
    .c(_0538_),
    .y(_0539_)
  );
  al_and3ftt _1217_ (
    .a(_0539_),
    .b(_0536_),
    .c(_0537_),
    .y(_0540_)
  );
  al_ao21 _1218_ (
    .a(_0534_),
    .b(_0540_),
    .c(_0278_),
    .y(_0541_)
  );
  al_nand3 _1219_ (
    .a(_0265_),
    .b(_0541_),
    .c(_0532_),
    .y(_0542_)
  );
  al_oai21 _1220_ (
    .a(_0641_),
    .b(_0642_),
    .c(_0441_),
    .y(_0543_)
  );
  al_aoi21ftf _1221_ (
    .a(_0247_),
    .b(N87),
    .c(_0439_),
    .y(_0544_)
  );
  al_aoi21 _1222_ (
    .a(_0544_),
    .b(_0543_),
    .c(_0309_),
    .y(_0545_)
  );
  al_and3 _1223_ (
    .a(_0542_),
    .b(_0545_),
    .c(_0524_),
    .y(_0546_)
  );
  al_nand2ft _1224_ (
    .a(_0546_),
    .b(_0523_),
    .y(N5045)
  );
  al_ao21ttf _1225_ (
    .a(_0507_),
    .b(_0508_),
    .c(_0496_),
    .y(_0547_)
  );
  al_nand3 _1226_ (
    .a(_0248_),
    .b(_0509_),
    .c(_0547_),
    .y(_0548_)
  );
  al_nand3 _1227_ (
    .a(_0246_),
    .b(_0507_),
    .c(_0508_),
    .y(_0549_)
  );
  al_nand3fft _1228_ (
    .a(_0417_),
    .b(_0502_),
    .c(_0503_),
    .y(_0550_)
  );
  al_and3ftt _1229_ (
    .a(N190),
    .b(N50),
    .c(_0274_),
    .y(_0551_)
  );
  al_aoi21 _1230_ (
    .a(N150),
    .b(_0344_),
    .c(_0551_),
    .y(_0552_)
  );
  al_and3 _1231_ (
    .a(N68),
    .b(N190),
    .c(_0266_),
    .y(_0553_)
  );
  al_aoi21 _1232_ (
    .a(N143),
    .b(_0279_),
    .c(_0553_),
    .y(_0554_)
  );
  al_and3ftt _1233_ (
    .a(N190),
    .b(N58),
    .c(_0268_),
    .y(_0555_)
  );
  al_aoi21 _1234_ (
    .a(N159),
    .b(_0290_),
    .c(_0555_),
    .y(_0556_)
  );
  al_and3 _1235_ (
    .a(_0373_),
    .b(_0273_),
    .c(_0556_),
    .y(_0557_)
  );
  al_and3 _1236_ (
    .a(_0552_),
    .b(_0554_),
    .c(_0557_),
    .y(_0558_)
  );
  al_and3 _1237_ (
    .a(N190),
    .b(N317),
    .c(_0274_),
    .y(_0559_)
  );
  al_aoi21 _1238_ (
    .a(N294),
    .b(_0269_),
    .c(_0559_),
    .y(_0560_)
  );
  al_aoi21ftf _1239_ (
    .a(_0365_),
    .b(_0289_),
    .c(_0560_),
    .y(_0561_)
  );
  al_and3 _1240_ (
    .a(N190),
    .b(N283),
    .c(_0266_),
    .y(_0562_)
  );
  al_aoi21 _1241_ (
    .a(N322),
    .b(_0279_),
    .c(_0562_),
    .y(_0563_)
  );
  al_aoi21ftf _1242_ (
    .a(_0343_),
    .b(_0272_),
    .c(_0563_),
    .y(_0564_)
  );
  al_nand3 _1243_ (
    .a(N190),
    .b(N311),
    .c(_0268_),
    .y(_0565_)
  );
  al_and3 _1244_ (
    .a(N33),
    .b(_0565_),
    .c(_0429_),
    .y(_0566_)
  );
  al_nand3 _1245_ (
    .a(_0566_),
    .b(_0561_),
    .c(_0564_),
    .y(_0567_)
  );
  al_ao21ttf _1246_ (
    .a(_0278_),
    .b(_0558_),
    .c(_0567_),
    .y(_0568_)
  );
  al_oai21ftt _1247_ (
    .a(_0020_),
    .b(_0019_),
    .c(_0441_),
    .y(_0569_)
  );
  al_or2ft _1248_ (
    .a(N97),
    .b(_0247_),
    .y(_0570_)
  );
  al_and3 _1249_ (
    .a(_0439_),
    .b(_0570_),
    .c(_0569_),
    .y(_0571_)
  );
  al_aoi21 _1250_ (
    .a(_0265_),
    .b(_0568_),
    .c(_0571_),
    .y(_0572_)
  );
  al_nand3 _1251_ (
    .a(_0300_),
    .b(_0572_),
    .c(_0550_),
    .y(_0573_)
  );
  al_nand3 _1252_ (
    .a(_0549_),
    .b(_0573_),
    .c(_0548_),
    .y(N5078)
  );
  al_nor3ftt _1253_ (
    .a(_0498_),
    .b(N5078),
    .c(N5045),
    .y(_0574_)
  );
  al_nand3 _1254_ (
    .a(_0574_),
    .b(_0414_),
    .c(_0354_),
    .y(N5192)
  );
  al_ao21ftf _1255_ (
    .a(_0244_),
    .b(_0384_),
    .c(_0308_),
    .y(_0575_)
  );
  al_ao21 _1256_ (
    .a(_0322_),
    .b(_0575_),
    .c(_0353_),
    .y(N5120)
  );
  al_or3 _1257_ (
    .a(N343),
    .b(N5102),
    .c(N5120),
    .y(_0576_)
  );
  al_nand3 _1258_ (
    .a(N213),
    .b(_0576_),
    .c(N5192),
    .y(N5231)
  );
  al_or3ftt _1259_ (
    .a(_0323_),
    .b(_0353_),
    .c(N5102),
    .y(_0577_)
  );
  al_aoi21ftf _1260_ (
    .a(_0353_),
    .b(_0323_),
    .c(N5102),
    .y(_0578_)
  );
  al_and2ft _1261_ (
    .a(_0578_),
    .b(_0577_),
    .y(_0579_)
  );
  al_ao21 _1262_ (
    .a(_0413_),
    .b(_0385_),
    .c(_0383_),
    .y(_0580_)
  );
  al_nand2ft _1263_ (
    .a(_0414_),
    .b(_0580_),
    .y(_0581_)
  );
  al_ao21 _1264_ (
    .a(_0493_),
    .b(_0497_),
    .c(_0451_),
    .y(_0582_)
  );
  al_nand2ft _1265_ (
    .a(_0498_),
    .b(_0582_),
    .y(_0583_)
  );
  al_aoi21 _1266_ (
    .a(_0510_),
    .b(_0509_),
    .c(_0522_),
    .y(_0584_)
  );
  al_nand3fft _1267_ (
    .a(_0584_),
    .b(_0546_),
    .c(N5078),
    .y(_0585_)
  );
  al_ao21ftt _1268_ (
    .a(_0546_),
    .b(_0523_),
    .c(N5078),
    .y(_0586_)
  );
  al_nand3 _1269_ (
    .a(_0583_),
    .b(_0585_),
    .c(_0586_),
    .y(_0587_)
  );
  al_or3 _1270_ (
    .a(_0584_),
    .b(_0546_),
    .c(N5078),
    .y(_0588_)
  );
  al_and2ft _1271_ (
    .a(_0498_),
    .b(_0582_),
    .y(_0589_)
  );
  al_ao21ftf _1272_ (
    .a(_0546_),
    .b(_0523_),
    .c(N5078),
    .y(_0590_)
  );
  al_nand3 _1273_ (
    .a(_0589_),
    .b(_0590_),
    .c(_0588_),
    .y(_0591_)
  );
  al_nand3 _1274_ (
    .a(_0587_),
    .b(_0591_),
    .c(_0581_),
    .y(_0592_)
  );
  al_and2ft _1275_ (
    .a(_0414_),
    .b(_0580_),
    .y(_0593_)
  );
  al_nand3 _1276_ (
    .a(_0583_),
    .b(_0590_),
    .c(_0588_),
    .y(_0594_)
  );
  al_nand3 _1277_ (
    .a(_0589_),
    .b(_0585_),
    .c(_0586_),
    .y(_0595_)
  );
  al_nand3 _1278_ (
    .a(_0594_),
    .b(_0595_),
    .c(_0593_),
    .y(_0596_)
  );
  al_and3ftt _1279_ (
    .a(_0579_),
    .b(_0592_),
    .c(_0596_),
    .y(_0597_)
  );
  al_nand3 _1280_ (
    .a(_0594_),
    .b(_0595_),
    .c(_0581_),
    .y(_0598_)
  );
  al_nand3 _1281_ (
    .a(_0587_),
    .b(_0591_),
    .c(_0593_),
    .y(_0599_)
  );
  al_nand3 _1282_ (
    .a(_0579_),
    .b(_0598_),
    .c(_0599_),
    .y(_0600_)
  );
  al_nand2ft _1283_ (
    .a(_0597_),
    .b(_0600_),
    .y(N5361)
  );
  al_nor2 _1284_ (
    .a(N77),
    .b(_0032_),
    .y(N1713)
  );
  al_and2ft _1285_ (
    .a(_0232_),
    .b(_0111_),
    .y(N4028)
  );
  al_ao21 _1286_ (
    .a(_0455_),
    .b(_0486_),
    .c(_0499_),
    .y(N4589)
  );
  al_and3fft _1287_ (
    .a(N116),
    .b(_0116_),
    .c(N1),
    .y(_0601_)
  );
  al_mux2l _1288_ (
    .a(_0623_),
    .b(_0601_),
    .s(_0248_),
    .y(_0602_)
  );
  al_ao21 _1289_ (
    .a(_0245_),
    .b(_0494_),
    .c(_0602_),
    .y(N4667)
  );
  al_inv _1290_ (
    .a(_0451_),
    .y(N4815)
  );
  al_inv _1291_ (
    .a(_0383_),
    .y(N4944)
  );
  al_or3fft _1292_ (
    .a(_0202_),
    .b(_0257_),
    .c(_0313_),
    .y(_0603_)
  );
  al_nand3 _1293_ (
    .a(_0111_),
    .b(_0207_),
    .c(_0218_),
    .y(_0604_)
  );
  al_ao21ttf _1294_ (
    .a(_0240_),
    .b(_0310_),
    .c(_0256_),
    .y(_0605_)
  );
  al_nand3ftt _1295_ (
    .a(_0307_),
    .b(_0604_),
    .c(_0605_),
    .y(_0606_)
  );
  al_ao21ttf _1296_ (
    .a(_0604_),
    .b(_0605_),
    .c(_0307_),
    .y(_0607_)
  );
  al_nand3 _1297_ (
    .a(_0313_),
    .b(_0606_),
    .c(_0607_),
    .y(_0608_)
  );
  al_oa21ftt _1298_ (
    .a(N13),
    .b(N20),
    .c(N1),
    .y(_0609_)
  );
  al_ao21 _1299_ (
    .a(_0603_),
    .b(_0608_),
    .c(_0609_),
    .y(_0610_)
  );
  al_ao21ttf _1300_ (
    .a(N58),
    .b(N68),
    .c(N77),
    .y(_0611_)
  );
  al_ao21 _1301_ (
    .a(N58),
    .b(N50),
    .c(N68),
    .y(_0612_)
  );
  al_and3ftt _1302_ (
    .a(N13),
    .b(N1),
    .c(_0612_),
    .y(_0613_)
  );
  al_ao21ftf _1303_ (
    .a(_0390_),
    .b(_0611_),
    .c(_0613_),
    .y(_0614_)
  );
  al_or3ftt _1304_ (
    .a(_0026_),
    .b(_0173_),
    .c(_0016_),
    .y(_0615_)
  );
  al_nand3 _1305_ (
    .a(_0614_),
    .b(_0615_),
    .c(_0610_),
    .y(N5002)
  );
  al_nand2 _1306_ (
    .a(_0493_),
    .b(_0497_),
    .y(N5047)
  );
  al_ao21ttf _1307_ (
    .a(_0384_),
    .b(_0260_),
    .c(_0413_),
    .y(N5121)
  );
  al_nand2ft _1308_ (
    .a(N343),
    .b(N213),
    .y(_0616_)
  );
  al_or3ftt _1309_ (
    .a(_0616_),
    .b(_0578_),
    .c(_0354_),
    .y(_0617_)
  );
  al_aoi21ftf _1310_ (
    .a(_0616_),
    .b(N350),
    .c(_0617_),
    .y(_0618_)
  );
  al_aoi21 _1311_ (
    .a(_0592_),
    .b(_0596_),
    .c(_0618_),
    .y(_0619_)
  );
  al_ao21ttf _1312_ (
    .a(_0598_),
    .b(_0599_),
    .c(_0618_),
    .y(_0620_)
  );
  al_nand2ft _1313_ (
    .a(_0619_),
    .b(_0620_),
    .y(N5360)
  );
  assign N1279 = N13;
  assign N1334 = N1;
  assign N1345 = N20;
  assign N1346 = N20;
  assign N1347 = N20;
  assign N1348 = N20;
  assign N1349 = N20;
  assign N1350 = N20;
  assign N1351 = N20;
  assign N1352 = N20;
  assign N1369 = N33;
  assign N1493 = N68;
  assign N1496 = N68;
  assign N1499 = N107;
  assign N1502 = N107;
  assign N1726 = N50;
  assign N1735 = N1947;
  assign N1736 = N45;
  assign N1737 = N45;
  assign N1849 = N33;
  assign N1851 = N33;
  assign N1853 = N33;
  assign N1855 = N33;
  assign N1857 = N33;
  assign N1859 = N33;
  assign N1861 = N33;
  assign N1863 = N33;
  assign N1939 = N58;
  assign N1941 = N68;
  assign N1942 = N77;
  assign N1943 = N87;
  assign N1944 = N97;
  assign N1945 = N107;
  assign N1946 = N116;
  assign N655 = N50;
  assign N670 = N58;
  assign N683 = N68;
  assign N690 = N68;
  assign N699 = N77;
  assign N706 = N77;
  assign N715 = N87;
  assign N727 = N97;
  assign N740 = N107;
  assign N753 = N116;
  assign N772 = N1;
  assign N782 = N13;
  assign N798 = N20;
  assign N821 = N33;
  assign N836 = N45;
  assign N845 = N58;
  assign N851 = N68;
  assign N858 = N87;
  assign N864 = N97;
  assign N874 = N1;
  assign N877 = N68;
  assign N880 = N107;
  assign N886 = N190;
  assign N917 = N179;
  assign N923 = N343;
  assign N926 = N226;
  assign N929 = N232;
  assign N932 = N238;
  assign N935 = N244;
  assign N938 = N250;
  assign N941 = N257;
  assign N944 = N264;
  assign N947 = N270;
  assign N950 = N50;
  assign N953 = N58;
  assign N956 = N58;
  assign N959 = N97;
  assign N962 = N97;
  assign N965 = N330;
endmodule
