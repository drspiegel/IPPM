
module c2670(N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N32, N33, N34, N35, N36, N37, N40, N43, N44, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N138, N139, N140, N141, N142, N219, N224, N227, N230, N231, N234, N237, N241, N246, N253, N256, N259, N262, N263, N266, N269, N272, N275, N278, N281, N284, N287, N290, N294, N297, N301, N305, N309, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N143_I, N144_I, N145_I, N146_I, N147_I, N148_I, N149_I, N150_I, N151_I, N152_I, N153_I, N154_I, N155_I, N156_I, N157_I, N158_I, N159_I, N160_I, N161_I, N162_I, N163_I, N164_I, N165_I, N166_I, N167_I, N168_I, N169_I, N170_I, N171_I, N172_I, N173_I, N174_I, N175_I, N176_I, N177_I, N178_I, N179_I, N180_I, N181_I, N182_I, N183_I, N184_I, N185_I, N186_I, N187_I, N188_I, N189_I, N190_I, N191_I, N192_I, N193_I, N194_I, N195_I, N196_I, N197_I, N198_I, N199_I, N200_I, N201_I, N202_I, N203_I, N204_I, N205_I, N206_I, N207_I, N208_I, N209_I, N210_I, N211_I, N212_I, N213_I, N214_I, N215_I, N216_I, N217_I, N218_I, N398, N400, N401, N419, N420, N456, N457, N458, N487, N488, N489, N490, N491, N492, N493, N494, N792, N799, N805, N1026, N1028, N1029, N1269, N1277, N1448, N1726, N1816, N1817, N1818, N1819, N1820, N1821, N1969, N1970, N1971, N2010, N2012, N2014, N2016, N2018, N2020, N2022, N2387, N2388, N2389, N2390, N2496, N2643, N2644, N2891, N2925, N2970, N2971, N3038, N3079, N3546, N3671, N3803, N3804, N3809, N3851, N3875, N3881, N3882, N143_O, N144_O, N145_O, N146_O, N147_O, N148_O, N149_O, N150_O, N151_O, N152_O, N153_O, N154_O, N155_O, N156_O, N157_O, N158_O, N159_O, N160_O, N161_O, N162_O, N163_O, N164_O, N165_O, N166_O, N167_O, N168_O, N169_O, N170_O, N171_O, N172_O, N173_O, N174_O, N175_O, N176_O, N177_O, N178_O, N179_O, N180_O, N181_O, N182_O, N183_O, N184_O, N185_O, N186_O, N187_O, N188_O, N189_O, N190_O, N191_O, N192_O, N193_O, N194_O, N195_O, N196_O, N197_O, N198_O, N199_O, N200_O, N201_O, N202_O, N203_O, N204_O, N205_O, N206_O, N207_O, N208_O, N209_O, N210_O, N211_O, N212_O, N213_O, N214_O, N215_O, N216_O, N217_O, N218_O);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  wire _332_;
  wire _333_;
  wire _334_;
  wire _335_;
  wire _336_;
  wire _337_;
  wire _338_;
  wire _339_;
  input N1;
  input N100;
  input N101;
  input N102;
  output N1026;
  output N1028;
  output N1029;
  input N103;
  wire N1034;
  wire N1037;
  input N104;
  input N105;
  input N106;
  input N107;
  wire N1070;
  input N108;
  input N11;
  input N111;
  input N112;
  input N113;
  input N114;
  input N115;
  input N116;
  input N117;
  input N118;
  input N119;
  wire N1190;
  wire N1195;
  input N120;
  input N123;
  input N124;
  input N125;
  input N126;
  output N1269;
  input N127;
  output N1277;
  input N128;
  input N129;
  input N130;
  input N131;
  input N132;
  input N135;
  input N136;
  input N137;
  input N138;
  input N139;
  input N14;
  input N140;
  input N141;
  input N142;
  input N143_I;
  output N143_O;
  output N1448;
  input N144_I;
  output N144_O;
  input N145_I;
  output N145_O;
  input N146_I;
  output N146_O;
  input N147_I;
  output N147_O;
  input N148_I;
  output N148_O;
  input N149_I;
  output N149_O;
  input N15;
  input N150_I;
  output N150_O;
  wire N1519;
  input N151_I;
  output N151_O;
  wire N1520;
  wire N1521;
  wire N1522;
  wire N1523;
  wire N1524;
  wire N1525;
  wire N1526;
  wire N1527;
  wire N1528;
  input N152_I;
  output N152_O;
  input N153_I;
  output N153_O;
  input N154_I;
  output N154_O;
  input N155_I;
  output N155_O;
  input N156_I;
  output N156_O;
  wire N1572;
  wire N1573;
  wire N1574;
  wire N1575;
  wire N1576;
  wire N1577;
  input N157_I;
  output N157_O;
  input N158_I;
  output N158_O;
  wire N1591;
  input N159_I;
  output N159_O;
  input N16;
  input N160_I;
  output N160_O;
  wire N1612;
  wire N1615;
  wire N1619;
  input N161_I;
  output N161_O;
  wire N1624;
  wire N1628;
  input N162_I;
  output N162_O;
  wire N1631;
  wire N1634;
  input N163_I;
  output N163_O;
  input N164_I;
  output N164_O;
  input N165_I;
  output N165_O;
  input N166_I;
  output N166_O;
  input N167_I;
  output N167_O;
  input N168_I;
  output N168_O;
  input N169_I;
  output N169_O;
  input N170_I;
  output N170_O;
  input N171_I;
  output N171_O;
  output N1726;
  input N172_I;
  output N172_O;
  input N173_I;
  output N173_O;
  input N174_I;
  output N174_O;
  input N175_I;
  output N175_O;
  input N176_I;
  output N176_O;
  input N177_I;
  output N177_O;
  input N178_I;
  output N178_O;
  input N179_I;
  output N179_O;
  input N180_I;
  output N180_O;
  output N1816;
  output N1817;
  output N1818;
  output N1819;
  input N181_I;
  output N181_O;
  output N1820;
  output N1821;
  input N182_I;
  output N182_O;
  input N183_I;
  output N183_O;
  wire N1848;
  input N184_I;
  output N184_O;
  wire N1852;
  wire N1856;
  input N185_I;
  output N185_O;
  wire N1863;
  input N186_I;
  output N186_O;
  wire N1870;
  wire N1875;
  input N187_I;
  output N187_O;
  wire N1880;
  input N188_I;
  output N188_O;
  wire N1897;
  input N189_I;
  output N189_O;
  input N19;
  input N190_I;
  output N190_O;
  input N191_I;
  output N191_O;
  input N192_I;
  output N192_O;
  input N193_I;
  output N193_O;
  input N194_I;
  output N194_O;
  input N195_I;
  output N195_O;
  output N1969;
  input N196_I;
  output N196_O;
  output N1970;
  output N1971;
  input N197_I;
  output N197_O;
  input N198_I;
  output N198_O;
  input N199_I;
  output N199_O;
  input N2;
  input N20;
  input N200_I;
  output N200_O;
  output N2010;
  output N2012;
  output N2014;
  output N2016;
  output N2018;
  input N201_I;
  output N201_O;
  output N2020;
  output N2022;
  input N202_I;
  output N202_O;
  input N203_I;
  output N203_O;
  input N204_I;
  output N204_O;
  input N205_I;
  output N205_O;
  input N206_I;
  output N206_O;
  input N207_I;
  output N207_O;
  input N208_I;
  output N208_O;
  input N209_I;
  output N209_O;
  input N21;
  input N210_I;
  output N210_O;
  input N211_I;
  output N211_O;
  input N212_I;
  output N212_O;
  wire N2135;
  input N213_I;
  output N213_O;
  wire N2141;
  input N214_I;
  output N214_O;
  input N215_I;
  output N215_O;
  input N216_I;
  output N216_O;
  wire N2175;
  input N217_I;
  output N217_O;
  input N218_I;
  output N218_O;
  input N219;
  wire N2194;
  input N22;
  wire N2234;
  wire N2235;
  input N224;
  wire N2266;
  wire N2269;
  input N227;
  input N23;
  input N230;
  input N231;
  input N234;
  wire N2367;
  input N237;
  output N2387;
  output N2388;
  output N2389;
  output N2390;
  input N24;
  input N241;
  wire N2437;
  wire N2443;
  input N246;
  wire N2460;
  wire N2475;
  wire N2481;
  output N2496;
  input N25;
  wire N2521;
  input N253;
  input N256;
  input N259;
  input N26;
  wire N2617;
  input N262;
  wire N2620;
  wire N2628;
  input N263;
  wire N2630;
  output N2643;
  output N2644;
  wire N2645;
  wire N2655;
  wire N2656;
  input N266;
  input N269;
  wire N2695;
  wire N2696;
  wire N2697;
  wire N2698;
  wire N2699;
  input N27;
  wire N2700;
  wire N2701;
  wire N2702;
  input N272;
  input N275;
  input N278;
  input N28;
  input N281;
  wire N2817;
  input N284;
  input N287;
  output N2891;
  input N29;
  input N290;
  output N2925;
  wire N2931;
  input N294;
  input N297;
  output N2970;
  output N2971;
  input N3;
  input N301;
  output N3038;
  input N305;
  output N3079;
  input N309;
  input N313;
  input N316;
  input N319;
  input N32;
  input N322;
  input N325;
  input N328;
  input N33;
  input N331;
  input N334;
  input N337;
  input N34;
  input N340;
  input N343;
  input N346;
  input N349;
  input N35;
  input N352;
  output N3546;
  input N355;
  input N36;
  wire N3600;
  output N3671;
  input N37;
  wire N3780;
  wire N3790;
  output N3803;
  output N3804;
  output N3809;
  wire N3840;
  wire N3843;
  output N3851;
  output N3875;
  wire N3877;
  output N3881;
  output N3882;
  output N398;
  input N4;
  input N40;
  output N400;
  output N401;
  output N419;
  output N420;
  input N43;
  input N44;
  output N456;
  output N457;
  output N458;
  input N47;
  input N48;
  output N487;
  output N488;
  output N489;
  input N49;
  output N490;
  output N491;
  output N492;
  output N493;
  output N494;
  wire N496;
  input N5;
  input N50;
  wire N500;
  wire N503;
  wire N506;
  wire N509;
  input N51;
  input N52;
  wire N521;
  input N53;
  input N54;
  input N55;
  wire N550;
  input N56;
  wire N562;
  input N57;
  wire N582;
  wire N594;
  input N6;
  input N60;
  input N61;
  wire N613;
  input N62;
  wire N625;
  input N63;
  wire N637;
  input N64;
  wire N643;
  input N65;
  input N66;
  input N67;
  input N68;
  input N69;
  wire N693;
  wire N699;
  input N7;
  input N72;
  input N73;
  wire N735;
  wire N738;
  input N74;
  wire N741;
  wire N744;
  wire N747;
  input N75;
  wire N750;
  wire N753;
  wire N756;
  wire N759;
  input N76;
  wire N762;
  wire N765;
  wire N768;
  input N77;
  wire N771;
  wire N774;
  wire N777;
  input N78;
  wire N780;
  wire N783;
  wire N786;
  input N79;
  output N792;
  output N799;
  input N8;
  input N80;
  output N805;
  input N81;
  input N82;
  input N85;
  input N86;
  input N87;
  input N88;
  input N89;
  input N90;
  input N91;
  input N92;
  input N93;
  input N94;
  input N95;
  input N96;
  input N99;
  al_inv _340_ (
    .a(N44),
    .y(N487)
  );
  al_inv _341_ (
    .a(N132),
    .y(N488)
  );
  al_inv _342_ (
    .a(N82),
    .y(N489)
  );
  al_inv _343_ (
    .a(N96),
    .y(N490)
  );
  al_inv _344_ (
    .a(N69),
    .y(N491)
  );
  al_inv _345_ (
    .a(N120),
    .y(N492)
  );
  al_inv _346_ (
    .a(N57),
    .y(N493)
  );
  al_inv _347_ (
    .a(N108),
    .y(N494)
  );
  al_and2 _348_ (
    .a(N309),
    .b(N305),
    .y(_000_)
  );
  al_nand3 _349_ (
    .a(N301),
    .b(N297),
    .c(_000_),
    .y(N792)
  );
  al_nand3 _350_ (
    .a(N2),
    .b(N15),
    .c(N237),
    .y(N799)
  );
  al_nand2 _351_ (
    .a(N237),
    .b(N7),
    .y(N1028)
  );
  al_nand3 _352_ (
    .a(N237),
    .b(N7),
    .c(N231),
    .y(N1029)
  );
  al_nand3 _353_ (
    .a(N237),
    .b(N7),
    .c(N325),
    .y(N1269)
  );
  al_and2 _354_ (
    .a(N69),
    .b(N120),
    .y(_001_)
  );
  al_and3 _355_ (
    .a(N57),
    .b(N108),
    .c(_001_),
    .y(_002_)
  );
  al_and2 _356_ (
    .a(N132),
    .b(N82),
    .y(_003_)
  );
  al_nand3 _357_ (
    .a(N44),
    .b(N96),
    .c(_003_),
    .y(_004_)
  );
  al_and2ft _358_ (
    .a(_004_),
    .b(_002_),
    .y(N1277)
  );
  al_inv _359_ (
    .a(N1277),
    .y(N1448)
  );
  al_nand2 _360_ (
    .a(N325),
    .b(_004_),
    .y(_005_)
  );
  al_aoi21ftf _361_ (
    .a(_002_),
    .b(N231),
    .c(_005_),
    .y(N1726)
  );
  al_and3 _362_ (
    .a(N237),
    .b(N224),
    .c(N1726),
    .y(_006_)
  );
  al_nand2 _363_ (
    .a(N36),
    .b(_006_),
    .y(N1970)
  );
  al_ao21ttf _364_ (
    .a(N1),
    .b(N3),
    .c(_006_),
    .y(N1971)
  );
  al_mux2l _365_ (
    .a(N53),
    .b(N91),
    .s(N227),
    .y(_007_)
  );
  al_and2ft _366_ (
    .a(N227),
    .b(N234),
    .y(_008_)
  );
  al_and3 _367_ (
    .a(N227),
    .b(N234),
    .c(N78),
    .y(_009_)
  );
  al_aoi21 _368_ (
    .a(N65),
    .b(_008_),
    .c(_009_),
    .y(_010_)
  );
  al_ao21ftf _369_ (
    .a(N234),
    .b(_007_),
    .c(_010_),
    .y(N2010)
  );
  al_mux2l _370_ (
    .a(N52),
    .b(N90),
    .s(N227),
    .y(_011_)
  );
  al_and3 _371_ (
    .a(N227),
    .b(N234),
    .c(N77),
    .y(_012_)
  );
  al_aoi21 _372_ (
    .a(N64),
    .b(_008_),
    .c(_012_),
    .y(_013_)
  );
  al_aoi21ftf _373_ (
    .a(N234),
    .b(_011_),
    .c(_013_),
    .y(N1821)
  );
  al_inv _374_ (
    .a(N1821),
    .y(N2012)
  );
  al_mux2l _375_ (
    .a(N50),
    .b(N88),
    .s(N227),
    .y(_014_)
  );
  al_and3 _376_ (
    .a(N227),
    .b(N234),
    .c(N75),
    .y(_015_)
  );
  al_aoi21 _377_ (
    .a(N62),
    .b(_008_),
    .c(_015_),
    .y(_016_)
  );
  al_aoi21ftf _378_ (
    .a(N234),
    .b(_014_),
    .c(_016_),
    .y(N1819)
  );
  al_inv _379_ (
    .a(N1819),
    .y(N2016)
  );
  al_and3ftt _380_ (
    .a(N74),
    .b(N227),
    .c(N234),
    .y(_017_)
  );
  al_mux2l _381_ (
    .a(N49),
    .b(N87),
    .s(N227),
    .y(_018_)
  );
  al_oai21ttf _382_ (
    .a(N234),
    .b(_018_),
    .c(_017_),
    .y(_019_)
  );
  al_inv _383_ (
    .a(_019_),
    .y(N2018)
  );
  al_mux2l _384_ (
    .a(N48),
    .b(N86),
    .s(N227),
    .y(_020_)
  );
  al_and3 _385_ (
    .a(N227),
    .b(N234),
    .c(N73),
    .y(_021_)
  );
  al_aoi21 _386_ (
    .a(N61),
    .b(_008_),
    .c(_021_),
    .y(_022_)
  );
  al_ao21ftf _387_ (
    .a(N234),
    .b(_020_),
    .c(_022_),
    .y(N2020)
  );
  al_mux2l _388_ (
    .a(N47),
    .b(N85),
    .s(N227),
    .y(_023_)
  );
  al_and3 _389_ (
    .a(N227),
    .b(N234),
    .c(N72),
    .y(_024_)
  );
  al_aoi21 _390_ (
    .a(N60),
    .b(_008_),
    .c(_024_),
    .y(_025_)
  );
  al_ao21ftf _391_ (
    .a(N234),
    .b(_023_),
    .c(_025_),
    .y(N2022)
  );
  al_nand3fft _392_ (
    .a(N319),
    .b(N322),
    .c(N138),
    .y(_026_)
  );
  al_nand3 _393_ (
    .a(N319),
    .b(N322),
    .c(N114),
    .y(_027_)
  );
  al_and3ftt _394_ (
    .a(N322),
    .b(N319),
    .c(N102),
    .y(_028_)
  );
  al_and2ft _395_ (
    .a(N319),
    .b(N322),
    .y(_029_)
  );
  al_aoi21 _396_ (
    .a(N126),
    .b(_029_),
    .c(_028_),
    .y(_030_)
  );
  al_nand3 _397_ (
    .a(_026_),
    .b(_027_),
    .c(_030_),
    .y(_031_)
  );
  al_inv _398_ (
    .a(_031_),
    .y(N1818)
  );
  al_mux2l _399_ (
    .a(N51),
    .b(N89),
    .s(N227),
    .y(_032_)
  );
  al_and3 _400_ (
    .a(N227),
    .b(N234),
    .c(N76),
    .y(_033_)
  );
  al_aoi21 _401_ (
    .a(N63),
    .b(_008_),
    .c(_033_),
    .y(_034_)
  );
  al_aoi21ftf _402_ (
    .a(N234),
    .b(_032_),
    .c(_034_),
    .y(N1820)
  );
  al_inv _403_ (
    .a(N1820),
    .y(N2014)
  );
  al_inv _404_ (
    .a(N124),
    .y(_035_)
  );
  al_nor2 _405_ (
    .a(N319),
    .b(N322),
    .y(_036_)
  );
  al_and2ft _406_ (
    .a(N322),
    .b(N319),
    .y(_037_)
  );
  al_and3 _407_ (
    .a(N319),
    .b(N322),
    .c(N112),
    .y(_038_)
  );
  al_aoi21 _408_ (
    .a(N100),
    .b(_037_),
    .c(_038_),
    .y(_039_)
  );
  al_ao21ttf _409_ (
    .a(N136),
    .b(_036_),
    .c(_039_),
    .y(_040_)
  );
  al_aoi21ftt _410_ (
    .a(_035_),
    .b(_029_),
    .c(_040_),
    .y(N1817)
  );
  al_and3fft _411_ (
    .a(N319),
    .b(N322),
    .c(N137),
    .y(_041_)
  );
  al_nand3ftt _412_ (
    .a(N322),
    .b(N319),
    .c(N101),
    .y(_042_)
  );
  al_nand3 _413_ (
    .a(N319),
    .b(N322),
    .c(N113),
    .y(_043_)
  );
  al_and3ftt _414_ (
    .a(N319),
    .b(N322),
    .c(N125),
    .y(_044_)
  );
  al_and3ftt _415_ (
    .a(_044_),
    .b(_042_),
    .c(_043_),
    .y(_045_)
  );
  al_and2ft _416_ (
    .a(_041_),
    .b(_045_),
    .y(N1816)
  );
  al_and2ft _417_ (
    .a(N263),
    .b(N352),
    .y(_046_)
  );
  al_nand2ft _418_ (
    .a(N352),
    .b(N263),
    .y(_047_)
  );
  al_nor2 _419_ (
    .a(N275),
    .b(N272),
    .y(_048_)
  );
  al_nand2 _420_ (
    .a(N275),
    .b(N272),
    .y(_049_)
  );
  al_nand2ft _421_ (
    .a(_048_),
    .b(_049_),
    .y(_050_)
  );
  al_and3ftt _422_ (
    .a(_046_),
    .b(_047_),
    .c(_050_),
    .y(_051_)
  );
  al_ao21ftt _423_ (
    .a(_046_),
    .b(_047_),
    .c(_050_),
    .y(_052_)
  );
  al_nand2ft _424_ (
    .a(_051_),
    .b(_052_),
    .y(_053_)
  );
  al_and2ft _425_ (
    .a(N266),
    .b(N269),
    .y(_054_)
  );
  al_nand2ft _426_ (
    .a(N269),
    .b(N266),
    .y(_055_)
  );
  al_nand2ft _427_ (
    .a(_054_),
    .b(_055_),
    .y(_056_)
  );
  al_and2ft _428_ (
    .a(N287),
    .b(N284),
    .y(_057_)
  );
  al_nand2ft _429_ (
    .a(N284),
    .b(N287),
    .y(_058_)
  );
  al_and3ftt _430_ (
    .a(_057_),
    .b(_058_),
    .c(_056_),
    .y(_059_)
  );
  al_ao21ftt _431_ (
    .a(_057_),
    .b(_058_),
    .c(_056_),
    .y(_060_)
  );
  al_nor2 _432_ (
    .a(N281),
    .b(N278),
    .y(_061_)
  );
  al_nand2 _433_ (
    .a(N281),
    .b(N278),
    .y(_062_)
  );
  al_nand2ft _434_ (
    .a(_061_),
    .b(_062_),
    .y(_063_)
  );
  al_nor3fft _435_ (
    .a(_063_),
    .b(_060_),
    .c(_059_),
    .y(_064_)
  );
  al_oai21ftf _436_ (
    .a(_060_),
    .b(_059_),
    .c(_063_),
    .y(_065_)
  );
  al_nand3fft _437_ (
    .a(_064_),
    .b(_053_),
    .c(_065_),
    .y(_066_)
  );
  al_aoi21ftf _438_ (
    .a(_064_),
    .b(_065_),
    .c(_053_),
    .y(_067_)
  );
  al_nor2ft _439_ (
    .a(_066_),
    .b(_067_),
    .y(_068_)
  );
  al_inv _440_ (
    .a(_068_),
    .y(N2971)
  );
  al_nand2 _441_ (
    .a(N301),
    .b(N297),
    .y(_069_)
  );
  al_nor2 _442_ (
    .a(N301),
    .b(N297),
    .y(_070_)
  );
  al_nand2ft _443_ (
    .a(_070_),
    .b(_069_),
    .y(_071_)
  );
  al_or2 _444_ (
    .a(N316),
    .b(N313),
    .y(_072_)
  );
  al_nand2 _445_ (
    .a(N316),
    .b(N313),
    .y(_073_)
  );
  al_and3 _446_ (
    .a(_072_),
    .b(_073_),
    .c(_071_),
    .y(_074_)
  );
  al_aoi21 _447_ (
    .a(_072_),
    .b(_073_),
    .c(_071_),
    .y(_075_)
  );
  al_or2 _448_ (
    .a(_074_),
    .b(_075_),
    .y(_076_)
  );
  al_nor2 _449_ (
    .a(N309),
    .b(N305),
    .y(_077_)
  );
  al_nand2ft _450_ (
    .a(N294),
    .b(N355),
    .y(_078_)
  );
  al_and2ft _451_ (
    .a(N355),
    .b(N294),
    .y(_079_)
  );
  al_and2ft _452_ (
    .a(_079_),
    .b(_078_),
    .y(_080_)
  );
  al_nand3fft _453_ (
    .a(_000_),
    .b(_077_),
    .c(_080_),
    .y(_081_)
  );
  al_oai21ttf _454_ (
    .a(_000_),
    .b(_077_),
    .c(_080_),
    .y(_082_)
  );
  al_or3fft _455_ (
    .a(_081_),
    .b(_082_),
    .c(_076_),
    .y(_083_)
  );
  al_aoi21ttf _456_ (
    .a(_081_),
    .b(_082_),
    .c(_076_),
    .y(_084_)
  );
  al_nand2ft _457_ (
    .a(_084_),
    .b(_083_),
    .y(N2970)
  );
  al_and3 _458_ (
    .a(N319),
    .b(N322),
    .c(N111),
    .y(_085_)
  );
  al_aoi21 _459_ (
    .a(N99),
    .b(_037_),
    .c(_085_),
    .y(_086_)
  );
  al_aoi21ttf _460_ (
    .a(N123),
    .b(_029_),
    .c(_086_),
    .y(_087_)
  );
  al_ao21ttf _461_ (
    .a(N135),
    .b(_036_),
    .c(_087_),
    .y(_088_)
  );
  al_oa21ttf _462_ (
    .a(N313),
    .b(_088_),
    .c(N316),
    .y(_089_)
  );
  al_ao21ttf _463_ (
    .a(N313),
    .b(_088_),
    .c(_089_),
    .y(N2891)
  );
  al_and2ft _464_ (
    .a(N259),
    .b(N256),
    .y(_090_)
  );
  al_nand2ft _465_ (
    .a(N256),
    .b(N259),
    .y(_091_)
  );
  al_and2ft _466_ (
    .a(N349),
    .b(N346),
    .y(_092_)
  );
  al_nand2ft _467_ (
    .a(N346),
    .b(N349),
    .y(_093_)
  );
  al_nand2ft _468_ (
    .a(_092_),
    .b(_093_),
    .y(_094_)
  );
  al_and3ftt _469_ (
    .a(_090_),
    .b(_091_),
    .c(_094_),
    .y(_095_)
  );
  al_ao21ftt _470_ (
    .a(_090_),
    .b(_091_),
    .c(_094_),
    .y(_096_)
  );
  al_nand2ft _471_ (
    .a(_095_),
    .b(_096_),
    .y(_097_)
  );
  al_and2ft _472_ (
    .a(N340),
    .b(N343),
    .y(_098_)
  );
  al_nand2ft _473_ (
    .a(N343),
    .b(N340),
    .y(_099_)
  );
  al_and2ft _474_ (
    .a(N337),
    .b(N334),
    .y(_100_)
  );
  al_nand2ft _475_ (
    .a(N334),
    .b(N337),
    .y(_101_)
  );
  al_nand2ft _476_ (
    .a(_100_),
    .b(_101_),
    .y(_102_)
  );
  al_nand3ftt _477_ (
    .a(_098_),
    .b(_099_),
    .c(_102_),
    .y(_103_)
  );
  al_ao21ftt _478_ (
    .a(_098_),
    .b(_099_),
    .c(_102_),
    .y(_104_)
  );
  al_nor2 _479_ (
    .a(N328),
    .b(N331),
    .y(_105_)
  );
  al_nand2 _480_ (
    .a(N328),
    .b(N331),
    .y(_106_)
  );
  al_nand2ft _481_ (
    .a(_105_),
    .b(_106_),
    .y(_107_)
  );
  al_nand3ftt _482_ (
    .a(_107_),
    .b(_103_),
    .c(_104_),
    .y(_108_)
  );
  al_ao21ttf _483_ (
    .a(_103_),
    .b(_104_),
    .c(_107_),
    .y(_109_)
  );
  al_nand3 _484_ (
    .a(_108_),
    .b(_097_),
    .c(_109_),
    .y(_110_)
  );
  al_ao21 _485_ (
    .a(_108_),
    .b(_109_),
    .c(_097_),
    .y(_111_)
  );
  al_nand3 _486_ (
    .a(N14),
    .b(_111_),
    .c(_110_),
    .y(_112_)
  );
  al_inv _487_ (
    .a(_112_),
    .y(N2925)
  );
  al_mux2l _488_ (
    .a(N54),
    .b(N92),
    .s(N227),
    .y(_113_)
  );
  al_and3 _489_ (
    .a(N227),
    .b(N234),
    .c(N79),
    .y(_114_)
  );
  al_aoi21 _490_ (
    .a(N66),
    .b(_008_),
    .c(_114_),
    .y(_115_)
  );
  al_aoi21ftf _491_ (
    .a(N234),
    .b(_113_),
    .c(_115_),
    .y(_116_)
  );
  al_inv _492_ (
    .a(_116_),
    .y(_117_)
  );
  al_mux2h _493_ (
    .a(N4),
    .b(_117_),
    .s(N16),
    .y(_118_)
  );
  al_nand2 _494_ (
    .a(N259),
    .b(_118_),
    .y(_119_)
  );
  al_inv _495_ (
    .a(N272),
    .y(_120_)
  );
  al_inv _496_ (
    .a(N22),
    .y(_121_)
  );
  al_mux2h _497_ (
    .a(_121_),
    .b(N1819),
    .s(N16),
    .y(_122_)
  );
  al_or2 _498_ (
    .a(_120_),
    .b(_122_),
    .y(_123_)
  );
  al_inv _499_ (
    .a(N301),
    .y(_124_)
  );
  al_nand3ftt _500_ (
    .a(N319),
    .b(N322),
    .c(N126),
    .y(_125_)
  );
  al_and3ftt _501_ (
    .a(_028_),
    .b(_027_),
    .c(_125_),
    .y(_126_)
  );
  al_nand3 _502_ (
    .a(N29),
    .b(_026_),
    .c(_126_),
    .y(_127_)
  );
  al_oai21 _503_ (
    .a(N29),
    .b(N27),
    .c(_127_),
    .y(_128_)
  );
  al_or2 _504_ (
    .a(_124_),
    .b(_128_),
    .y(_129_)
  );
  al_nand3 _505_ (
    .a(_123_),
    .b(_129_),
    .c(_119_),
    .y(_130_)
  );
  al_inv _506_ (
    .a(N275),
    .y(_131_)
  );
  al_inv _507_ (
    .a(N23),
    .y(_132_)
  );
  al_mux2h _508_ (
    .a(_132_),
    .b(_019_),
    .s(N16),
    .y(_133_)
  );
  al_and2 _509_ (
    .a(_131_),
    .b(_133_),
    .y(_134_)
  );
  al_inv _510_ (
    .a(N5),
    .y(_135_)
  );
  al_mux2h _511_ (
    .a(_135_),
    .b(N1821),
    .s(N16),
    .y(_136_)
  );
  al_oai21ftf _512_ (
    .a(N266),
    .b(_136_),
    .c(_134_),
    .y(_137_)
  );
  al_mux2h _513_ (
    .a(N6),
    .b(N2020),
    .s(N16),
    .y(_138_)
  );
  al_nor2 _514_ (
    .a(N278),
    .b(_138_),
    .y(_139_)
  );
  al_inv _515_ (
    .a(N284),
    .y(_140_)
  );
  al_inv _516_ (
    .a(N25),
    .y(_141_)
  );
  al_inv _517_ (
    .a(N131),
    .y(_142_)
  );
  al_and2 _518_ (
    .a(N319),
    .b(N322),
    .y(_143_)
  );
  al_and3ftt _519_ (
    .a(N319),
    .b(N322),
    .c(N119),
    .y(_144_)
  );
  al_aoi21 _520_ (
    .a(N95),
    .b(_037_),
    .c(_144_),
    .y(_145_)
  );
  al_aoi21ttf _521_ (
    .a(N107),
    .b(_143_),
    .c(_145_),
    .y(_146_)
  );
  al_aoi21ftf _522_ (
    .a(_142_),
    .b(_036_),
    .c(_146_),
    .y(_147_)
  );
  al_mux2h _523_ (
    .a(_141_),
    .b(_147_),
    .s(N29),
    .y(_148_)
  );
  al_or2 _524_ (
    .a(_140_),
    .b(_148_),
    .y(_149_)
  );
  al_nand3fft _525_ (
    .a(_137_),
    .b(_139_),
    .c(_149_),
    .y(_150_)
  );
  al_nand2ft _526_ (
    .a(N266),
    .b(_136_),
    .y(_151_)
  );
  al_and2 _527_ (
    .a(N278),
    .b(_138_),
    .y(_152_)
  );
  al_inv _528_ (
    .a(N19),
    .y(_153_)
  );
  al_mux2l _529_ (
    .a(N43),
    .b(N81),
    .s(N227),
    .y(_154_)
  );
  al_and3 _530_ (
    .a(N227),
    .b(N234),
    .c(N68),
    .y(_155_)
  );
  al_aoi21 _531_ (
    .a(N56),
    .b(_008_),
    .c(_155_),
    .y(_156_)
  );
  al_aoi21ftf _532_ (
    .a(N234),
    .b(_154_),
    .c(_156_),
    .y(_157_)
  );
  al_mux2h _533_ (
    .a(_153_),
    .b(_157_),
    .s(N16),
    .y(_158_)
  );
  al_nor2 _534_ (
    .a(_131_),
    .b(_133_),
    .y(_159_)
  );
  al_oa21ftf _535_ (
    .a(N256),
    .b(_158_),
    .c(_159_),
    .y(_160_)
  );
  al_and3ftt _536_ (
    .a(_152_),
    .b(_151_),
    .c(_160_),
    .y(_161_)
  );
  al_nor3ftt _537_ (
    .a(_161_),
    .b(_150_),
    .c(_130_),
    .y(_162_)
  );
  al_and3ftt _538_ (
    .a(N319),
    .b(N322),
    .c(N127),
    .y(_163_)
  );
  al_and3fft _539_ (
    .a(N319),
    .b(N322),
    .c(N139),
    .y(_164_)
  );
  al_and3 _540_ (
    .a(N319),
    .b(N322),
    .c(N115),
    .y(_165_)
  );
  al_aoi21 _541_ (
    .a(N103),
    .b(_037_),
    .c(_165_),
    .y(_166_)
  );
  al_nand3fft _542_ (
    .a(_163_),
    .b(_164_),
    .c(_166_),
    .y(_167_)
  );
  al_mux2h _543_ (
    .a(N33),
    .b(_167_),
    .s(N29),
    .y(_168_)
  );
  al_or2 _544_ (
    .a(N297),
    .b(_168_),
    .y(_169_)
  );
  al_and2 _545_ (
    .a(N297),
    .b(_168_),
    .y(_170_)
  );
  al_inv _546_ (
    .a(N294),
    .y(_171_)
  );
  al_and3 _547_ (
    .a(N319),
    .b(N322),
    .c(N116),
    .y(_172_)
  );
  al_aoi21 _548_ (
    .a(N104),
    .b(_037_),
    .c(_172_),
    .y(_173_)
  );
  al_aoi21ttf _549_ (
    .a(N128),
    .b(_029_),
    .c(_173_),
    .y(_174_)
  );
  al_ao21ttf _550_ (
    .a(N140),
    .b(_036_),
    .c(_174_),
    .y(_175_)
  );
  al_mux2h _551_ (
    .a(N26),
    .b(_175_),
    .s(N29),
    .y(_176_)
  );
  al_and2 _552_ (
    .a(_171_),
    .b(_176_),
    .y(_177_)
  );
  al_or2 _553_ (
    .a(_171_),
    .b(_176_),
    .y(_178_)
  );
  al_inv _554_ (
    .a(N287),
    .y(_179_)
  );
  al_and3ftt _555_ (
    .a(N319),
    .b(N322),
    .c(N129),
    .y(_180_)
  );
  al_aoi21 _556_ (
    .a(N105),
    .b(_037_),
    .c(_180_),
    .y(_181_)
  );
  al_aoi21ttf _557_ (
    .a(N117),
    .b(_143_),
    .c(_181_),
    .y(_182_)
  );
  al_ao21ttf _558_ (
    .a(N141),
    .b(_036_),
    .c(_182_),
    .y(_183_)
  );
  al_mux2h _559_ (
    .a(N32),
    .b(_183_),
    .s(N29),
    .y(_184_)
  );
  al_and2 _560_ (
    .a(_179_),
    .b(_184_),
    .y(_185_)
  );
  al_or2 _561_ (
    .a(_179_),
    .b(_184_),
    .y(_186_)
  );
  al_nand2ft _562_ (
    .a(_185_),
    .b(_186_),
    .y(_187_)
  );
  al_aoi21ftf _563_ (
    .a(_177_),
    .b(_178_),
    .c(_187_),
    .y(_188_)
  );
  al_and3ftt _564_ (
    .a(_170_),
    .b(_169_),
    .c(_188_),
    .y(_189_)
  );
  al_mux2h _565_ (
    .a(N24),
    .b(N2022),
    .s(N16),
    .y(_190_)
  );
  al_or2 _566_ (
    .a(N281),
    .b(_190_),
    .y(_191_)
  );
  al_nand3ftt _567_ (
    .a(_041_),
    .b(N29),
    .c(_045_),
    .y(_192_)
  );
  al_oa21 _568_ (
    .a(N29),
    .b(N34),
    .c(_192_),
    .y(_193_)
  );
  al_oa21 _569_ (
    .a(N305),
    .b(_193_),
    .c(_191_),
    .y(_194_)
  );
  al_and2ft _570_ (
    .a(N16),
    .b(N20),
    .y(_195_)
  );
  al_aoi21 _571_ (
    .a(N16),
    .b(N2010),
    .c(_195_),
    .y(_196_)
  );
  al_and2 _572_ (
    .a(N263),
    .b(_196_),
    .y(_197_)
  );
  al_or2 _573_ (
    .a(N263),
    .b(_196_),
    .y(_198_)
  );
  al_aoi21ftf _574_ (
    .a(_197_),
    .b(_198_),
    .c(_194_),
    .y(_199_)
  );
  al_oai21 _575_ (
    .a(N29),
    .b(N28),
    .c(N11),
    .y(_200_)
  );
  al_oai21ftf _576_ (
    .a(N29),
    .b(_088_),
    .c(_200_),
    .y(_201_)
  );
  al_oa21ttf _577_ (
    .a(N259),
    .b(_118_),
    .c(_201_),
    .y(_202_)
  );
  al_nor2 _578_ (
    .a(N29),
    .b(N35),
    .y(_203_)
  );
  al_aoi21 _579_ (
    .a(N29),
    .b(N1817),
    .c(_203_),
    .y(_204_)
  );
  al_or2 _580_ (
    .a(N309),
    .b(_204_),
    .y(_205_)
  );
  al_nand2 _581_ (
    .a(N309),
    .b(_204_),
    .y(_206_)
  );
  al_and3 _582_ (
    .a(_205_),
    .b(_206_),
    .c(_202_),
    .y(_207_)
  );
  al_nand2 _583_ (
    .a(N281),
    .b(_190_),
    .y(_208_)
  );
  al_aoi21ftf _584_ (
    .a(N256),
    .b(_158_),
    .c(_208_),
    .y(_209_)
  );
  al_mux2h _585_ (
    .a(N21),
    .b(N2014),
    .s(N16),
    .y(_210_)
  );
  al_or2 _586_ (
    .a(N269),
    .b(_210_),
    .y(_211_)
  );
  al_nand2 _587_ (
    .a(N305),
    .b(_193_),
    .y(_212_)
  );
  al_nand3 _588_ (
    .a(_209_),
    .b(_212_),
    .c(_211_),
    .y(_213_)
  );
  al_nand2 _589_ (
    .a(N269),
    .b(_210_),
    .y(_214_)
  );
  al_aoi21ftf _590_ (
    .a(N284),
    .b(_148_),
    .c(_214_),
    .y(_215_)
  );
  al_nand2 _591_ (
    .a(_124_),
    .b(_128_),
    .y(_216_)
  );
  al_aoi21ftf _592_ (
    .a(N272),
    .b(_122_),
    .c(_216_),
    .y(_217_)
  );
  al_nor3fft _593_ (
    .a(_217_),
    .b(_215_),
    .c(_213_),
    .y(_218_)
  );
  al_and3 _594_ (
    .a(_199_),
    .b(_207_),
    .c(_218_),
    .y(_219_)
  );
  al_and3 _595_ (
    .a(_162_),
    .b(_189_),
    .c(_219_),
    .y(N3038)
  );
  al_inv _596_ (
    .a(N3038),
    .y(N3079)
  );
  al_inv _597_ (
    .a(N37),
    .y(_220_)
  );
  al_or2 _598_ (
    .a(N1816),
    .b(_088_),
    .y(_221_)
  );
  al_nand2 _599_ (
    .a(N1816),
    .b(_088_),
    .y(_222_)
  );
  al_and3 _600_ (
    .a(N1817),
    .b(_222_),
    .c(_221_),
    .y(_223_)
  );
  al_ao21 _601_ (
    .a(_222_),
    .b(_221_),
    .c(N1817),
    .y(_224_)
  );
  al_and2ft _602_ (
    .a(_223_),
    .b(_224_),
    .y(_225_)
  );
  al_and3ftt _603_ (
    .a(N322),
    .b(N319),
    .c(N106),
    .y(_226_)
  );
  al_and3 _604_ (
    .a(N319),
    .b(N322),
    .c(N118),
    .y(_227_)
  );
  al_and3fft _605_ (
    .a(N319),
    .b(N322),
    .c(N142),
    .y(_228_)
  );
  al_aoi21 _606_ (
    .a(N130),
    .b(_029_),
    .c(_228_),
    .y(_229_)
  );
  al_nand3fft _607_ (
    .a(_226_),
    .b(_227_),
    .c(_229_),
    .y(_230_)
  );
  al_and2ft _608_ (
    .a(_230_),
    .b(_167_),
    .y(_231_)
  );
  al_nand2ft _609_ (
    .a(_167_),
    .b(_230_),
    .y(_232_)
  );
  al_nand2ft _610_ (
    .a(_231_),
    .b(_232_),
    .y(_233_)
  );
  al_nand2ft _611_ (
    .a(_147_),
    .b(_183_),
    .y(_234_)
  );
  al_and2ft _612_ (
    .a(_183_),
    .b(_147_),
    .y(_235_)
  );
  al_oai21ftf _613_ (
    .a(_234_),
    .b(_235_),
    .c(_233_),
    .y(_236_)
  );
  al_nand3ftt _614_ (
    .a(_235_),
    .b(_234_),
    .c(_233_),
    .y(_237_)
  );
  al_and2ft _615_ (
    .a(_031_),
    .b(_175_),
    .y(_238_)
  );
  al_or2ft _616_ (
    .a(_031_),
    .b(_175_),
    .y(_239_)
  );
  al_nand2ft _617_ (
    .a(_238_),
    .b(_239_),
    .y(_240_)
  );
  al_ao21 _618_ (
    .a(_237_),
    .b(_236_),
    .c(_240_),
    .y(_241_)
  );
  al_nand3 _619_ (
    .a(_240_),
    .b(_237_),
    .c(_236_),
    .y(_242_)
  );
  al_ao21 _620_ (
    .a(_242_),
    .b(_241_),
    .c(_225_),
    .y(_243_)
  );
  al_nand3 _621_ (
    .a(_225_),
    .b(_242_),
    .c(_241_),
    .y(_244_)
  );
  al_and3 _622_ (
    .a(_220_),
    .b(_244_),
    .c(_243_),
    .y(N3671)
  );
  al_nand2ft _623_ (
    .a(N2020),
    .b(N2022),
    .y(_245_)
  );
  al_and2ft _624_ (
    .a(N2022),
    .b(N2020),
    .y(_246_)
  );
  al_or2 _625_ (
    .a(_019_),
    .b(N1819),
    .y(_247_)
  );
  al_and2 _626_ (
    .a(_019_),
    .b(N1819),
    .y(_248_)
  );
  al_nand2ft _627_ (
    .a(_248_),
    .b(_247_),
    .y(_249_)
  );
  al_aoi21ftf _628_ (
    .a(_246_),
    .b(_245_),
    .c(_249_),
    .y(_250_)
  );
  al_and3fft _629_ (
    .a(_246_),
    .b(_249_),
    .c(_245_),
    .y(_251_)
  );
  al_or2 _630_ (
    .a(_250_),
    .b(_251_),
    .y(_252_)
  );
  al_mux2l _631_ (
    .a(N55),
    .b(N93),
    .s(N227),
    .y(_253_)
  );
  al_and3 _632_ (
    .a(N227),
    .b(N234),
    .c(N80),
    .y(_254_)
  );
  al_aoi21 _633_ (
    .a(N67),
    .b(_008_),
    .c(_254_),
    .y(_255_)
  );
  al_ao21ftf _634_ (
    .a(N234),
    .b(_253_),
    .c(_255_),
    .y(_256_)
  );
  al_and2ft _635_ (
    .a(_256_),
    .b(_157_),
    .y(_257_)
  );
  al_nand2ft _636_ (
    .a(_157_),
    .b(_256_),
    .y(_258_)
  );
  al_nand2ft _637_ (
    .a(_257_),
    .b(_258_),
    .y(_259_)
  );
  al_and2ft _638_ (
    .a(N2010),
    .b(_116_),
    .y(_260_)
  );
  al_nand2ft _639_ (
    .a(_116_),
    .b(N2010),
    .y(_261_)
  );
  al_nand2 _640_ (
    .a(N1821),
    .b(N1820),
    .y(_262_)
  );
  al_nor2 _641_ (
    .a(N1821),
    .b(N1820),
    .y(_263_)
  );
  al_nand2ft _642_ (
    .a(_263_),
    .b(_262_),
    .y(_264_)
  );
  al_nand3ftt _643_ (
    .a(_260_),
    .b(_261_),
    .c(_264_),
    .y(_265_)
  );
  al_ao21ftt _644_ (
    .a(_260_),
    .b(_261_),
    .c(_264_),
    .y(_266_)
  );
  al_ao21 _645_ (
    .a(_265_),
    .b(_266_),
    .c(_259_),
    .y(_267_)
  );
  al_nand3 _646_ (
    .a(_259_),
    .b(_265_),
    .c(_266_),
    .y(_268_)
  );
  al_ao21ttf _647_ (
    .a(_268_),
    .b(_267_),
    .c(_252_),
    .y(_269_)
  );
  al_and3ftt _648_ (
    .a(_252_),
    .b(_268_),
    .c(_267_),
    .y(_270_)
  );
  al_nor3fft _649_ (
    .a(_220_),
    .b(_269_),
    .c(_270_),
    .y(N3809)
  );
  al_nor3fft _650_ (
    .a(N1726),
    .b(_083_),
    .c(_084_),
    .y(_271_)
  );
  al_and3 _651_ (
    .a(_271_),
    .b(_112_),
    .c(_068_),
    .y(_272_)
  );
  al_nor3ftt _652_ (
    .a(_272_),
    .b(N3671),
    .c(N3809),
    .y(N3881)
  );
  al_inv _653_ (
    .a(N3881),
    .y(N3882)
  );
  al_and2 _654_ (
    .a(N94),
    .b(N219),
    .y(N1026)
  );
  al_nand2 _655_ (
    .a(N241),
    .b(_157_),
    .y(N1969)
  );
  al_mux2l _656_ (
    .a(N2012),
    .b(_117_),
    .s(N246),
    .y(N2387)
  );
  al_mux2h _657_ (
    .a(N2010),
    .b(N2014),
    .s(N246),
    .y(N2389)
  );
  al_ao21ftf _658_ (
    .a(N241),
    .b(N230),
    .c(_116_),
    .y(N2496)
  );
  al_inv _659_ (
    .a(N246),
    .y(_273_)
  );
  al_nand3fft _660_ (
    .a(N230),
    .b(_273_),
    .c(_116_),
    .y(_274_)
  );
  al_aoi21ftf _661_ (
    .a(N246),
    .b(_157_),
    .c(_274_),
    .y(N2643)
  );
  al_nand3 _662_ (
    .a(N230),
    .b(_116_),
    .c(_259_),
    .y(_275_)
  );
  al_ao21ftt _663_ (
    .a(_117_),
    .b(N230),
    .c(_259_),
    .y(_276_)
  );
  al_nand3ftt _664_ (
    .a(N241),
    .b(_275_),
    .c(_276_),
    .y(_277_)
  );
  al_ao21ttf _665_ (
    .a(N241),
    .b(_256_),
    .c(_277_),
    .y(N3546)
  );
  al_and3 _666_ (
    .a(N2010),
    .b(_275_),
    .c(_276_),
    .y(_278_)
  );
  al_ao21 _667_ (
    .a(_275_),
    .b(_276_),
    .c(N2010),
    .y(_279_)
  );
  al_ao21ftt _668_ (
    .a(_278_),
    .b(_279_),
    .c(_252_),
    .y(_280_)
  );
  al_or3fft _669_ (
    .a(_252_),
    .b(_279_),
    .c(_278_),
    .y(_281_)
  );
  al_nand3 _670_ (
    .a(N246),
    .b(_281_),
    .c(_280_),
    .y(_282_)
  );
  al_aoi21ftf _671_ (
    .a(_256_),
    .b(_273_),
    .c(_282_),
    .y(N3803)
  );
  al_aoi21 _672_ (
    .a(_026_),
    .b(_126_),
    .c(N262),
    .y(_283_)
  );
  al_and3ftt _673_ (
    .a(_041_),
    .b(N40),
    .c(_045_),
    .y(_284_)
  );
  al_nand3 _674_ (
    .a(N301),
    .b(_284_),
    .c(_283_),
    .y(_285_)
  );
  al_ao21ttf _675_ (
    .a(_284_),
    .b(_283_),
    .c(N266),
    .y(_286_)
  );
  al_aoi21 _676_ (
    .a(_285_),
    .b(_286_),
    .c(N1821),
    .y(_287_)
  );
  al_inv _677_ (
    .a(N262),
    .y(_288_)
  );
  al_nand3 _678_ (
    .a(_288_),
    .b(_031_),
    .c(_284_),
    .y(_289_)
  );
  al_nand3 _679_ (
    .a(_171_),
    .b(_284_),
    .c(_283_),
    .y(_290_)
  );
  al_ao21ftf _680_ (
    .a(N259),
    .b(_289_),
    .c(_290_),
    .y(_291_)
  );
  al_nand3 _681_ (
    .a(N287),
    .b(_284_),
    .c(_283_),
    .y(_292_)
  );
  al_ao21ttf _682_ (
    .a(_284_),
    .b(_283_),
    .c(N256),
    .y(_293_)
  );
  al_nand3 _683_ (
    .a(_157_),
    .b(_292_),
    .c(_293_),
    .y(_294_)
  );
  al_ao21ttf _684_ (
    .a(_116_),
    .b(_291_),
    .c(_294_),
    .y(_295_)
  );
  al_ao21 _685_ (
    .a(_284_),
    .b(_283_),
    .c(N263),
    .y(_296_)
  );
  al_nand3ftt _686_ (
    .a(N297),
    .b(_284_),
    .c(_283_),
    .y(_297_)
  );
  al_nand3 _687_ (
    .a(N2010),
    .b(_297_),
    .c(_296_),
    .y(_298_)
  );
  al_ao21 _688_ (
    .a(_284_),
    .b(_283_),
    .c(N259),
    .y(_299_)
  );
  al_nand3ftt _689_ (
    .a(_116_),
    .b(_290_),
    .c(_299_),
    .y(_300_)
  );
  al_nand3 _690_ (
    .a(_298_),
    .b(_300_),
    .c(_295_),
    .y(_301_)
  );
  al_ao21ftf _691_ (
    .a(N263),
    .b(_289_),
    .c(_297_),
    .y(_302_)
  );
  al_nand3 _692_ (
    .a(N1821),
    .b(_285_),
    .c(_286_),
    .y(_303_)
  );
  al_aoi21ftf _693_ (
    .a(N2010),
    .b(_302_),
    .c(_303_),
    .y(_304_)
  );
  al_ao21 _694_ (
    .a(_304_),
    .b(_301_),
    .c(_287_),
    .y(_305_)
  );
  al_mux2l _695_ (
    .a(N269),
    .b(N305),
    .s(_289_),
    .y(_306_)
  );
  al_or3fft _696_ (
    .a(N8),
    .b(N1820),
    .c(_306_),
    .y(_307_)
  );
  al_inv _697_ (
    .a(N8),
    .y(_308_)
  );
  al_inv _698_ (
    .a(N309),
    .y(_309_)
  );
  al_mux2l _699_ (
    .a(_120_),
    .b(_309_),
    .s(_289_),
    .y(_310_)
  );
  al_or2 _700_ (
    .a(N1819),
    .b(_310_),
    .y(_311_)
  );
  al_nand2 _701_ (
    .a(N2014),
    .b(_306_),
    .y(_312_)
  );
  al_aoi21 _702_ (
    .a(_312_),
    .b(_311_),
    .c(_308_),
    .y(_313_)
  );
  al_ao21 _703_ (
    .a(_307_),
    .b(_305_),
    .c(_313_),
    .y(_314_)
  );
  al_nand3fft _704_ (
    .a(_308_),
    .b(N2016),
    .c(_310_),
    .y(_315_)
  );
  al_aoi21 _705_ (
    .a(_284_),
    .b(_283_),
    .c(_308_),
    .y(_316_)
  );
  al_and3 _706_ (
    .a(N275),
    .b(N2018),
    .c(_316_),
    .y(_317_)
  );
  al_ao21 _707_ (
    .a(_315_),
    .b(_314_),
    .c(_317_),
    .y(_318_)
  );
  al_and2 _708_ (
    .a(_131_),
    .b(_019_),
    .y(_319_)
  );
  al_oai21ttf _709_ (
    .a(N278),
    .b(N2020),
    .c(_319_),
    .y(_320_)
  );
  al_nand3 _710_ (
    .a(N8),
    .b(_289_),
    .c(_320_),
    .y(_321_)
  );
  al_aoi21ttf _711_ (
    .a(_288_),
    .b(_031_),
    .c(_284_),
    .y(_322_)
  );
  al_nand3 _712_ (
    .a(N287),
    .b(_183_),
    .c(_322_),
    .y(_323_)
  );
  al_and2 _713_ (
    .a(N281),
    .b(N2022),
    .y(_324_)
  );
  al_oai21ftf _714_ (
    .a(N284),
    .b(_147_),
    .c(_324_),
    .y(_325_)
  );
  al_and3fft _715_ (
    .a(N281),
    .b(N2022),
    .c(_322_),
    .y(_326_)
  );
  al_aoi21 _716_ (
    .a(_322_),
    .b(_325_),
    .c(_326_),
    .y(_327_)
  );
  al_nand3 _717_ (
    .a(N278),
    .b(N2020),
    .c(_316_),
    .y(_328_)
  );
  al_and3ftt _718_ (
    .a(_183_),
    .b(_179_),
    .c(_322_),
    .y(_329_)
  );
  al_and3 _719_ (
    .a(_140_),
    .b(_147_),
    .c(_322_),
    .y(_330_)
  );
  al_and3fft _720_ (
    .a(_329_),
    .b(_330_),
    .c(_328_),
    .y(_331_)
  );
  al_nand3 _721_ (
    .a(_323_),
    .b(_327_),
    .c(_331_),
    .y(_332_)
  );
  al_ao21 _722_ (
    .a(_321_),
    .b(_318_),
    .c(_332_),
    .y(_333_)
  );
  al_nor2 _723_ (
    .a(_140_),
    .b(_147_),
    .y(_334_)
  );
  al_nand2ft _724_ (
    .a(_334_),
    .b(_326_),
    .y(_335_)
  );
  al_nand3fft _725_ (
    .a(_329_),
    .b(_330_),
    .c(_335_),
    .y(_336_)
  );
  al_and3ftt _726_ (
    .a(_175_),
    .b(_171_),
    .c(_322_),
    .y(_337_)
  );
  al_aoi21 _727_ (
    .a(_323_),
    .b(_336_),
    .c(_337_),
    .y(_338_)
  );
  al_and3 _728_ (
    .a(N294),
    .b(_175_),
    .c(_322_),
    .y(_339_)
  );
  al_aoi21 _729_ (
    .a(_338_),
    .b(_333_),
    .c(_339_),
    .y(N3851)
  );
  assign N1034 = N1277;
  assign N1037 = N8;
  assign N1070 = N8;
  assign N1190 = N8;
  assign N1195 = N8;
  assign N143_O = N143_I;
  assign N144_O = N144_I;
  assign N145_O = N145_I;
  assign N146_O = N146_I;
  assign N147_O = N147_I;
  assign N148_O = N148_I;
  assign N149_O = N149_I;
  assign N150_O = N150_I;
  assign N1519 = N256;
  assign N151_O = N151_I;
  assign N1520 = N259;
  assign N1521 = N263;
  assign N1522 = N266;
  assign N1523 = N269;
  assign N1524 = N272;
  assign N1525 = N275;
  assign N1526 = N278;
  assign N1527 = N281;
  assign N1528 = N284;
  assign N152_O = N152_I;
  assign N153_O = N153_I;
  assign N154_O = N154_I;
  assign N155_O = N155_I;
  assign N156_O = N156_I;
  assign N1572 = N287;
  assign N1573 = N294;
  assign N1574 = N297;
  assign N1575 = N301;
  assign N1576 = N305;
  assign N1577 = N309;
  assign N157_O = N157_I;
  assign N158_O = N158_I;
  assign N1591 = N1726;
  assign N159_O = N159_I;
  assign N160_O = N160_I;
  assign N1612 = N2010;
  assign N1615 = N2012;
  assign N1619 = N2014;
  assign N161_O = N161_I;
  assign N1624 = N2016;
  assign N1628 = N2018;
  assign N162_O = N162_I;
  assign N1631 = N2020;
  assign N1634 = N2022;
  assign N163_O = N163_I;
  assign N164_O = N164_I;
  assign N165_O = N165_I;
  assign N166_O = N166_I;
  assign N167_O = N167_I;
  assign N168_O = N168_I;
  assign N169_O = N169_I;
  assign N170_O = N170_I;
  assign N171_O = N171_I;
  assign N172_O = N172_I;
  assign N173_O = N173_I;
  assign N174_O = N174_I;
  assign N175_O = N175_I;
  assign N176_O = N176_I;
  assign N177_O = N177_I;
  assign N178_O = N178_I;
  assign N179_O = N179_I;
  assign N180_O = N180_I;
  assign N181_O = N181_I;
  assign N182_O = N182_I;
  assign N183_O = N183_I;
  assign N1848 = N2010;
  assign N184_O = N184_I;
  assign N1852 = N2012;
  assign N1856 = N2014;
  assign N185_O = N185_I;
  assign N1863 = N2016;
  assign N186_O = N186_I;
  assign N1870 = N2018;
  assign N1875 = N2020;
  assign N187_O = N187_I;
  assign N1880 = N2022;
  assign N188_O = N188_I;
  assign N1897 = N1816;
  assign N189_O = N189_I;
  assign N190_O = N190_I;
  assign N191_O = N191_I;
  assign N192_O = N192_I;
  assign N193_O = N193_I;
  assign N194_O = N194_I;
  assign N195_O = N195_I;
  assign N196_O = N196_I;
  assign N197_O = N197_I;
  assign N198_O = N198_I;
  assign N199_O = N199_I;
  assign N200_O = N200_I;
  assign N201_O = N201_I;
  assign N202_O = N202_I;
  assign N203_O = N203_I;
  assign N204_O = N204_I;
  assign N205_O = N205_I;
  assign N206_O = N206_I;
  assign N207_O = N207_I;
  assign N208_O = N208_I;
  assign N209_O = N209_I;
  assign N210_O = N210_I;
  assign N211_O = N211_I;
  assign N212_O = N212_I;
  assign N2135 = N1821;
  assign N213_O = N213_I;
  assign N2141 = N1819;
  assign N214_O = N214_I;
  assign N215_O = N215_I;
  assign N216_O = N216_I;
  assign N2175 = N1818;
  assign N217_O = N217_I;
  assign N218_O = N218_I;
  assign N2194 = N1820;
  assign N2234 = N1817;
  assign N2235 = N1816;
  assign N2266 = N2387;
  assign N2269 = N2389;
  assign N2367 = N2014;
  assign N2388 = N2387;
  assign N2390 = N2389;
  assign N2437 = N1821;
  assign N2443 = N1819;
  assign N2460 = N1819;
  assign N2475 = N1821;
  assign N2481 = N1821;
  assign N2521 = N2643;
  assign N2617 = N2010;
  assign N2620 = N2012;
  assign N2628 = N2010;
  assign N2630 = N2010;
  assign N2644 = N2643;
  assign N2645 = N2012;
  assign N2655 = N2010;
  assign N2656 = N2012;
  assign N2695 = N2018;
  assign N2696 = N2016;
  assign N2697 = N2022;
  assign N2698 = N2020;
  assign N2699 = N2018;
  assign N2700 = N2016;
  assign N2701 = N2022;
  assign N2702 = N2020;
  assign N2817 = N2925;
  assign N2931 = N3038;
  assign N3600 = N3671;
  assign N3780 = N3803;
  assign N3790 = N3809;
  assign N3804 = N3803;
  assign N3840 = N3851;
  assign N3843 = N3851;
  assign N3875 = 1'b0;
  assign N3877 = N3881;
  assign N398 = N219;
  assign N400 = N219;
  assign N401 = N219;
  assign N419 = N253;
  assign N420 = N253;
  assign N456 = N290;
  assign N457 = N290;
  assign N458 = N290;
  assign N496 = N237;
  assign N500 = N219;
  assign N503 = N8;
  assign N506 = N8;
  assign N509 = N227;
  assign N521 = N234;
  assign N550 = N227;
  assign N562 = N234;
  assign N582 = N319;
  assign N594 = N322;
  assign N613 = N319;
  assign N625 = N322;
  assign N637 = N16;
  assign N643 = N16;
  assign N693 = N29;
  assign N699 = N29;
  assign N735 = N259;
  assign N738 = N256;
  assign N741 = N263;
  assign N744 = N269;
  assign N747 = N266;
  assign N750 = N275;
  assign N753 = N272;
  assign N756 = N281;
  assign N759 = N278;
  assign N762 = N287;
  assign N765 = N284;
  assign N768 = N294;
  assign N771 = N301;
  assign N774 = N297;
  assign N777 = N309;
  assign N780 = N305;
  assign N783 = N316;
  assign N786 = N313;
  assign N805 = N219;
endmodule
