
module c1355(G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  input G1;
  input G10;
  input G11;
  input G12;
  input G13;
  output G1324;
  output G1325;
  output G1326;
  output G1327;
  output G1328;
  output G1329;
  output G1330;
  output G1331;
  output G1332;
  output G1333;
  output G1334;
  output G1335;
  output G1336;
  output G1337;
  output G1338;
  output G1339;
  output G1340;
  output G1341;
  output G1342;
  output G1343;
  output G1344;
  output G1345;
  output G1346;
  output G1347;
  output G1348;
  output G1349;
  output G1350;
  output G1351;
  output G1352;
  output G1353;
  output G1354;
  output G1355;
  input G14;
  input G15;
  input G16;
  input G17;
  input G18;
  input G19;
  input G2;
  input G20;
  input G21;
  input G22;
  input G23;
  input G24;
  input G25;
  input G26;
  input G27;
  input G28;
  input G29;
  input G3;
  input G30;
  input G31;
  input G32;
  input G33;
  input G34;
  input G35;
  input G36;
  input G37;
  input G38;
  input G39;
  input G4;
  input G40;
  input G41;
  input G5;
  input G6;
  input G7;
  input G8;
  input G9;
  al_and2 _299_ (
    .a(G33),
    .b(G41),
    .y(_273_)
  );
  al_and2ft _300_ (
    .a(G19),
    .b(G20),
    .y(_274_)
  );
  al_nand2ft _301_ (
    .a(G20),
    .b(G19),
    .y(_275_)
  );
  al_nand2ft _302_ (
    .a(_274_),
    .b(_275_),
    .y(_276_)
  );
  al_nand2ft _303_ (
    .a(G18),
    .b(G17),
    .y(_277_)
  );
  al_nand2ft _304_ (
    .a(G17),
    .b(G18),
    .y(_278_)
  );
  al_ao21 _305_ (
    .a(_277_),
    .b(_278_),
    .c(_276_),
    .y(_279_)
  );
  al_nand3 _306_ (
    .a(_277_),
    .b(_278_),
    .c(_276_),
    .y(_280_)
  );
  al_and3ftt _307_ (
    .a(_273_),
    .b(_280_),
    .c(_279_),
    .y(_281_)
  );
  al_inv _308_ (
    .a(_273_),
    .y(_282_)
  );
  al_ao21 _309_ (
    .a(_280_),
    .b(_279_),
    .c(_282_),
    .y(_283_)
  );
  al_nand2ft _310_ (
    .a(_281_),
    .b(_283_),
    .y(_284_)
  );
  al_and2ft _311_ (
    .a(G23),
    .b(G24),
    .y(_285_)
  );
  al_nand2ft _312_ (
    .a(G24),
    .b(G23),
    .y(_286_)
  );
  al_and2ft _313_ (
    .a(G22),
    .b(G21),
    .y(_287_)
  );
  al_nand2ft _314_ (
    .a(G21),
    .b(G22),
    .y(_288_)
  );
  al_nand2ft _315_ (
    .a(_287_),
    .b(_288_),
    .y(_289_)
  );
  al_and3fft _316_ (
    .a(_285_),
    .b(_289_),
    .c(_286_),
    .y(_290_)
  );
  al_ao21ftf _317_ (
    .a(_285_),
    .b(_286_),
    .c(_289_),
    .y(_291_)
  );
  al_and2ft _318_ (
    .a(G13),
    .b(G9),
    .y(_292_)
  );
  al_nand2ft _319_ (
    .a(G9),
    .b(G13),
    .y(_293_)
  );
  al_and2ft _320_ (
    .a(G5),
    .b(G1),
    .y(_294_)
  );
  al_nand2ft _321_ (
    .a(G1),
    .b(G5),
    .y(_295_)
  );
  al_nand2ft _322_ (
    .a(_294_),
    .b(_295_),
    .y(_296_)
  );
  al_and3ftt _323_ (
    .a(_292_),
    .b(_293_),
    .c(_296_),
    .y(_297_)
  );
  al_ao21ftt _324_ (
    .a(_292_),
    .b(_293_),
    .c(_296_),
    .y(_298_)
  );
  al_and2ft _325_ (
    .a(_297_),
    .b(_298_),
    .y(_000_)
  );
  al_nand3ftt _326_ (
    .a(_290_),
    .b(_291_),
    .c(_000_),
    .y(_001_)
  );
  al_and3ftt _327_ (
    .a(_285_),
    .b(_286_),
    .c(_289_),
    .y(_002_)
  );
  al_aoi21ftt _328_ (
    .a(_285_),
    .b(_286_),
    .c(_289_),
    .y(_003_)
  );
  al_nand2ft _329_ (
    .a(_297_),
    .b(_298_),
    .y(_004_)
  );
  al_nand3fft _330_ (
    .a(_002_),
    .b(_003_),
    .c(_004_),
    .y(_005_)
  );
  al_aoi21ttf _331_ (
    .a(_005_),
    .b(_001_),
    .c(_284_),
    .y(_006_)
  );
  al_nand3ftt _332_ (
    .a(_290_),
    .b(_291_),
    .c(_004_),
    .y(_007_)
  );
  al_nand3fft _333_ (
    .a(_002_),
    .b(_003_),
    .c(_000_),
    .y(_008_)
  );
  al_ao21 _334_ (
    .a(_007_),
    .b(_008_),
    .c(_284_),
    .y(_009_)
  );
  al_nand2ft _335_ (
    .a(_006_),
    .b(_009_),
    .y(_010_)
  );
  al_and2ft _336_ (
    .a(G3),
    .b(G4),
    .y(_011_)
  );
  al_nand2ft _337_ (
    .a(G4),
    .b(G3),
    .y(_012_)
  );
  al_nand2ft _338_ (
    .a(_011_),
    .b(_012_),
    .y(_013_)
  );
  al_nand2ft _339_ (
    .a(G2),
    .b(G1),
    .y(_014_)
  );
  al_nand2ft _340_ (
    .a(G1),
    .b(G2),
    .y(_015_)
  );
  al_ao21 _341_ (
    .a(_014_),
    .b(_015_),
    .c(_013_),
    .y(_016_)
  );
  al_nand3 _342_ (
    .a(_014_),
    .b(_015_),
    .c(_013_),
    .y(_017_)
  );
  al_nand2 _343_ (
    .a(G41),
    .b(G37),
    .y(_018_)
  );
  al_and3 _344_ (
    .a(_018_),
    .b(_017_),
    .c(_016_),
    .y(_019_)
  );
  al_ao21 _345_ (
    .a(_017_),
    .b(_016_),
    .c(_018_),
    .y(_020_)
  );
  al_nand2ft _346_ (
    .a(_019_),
    .b(_020_),
    .y(_021_)
  );
  al_and2ft _347_ (
    .a(G7),
    .b(G8),
    .y(_022_)
  );
  al_nand2ft _348_ (
    .a(G8),
    .b(G7),
    .y(_023_)
  );
  al_and2ft _349_ (
    .a(G6),
    .b(G5),
    .y(_024_)
  );
  al_nand2ft _350_ (
    .a(G5),
    .b(G6),
    .y(_025_)
  );
  al_nand2ft _351_ (
    .a(_024_),
    .b(_025_),
    .y(_026_)
  );
  al_and3fft _352_ (
    .a(_022_),
    .b(_026_),
    .c(_023_),
    .y(_027_)
  );
  al_aoi21ftf _353_ (
    .a(_022_),
    .b(_023_),
    .c(_026_),
    .y(_028_)
  );
  al_or2 _354_ (
    .a(_028_),
    .b(_027_),
    .y(_029_)
  );
  al_and2ft _355_ (
    .a(G21),
    .b(G17),
    .y(_030_)
  );
  al_and2ft _356_ (
    .a(G17),
    .b(G21),
    .y(_031_)
  );
  al_and2ft _357_ (
    .a(G29),
    .b(G25),
    .y(_032_)
  );
  al_nand2ft _358_ (
    .a(G25),
    .b(G29),
    .y(_033_)
  );
  al_nand2ft _359_ (
    .a(_032_),
    .b(_033_),
    .y(_034_)
  );
  al_oa21ttf _360_ (
    .a(_030_),
    .b(_031_),
    .c(_034_),
    .y(_035_)
  );
  al_nand3fft _361_ (
    .a(_030_),
    .b(_031_),
    .c(_034_),
    .y(_036_)
  );
  al_ao21ftt _362_ (
    .a(_035_),
    .b(_036_),
    .c(_029_),
    .y(_037_)
  );
  al_nand3ftt _363_ (
    .a(_035_),
    .b(_036_),
    .c(_029_),
    .y(_038_)
  );
  al_nand3 _364_ (
    .a(_037_),
    .b(_021_),
    .c(_038_),
    .y(_039_)
  );
  al_aoi21 _365_ (
    .a(_038_),
    .b(_037_),
    .c(_021_),
    .y(_040_)
  );
  al_nand2ft _366_ (
    .a(_040_),
    .b(_039_),
    .y(_041_)
  );
  al_and2ft _367_ (
    .a(G11),
    .b(G12),
    .y(_042_)
  );
  al_nand2ft _368_ (
    .a(G12),
    .b(G11),
    .y(_043_)
  );
  al_and2ft _369_ (
    .a(G10),
    .b(G9),
    .y(_044_)
  );
  al_nand2ft _370_ (
    .a(G9),
    .b(G10),
    .y(_045_)
  );
  al_nand2ft _371_ (
    .a(_044_),
    .b(_045_),
    .y(_046_)
  );
  al_and3ftt _372_ (
    .a(_042_),
    .b(_043_),
    .c(_046_),
    .y(_047_)
  );
  al_aoi21ftt _373_ (
    .a(_042_),
    .b(_043_),
    .c(_046_),
    .y(_048_)
  );
  al_nand2 _374_ (
    .a(G41),
    .b(G38),
    .y(_049_)
  );
  al_nor3ftt _375_ (
    .a(_049_),
    .b(_047_),
    .c(_048_),
    .y(_050_)
  );
  al_and3fft _376_ (
    .a(_042_),
    .b(_046_),
    .c(_043_),
    .y(_051_)
  );
  al_aoi21ftf _377_ (
    .a(_042_),
    .b(_043_),
    .c(_046_),
    .y(_052_)
  );
  al_or3 _378_ (
    .a(_049_),
    .b(_052_),
    .c(_051_),
    .y(_053_)
  );
  al_and2ft _379_ (
    .a(_050_),
    .b(_053_),
    .y(_054_)
  );
  al_and2ft _380_ (
    .a(G15),
    .b(G16),
    .y(_055_)
  );
  al_nand2ft _381_ (
    .a(G16),
    .b(G15),
    .y(_056_)
  );
  al_and2ft _382_ (
    .a(G14),
    .b(G13),
    .y(_057_)
  );
  al_nand2ft _383_ (
    .a(G13),
    .b(G14),
    .y(_058_)
  );
  al_nand2ft _384_ (
    .a(_057_),
    .b(_058_),
    .y(_059_)
  );
  al_and3ftt _385_ (
    .a(_055_),
    .b(_056_),
    .c(_059_),
    .y(_060_)
  );
  al_aoi21ftt _386_ (
    .a(_055_),
    .b(_056_),
    .c(_059_),
    .y(_061_)
  );
  al_or2 _387_ (
    .a(_060_),
    .b(_061_),
    .y(_062_)
  );
  al_and2ft _388_ (
    .a(G22),
    .b(G18),
    .y(_063_)
  );
  al_nand2ft _389_ (
    .a(G18),
    .b(G22),
    .y(_064_)
  );
  al_nand2ft _390_ (
    .a(_063_),
    .b(_064_),
    .y(_065_)
  );
  al_and2ft _391_ (
    .a(G30),
    .b(G26),
    .y(_066_)
  );
  al_nand2ft _392_ (
    .a(G26),
    .b(G30),
    .y(_067_)
  );
  al_and3ftt _393_ (
    .a(_066_),
    .b(_067_),
    .c(_065_),
    .y(_068_)
  );
  al_ao21ftt _394_ (
    .a(_066_),
    .b(_067_),
    .c(_065_),
    .y(_069_)
  );
  al_nand3ftt _395_ (
    .a(_068_),
    .b(_069_),
    .c(_062_),
    .y(_070_)
  );
  al_nor2 _396_ (
    .a(_060_),
    .b(_061_),
    .y(_071_)
  );
  al_ao21ftf _397_ (
    .a(_068_),
    .b(_069_),
    .c(_071_),
    .y(_072_)
  );
  al_ao21 _398_ (
    .a(_070_),
    .b(_072_),
    .c(_054_),
    .y(_073_)
  );
  al_nand3 _399_ (
    .a(_070_),
    .b(_072_),
    .c(_054_),
    .y(_074_)
  );
  al_and3 _400_ (
    .a(_073_),
    .b(_074_),
    .c(_041_),
    .y(_075_)
  );
  al_and2 _401_ (
    .a(G41),
    .b(G39),
    .y(_076_)
  );
  al_ao21 _402_ (
    .a(_017_),
    .b(_016_),
    .c(_076_),
    .y(_077_)
  );
  al_and3 _403_ (
    .a(_076_),
    .b(_017_),
    .c(_016_),
    .y(_078_)
  );
  al_nand2ft _404_ (
    .a(_078_),
    .b(_077_),
    .y(_079_)
  );
  al_nand2 _405_ (
    .a(G19),
    .b(G23),
    .y(_080_)
  );
  al_or2 _406_ (
    .a(G19),
    .b(G23),
    .y(_081_)
  );
  al_and2ft _407_ (
    .a(G31),
    .b(G27),
    .y(_082_)
  );
  al_nand2ft _408_ (
    .a(G27),
    .b(G31),
    .y(_083_)
  );
  al_nand2ft _409_ (
    .a(_082_),
    .b(_083_),
    .y(_084_)
  );
  al_ao21 _410_ (
    .a(_080_),
    .b(_081_),
    .c(_084_),
    .y(_085_)
  );
  al_and3 _411_ (
    .a(_080_),
    .b(_081_),
    .c(_084_),
    .y(_086_)
  );
  al_nand2ft _412_ (
    .a(_086_),
    .b(_085_),
    .y(_087_)
  );
  al_nand3fft _413_ (
    .a(_051_),
    .b(_052_),
    .c(_087_),
    .y(_088_)
  );
  al_and2ft _414_ (
    .a(_086_),
    .b(_085_),
    .y(_089_)
  );
  al_nand3fft _415_ (
    .a(_047_),
    .b(_048_),
    .c(_089_),
    .y(_090_)
  );
  al_aoi21 _416_ (
    .a(_088_),
    .b(_090_),
    .c(_079_),
    .y(_091_)
  );
  al_nand3 _417_ (
    .a(_088_),
    .b(_079_),
    .c(_090_),
    .y(_092_)
  );
  al_nand2ft _418_ (
    .a(_091_),
    .b(_092_),
    .y(_093_)
  );
  al_ao21ftf _419_ (
    .a(_022_),
    .b(_023_),
    .c(_026_),
    .y(_094_)
  );
  al_and2 _420_ (
    .a(G41),
    .b(G40),
    .y(_095_)
  );
  al_oai21ftf _421_ (
    .a(_094_),
    .b(_027_),
    .c(_095_),
    .y(_096_)
  );
  al_nor3fft _422_ (
    .a(_095_),
    .b(_094_),
    .c(_027_),
    .y(_097_)
  );
  al_nand2ft _423_ (
    .a(_097_),
    .b(_096_),
    .y(_098_)
  );
  al_and2ft _424_ (
    .a(G24),
    .b(G20),
    .y(_099_)
  );
  al_nand2ft _425_ (
    .a(G20),
    .b(G24),
    .y(_100_)
  );
  al_nand2ft _426_ (
    .a(_099_),
    .b(_100_),
    .y(_101_)
  );
  al_and2ft _427_ (
    .a(G32),
    .b(G28),
    .y(_102_)
  );
  al_nand2ft _428_ (
    .a(G28),
    .b(G32),
    .y(_103_)
  );
  al_and3ftt _429_ (
    .a(_102_),
    .b(_103_),
    .c(_101_),
    .y(_104_)
  );
  al_ao21ftt _430_ (
    .a(_102_),
    .b(_103_),
    .c(_101_),
    .y(_105_)
  );
  al_ao21ftf _431_ (
    .a(_104_),
    .b(_105_),
    .c(_062_),
    .y(_106_)
  );
  al_nand3ftt _432_ (
    .a(_104_),
    .b(_105_),
    .c(_071_),
    .y(_107_)
  );
  al_nand3 _433_ (
    .a(_106_),
    .b(_098_),
    .c(_107_),
    .y(_108_)
  );
  al_ao21 _434_ (
    .a(_106_),
    .b(_107_),
    .c(_098_),
    .y(_109_)
  );
  al_and3 _435_ (
    .a(_108_),
    .b(_109_),
    .c(_093_),
    .y(_110_)
  );
  al_nand2 _436_ (
    .a(G41),
    .b(G35),
    .y(_111_)
  );
  al_and3 _437_ (
    .a(_111_),
    .b(_280_),
    .c(_279_),
    .y(_112_)
  );
  al_ao21 _438_ (
    .a(_280_),
    .b(_279_),
    .c(_111_),
    .y(_113_)
  );
  al_nand2ft _439_ (
    .a(_112_),
    .b(_113_),
    .y(_114_)
  );
  al_and2ft _440_ (
    .a(G27),
    .b(G28),
    .y(_115_)
  );
  al_nand2ft _441_ (
    .a(G28),
    .b(G27),
    .y(_116_)
  );
  al_and2ft _442_ (
    .a(G26),
    .b(G25),
    .y(_117_)
  );
  al_nand2ft _443_ (
    .a(G25),
    .b(G26),
    .y(_118_)
  );
  al_nand2ft _444_ (
    .a(_117_),
    .b(_118_),
    .y(_119_)
  );
  al_and3ftt _445_ (
    .a(_115_),
    .b(_116_),
    .c(_119_),
    .y(_120_)
  );
  al_aoi21ftt _446_ (
    .a(_115_),
    .b(_116_),
    .c(_119_),
    .y(_121_)
  );
  al_or2 _447_ (
    .a(_120_),
    .b(_121_),
    .y(_122_)
  );
  al_and2ft _448_ (
    .a(G7),
    .b(G3),
    .y(_123_)
  );
  al_nand2ft _449_ (
    .a(G3),
    .b(G7),
    .y(_124_)
  );
  al_nand2ft _450_ (
    .a(_123_),
    .b(_124_),
    .y(_125_)
  );
  al_and2ft _451_ (
    .a(G15),
    .b(G11),
    .y(_126_)
  );
  al_nand2ft _452_ (
    .a(G11),
    .b(G15),
    .y(_127_)
  );
  al_and3ftt _453_ (
    .a(_126_),
    .b(_127_),
    .c(_125_),
    .y(_128_)
  );
  al_ao21ftt _454_ (
    .a(_126_),
    .b(_127_),
    .c(_125_),
    .y(_129_)
  );
  al_ao21ftf _455_ (
    .a(_128_),
    .b(_129_),
    .c(_122_),
    .y(_130_)
  );
  al_nor2 _456_ (
    .a(_120_),
    .b(_121_),
    .y(_131_)
  );
  al_nand3ftt _457_ (
    .a(_128_),
    .b(_129_),
    .c(_131_),
    .y(_132_)
  );
  al_nand3 _458_ (
    .a(_130_),
    .b(_132_),
    .c(_114_),
    .y(_133_)
  );
  al_aoi21 _459_ (
    .a(_130_),
    .b(_132_),
    .c(_114_),
    .y(_134_)
  );
  al_nand2ft _460_ (
    .a(_134_),
    .b(_133_),
    .y(_135_)
  );
  al_and2 _461_ (
    .a(G41),
    .b(G34),
    .y(_136_)
  );
  al_and2ft _462_ (
    .a(G31),
    .b(G32),
    .y(_137_)
  );
  al_nand2ft _463_ (
    .a(G32),
    .b(G31),
    .y(_138_)
  );
  al_and2ft _464_ (
    .a(G30),
    .b(G29),
    .y(_139_)
  );
  al_nand2ft _465_ (
    .a(G29),
    .b(G30),
    .y(_140_)
  );
  al_nand2ft _466_ (
    .a(_139_),
    .b(_140_),
    .y(_141_)
  );
  al_nand3ftt _467_ (
    .a(_137_),
    .b(_138_),
    .c(_141_),
    .y(_142_)
  );
  al_aoi21ftt _468_ (
    .a(_137_),
    .b(_138_),
    .c(_141_),
    .y(_143_)
  );
  al_and3fft _469_ (
    .a(_136_),
    .b(_143_),
    .c(_142_),
    .y(_144_)
  );
  al_and3fft _470_ (
    .a(_137_),
    .b(_141_),
    .c(_138_),
    .y(_145_)
  );
  al_ao21ftf _471_ (
    .a(_137_),
    .b(_138_),
    .c(_141_),
    .y(_146_)
  );
  al_or3fft _472_ (
    .a(_136_),
    .b(_146_),
    .c(_145_),
    .y(_147_)
  );
  al_or2ft _473_ (
    .a(_147_),
    .b(_144_),
    .y(_148_)
  );
  al_and2ft _474_ (
    .a(G14),
    .b(G10),
    .y(_149_)
  );
  al_nand2ft _475_ (
    .a(G10),
    .b(G14),
    .y(_150_)
  );
  al_nand2ft _476_ (
    .a(_149_),
    .b(_150_),
    .y(_151_)
  );
  al_nand2 _477_ (
    .a(G2),
    .b(G6),
    .y(_152_)
  );
  al_nor2 _478_ (
    .a(G2),
    .b(G6),
    .y(_153_)
  );
  al_and3fft _479_ (
    .a(_153_),
    .b(_151_),
    .c(_152_),
    .y(_154_)
  );
  al_ao21ftf _480_ (
    .a(_153_),
    .b(_152_),
    .c(_151_),
    .y(_155_)
  );
  al_nand3ftt _481_ (
    .a(_154_),
    .b(_155_),
    .c(_122_),
    .y(_156_)
  );
  al_ao21ftf _482_ (
    .a(_154_),
    .b(_155_),
    .c(_131_),
    .y(_157_)
  );
  al_and3 _483_ (
    .a(_156_),
    .b(_148_),
    .c(_157_),
    .y(_158_)
  );
  al_ao21 _484_ (
    .a(_156_),
    .b(_157_),
    .c(_148_),
    .y(_159_)
  );
  al_or2ft _485_ (
    .a(_159_),
    .b(_158_),
    .y(_160_)
  );
  al_or3 _486_ (
    .a(_010_),
    .b(_160_),
    .c(_135_),
    .y(_161_)
  );
  al_aoi21ftf _487_ (
    .a(_158_),
    .b(_159_),
    .c(_010_),
    .y(_162_)
  );
  al_ao21ftf _488_ (
    .a(_135_),
    .b(_162_),
    .c(_161_),
    .y(_163_)
  );
  al_and2 _489_ (
    .a(G41),
    .b(G36),
    .y(_164_)
  );
  al_and3fft _490_ (
    .a(_164_),
    .b(_290_),
    .c(_291_),
    .y(_165_)
  );
  al_or3ftt _491_ (
    .a(_164_),
    .b(_002_),
    .c(_003_),
    .y(_166_)
  );
  al_nand2ft _492_ (
    .a(_165_),
    .b(_166_),
    .y(_167_)
  );
  al_and2ft _493_ (
    .a(G8),
    .b(G4),
    .y(_168_)
  );
  al_nand2ft _494_ (
    .a(G4),
    .b(G8),
    .y(_169_)
  );
  al_nand2ft _495_ (
    .a(_168_),
    .b(_169_),
    .y(_170_)
  );
  al_and2ft _496_ (
    .a(G16),
    .b(G12),
    .y(_171_)
  );
  al_nand2ft _497_ (
    .a(G12),
    .b(G16),
    .y(_172_)
  );
  al_and3ftt _498_ (
    .a(_171_),
    .b(_172_),
    .c(_170_),
    .y(_173_)
  );
  al_ao21ftt _499_ (
    .a(_171_),
    .b(_172_),
    .c(_170_),
    .y(_174_)
  );
  al_nand2ft _500_ (
    .a(_173_),
    .b(_174_),
    .y(_175_)
  );
  al_or3ftt _501_ (
    .a(_146_),
    .b(_145_),
    .c(_175_),
    .y(_176_)
  );
  al_nand3ftt _502_ (
    .a(_143_),
    .b(_142_),
    .c(_175_),
    .y(_177_)
  );
  al_ao21 _503_ (
    .a(_177_),
    .b(_176_),
    .c(_167_),
    .y(_178_)
  );
  al_nand3 _504_ (
    .a(_177_),
    .b(_167_),
    .c(_176_),
    .y(_179_)
  );
  al_and2 _505_ (
    .a(_178_),
    .b(_179_),
    .y(_180_)
  );
  al_and3 _506_ (
    .a(_178_),
    .b(_179_),
    .c(_135_),
    .y(_181_)
  );
  al_ao21 _507_ (
    .a(_178_),
    .b(_179_),
    .c(_135_),
    .y(_182_)
  );
  al_and3ftt _508_ (
    .a(_006_),
    .b(_009_),
    .c(_160_),
    .y(_183_)
  );
  al_oa21ftt _509_ (
    .a(_182_),
    .b(_181_),
    .c(_183_),
    .y(_184_)
  );
  al_ao21 _510_ (
    .a(_180_),
    .b(_163_),
    .c(_184_),
    .y(_185_)
  );
  al_and3 _511_ (
    .a(_075_),
    .b(_110_),
    .c(_185_),
    .y(_186_)
  );
  al_and3 _512_ (
    .a(G1),
    .b(_010_),
    .c(_186_),
    .y(_187_)
  );
  al_ao21 _513_ (
    .a(_010_),
    .b(_186_),
    .c(G1),
    .y(_188_)
  );
  al_nand2ft _514_ (
    .a(_187_),
    .b(_188_),
    .y(G1324)
  );
  al_inv _515_ (
    .a(_160_),
    .y(_189_)
  );
  al_and3 _516_ (
    .a(G2),
    .b(_189_),
    .c(_186_),
    .y(_190_)
  );
  al_ao21 _517_ (
    .a(_189_),
    .b(_186_),
    .c(G2),
    .y(_191_)
  );
  al_nand2ft _518_ (
    .a(_190_),
    .b(_191_),
    .y(G1325)
  );
  al_ao21 _519_ (
    .a(_135_),
    .b(_186_),
    .c(G3),
    .y(_192_)
  );
  al_and3 _520_ (
    .a(G3),
    .b(_135_),
    .c(_186_),
    .y(_193_)
  );
  al_nand2ft _521_ (
    .a(_193_),
    .b(_192_),
    .y(G1326)
  );
  al_ao21ftt _522_ (
    .a(_180_),
    .b(_186_),
    .c(G4),
    .y(_194_)
  );
  al_and3ftt _523_ (
    .a(_180_),
    .b(G4),
    .c(_186_),
    .y(_195_)
  );
  al_nand2ft _524_ (
    .a(_195_),
    .b(_194_),
    .y(G1327)
  );
  al_nand2 _525_ (
    .a(_109_),
    .b(_108_),
    .y(_196_)
  );
  al_nand3ftt _526_ (
    .a(_091_),
    .b(_092_),
    .c(_196_),
    .y(_197_)
  );
  al_inv _527_ (
    .a(_197_),
    .y(_198_)
  );
  al_and3 _528_ (
    .a(_075_),
    .b(_198_),
    .c(_185_),
    .y(_199_)
  );
  al_and3 _529_ (
    .a(G5),
    .b(_010_),
    .c(_199_),
    .y(_200_)
  );
  al_ao21 _530_ (
    .a(_010_),
    .b(_199_),
    .c(G5),
    .y(_201_)
  );
  al_nand2ft _531_ (
    .a(_200_),
    .b(_201_),
    .y(G1328)
  );
  al_and3 _532_ (
    .a(G6),
    .b(_189_),
    .c(_199_),
    .y(_202_)
  );
  al_ao21 _533_ (
    .a(_189_),
    .b(_199_),
    .c(G6),
    .y(_203_)
  );
  al_nand2ft _534_ (
    .a(_202_),
    .b(_203_),
    .y(G1329)
  );
  al_ao21 _535_ (
    .a(_135_),
    .b(_199_),
    .c(G7),
    .y(_204_)
  );
  al_and3 _536_ (
    .a(G7),
    .b(_135_),
    .c(_199_),
    .y(_205_)
  );
  al_nand2ft _537_ (
    .a(_205_),
    .b(_204_),
    .y(G1330)
  );
  al_ao21ftt _538_ (
    .a(_180_),
    .b(_199_),
    .c(G8),
    .y(_206_)
  );
  al_and3ftt _539_ (
    .a(_180_),
    .b(G8),
    .c(_199_),
    .y(_207_)
  );
  al_nand2ft _540_ (
    .a(_207_),
    .b(_206_),
    .y(G1331)
  );
  al_nand2 _541_ (
    .a(_073_),
    .b(_074_),
    .y(_208_)
  );
  al_and3ftt _542_ (
    .a(_040_),
    .b(_039_),
    .c(_208_),
    .y(_209_)
  );
  al_and3 _543_ (
    .a(_110_),
    .b(_209_),
    .c(_185_),
    .y(_210_)
  );
  al_and3 _544_ (
    .a(G9),
    .b(_010_),
    .c(_210_),
    .y(_211_)
  );
  al_ao21 _545_ (
    .a(_010_),
    .b(_210_),
    .c(G9),
    .y(_212_)
  );
  al_nand2ft _546_ (
    .a(_211_),
    .b(_212_),
    .y(G1332)
  );
  al_and3 _547_ (
    .a(G10),
    .b(_189_),
    .c(_210_),
    .y(_213_)
  );
  al_ao21 _548_ (
    .a(_189_),
    .b(_210_),
    .c(G10),
    .y(_214_)
  );
  al_nand2ft _549_ (
    .a(_213_),
    .b(_214_),
    .y(G1333)
  );
  al_ao21 _550_ (
    .a(_135_),
    .b(_210_),
    .c(G11),
    .y(_215_)
  );
  al_and3 _551_ (
    .a(G11),
    .b(_135_),
    .c(_210_),
    .y(_216_)
  );
  al_nand2ft _552_ (
    .a(_216_),
    .b(_215_),
    .y(G1334)
  );
  al_ao21ftt _553_ (
    .a(_180_),
    .b(_210_),
    .c(G12),
    .y(_217_)
  );
  al_and3ftt _554_ (
    .a(_180_),
    .b(G12),
    .c(_210_),
    .y(_218_)
  );
  al_nand2ft _555_ (
    .a(_218_),
    .b(_217_),
    .y(G1335)
  );
  al_and3 _556_ (
    .a(_198_),
    .b(_209_),
    .c(_185_),
    .y(_219_)
  );
  al_ao21 _557_ (
    .a(_010_),
    .b(_219_),
    .c(G13),
    .y(_220_)
  );
  al_and3 _558_ (
    .a(G13),
    .b(_010_),
    .c(_219_),
    .y(_221_)
  );
  al_nand2ft _559_ (
    .a(_221_),
    .b(_220_),
    .y(G1336)
  );
  al_ao21 _560_ (
    .a(_189_),
    .b(_219_),
    .c(G14),
    .y(_222_)
  );
  al_and3 _561_ (
    .a(G14),
    .b(_189_),
    .c(_219_),
    .y(_223_)
  );
  al_nand2ft _562_ (
    .a(_223_),
    .b(_222_),
    .y(G1337)
  );
  al_ao21 _563_ (
    .a(_135_),
    .b(_219_),
    .c(G15),
    .y(_224_)
  );
  al_and3 _564_ (
    .a(G15),
    .b(_135_),
    .c(_219_),
    .y(_225_)
  );
  al_nand2ft _565_ (
    .a(_225_),
    .b(_224_),
    .y(G1338)
  );
  al_ao21ftt _566_ (
    .a(_180_),
    .b(_219_),
    .c(G16),
    .y(_226_)
  );
  al_and3ftt _567_ (
    .a(_180_),
    .b(G16),
    .c(_219_),
    .y(_227_)
  );
  al_nand2ft _568_ (
    .a(_227_),
    .b(_226_),
    .y(G1339)
  );
  al_or3fft _569_ (
    .a(_108_),
    .b(_109_),
    .c(_093_),
    .y(_228_)
  );
  al_oai21ttf _570_ (
    .a(_075_),
    .b(_209_),
    .c(_228_),
    .y(_229_)
  );
  al_nand2ft _571_ (
    .a(_110_),
    .b(_197_),
    .y(_230_)
  );
  al_nor3fft _572_ (
    .a(_073_),
    .b(_074_),
    .c(_041_),
    .y(_231_)
  );
  al_ao21ttf _573_ (
    .a(_231_),
    .b(_230_),
    .c(_229_),
    .y(_232_)
  );
  al_and3 _574_ (
    .a(_162_),
    .b(_181_),
    .c(_232_),
    .y(_233_)
  );
  al_ao21 _575_ (
    .a(_041_),
    .b(_233_),
    .c(G17),
    .y(_234_)
  );
  al_and3 _576_ (
    .a(G17),
    .b(_041_),
    .c(_233_),
    .y(_235_)
  );
  al_nand2ft _577_ (
    .a(_235_),
    .b(_234_),
    .y(G1340)
  );
  al_ao21 _578_ (
    .a(_208_),
    .b(_233_),
    .c(G18),
    .y(_236_)
  );
  al_and3 _579_ (
    .a(G18),
    .b(_208_),
    .c(_233_),
    .y(_237_)
  );
  al_nand2ft _580_ (
    .a(_237_),
    .b(_236_),
    .y(G1341)
  );
  al_ao21 _581_ (
    .a(_093_),
    .b(_233_),
    .c(G19),
    .y(_238_)
  );
  al_and3 _582_ (
    .a(G19),
    .b(_093_),
    .c(_233_),
    .y(_239_)
  );
  al_nand2ft _583_ (
    .a(_239_),
    .b(_238_),
    .y(G1342)
  );
  al_ao21 _584_ (
    .a(_196_),
    .b(_233_),
    .c(G20),
    .y(_240_)
  );
  al_and3 _585_ (
    .a(G20),
    .b(_196_),
    .c(_233_),
    .y(_241_)
  );
  al_nand2ft _586_ (
    .a(_241_),
    .b(_240_),
    .y(G1343)
  );
  al_oai21ftt _587_ (
    .a(_197_),
    .b(_110_),
    .c(_231_),
    .y(_242_)
  );
  al_or3ftt _588_ (
    .a(_162_),
    .b(_135_),
    .c(_180_),
    .y(_243_)
  );
  al_aoi21 _589_ (
    .a(_242_),
    .b(_229_),
    .c(_243_),
    .y(_244_)
  );
  al_ao21 _590_ (
    .a(_041_),
    .b(_244_),
    .c(G21),
    .y(_245_)
  );
  al_and3 _591_ (
    .a(G21),
    .b(_041_),
    .c(_244_),
    .y(_246_)
  );
  al_nand2ft _592_ (
    .a(_246_),
    .b(_245_),
    .y(G1344)
  );
  al_ao21 _593_ (
    .a(_208_),
    .b(_244_),
    .c(G22),
    .y(_247_)
  );
  al_and3 _594_ (
    .a(G22),
    .b(_208_),
    .c(_244_),
    .y(_248_)
  );
  al_nand2ft _595_ (
    .a(_248_),
    .b(_247_),
    .y(G1345)
  );
  al_ao21 _596_ (
    .a(_093_),
    .b(_244_),
    .c(G23),
    .y(_249_)
  );
  al_and3 _597_ (
    .a(G23),
    .b(_093_),
    .c(_244_),
    .y(_250_)
  );
  al_nand2ft _598_ (
    .a(_250_),
    .b(_249_),
    .y(G1346)
  );
  al_ao21 _599_ (
    .a(_196_),
    .b(_244_),
    .c(G24),
    .y(_251_)
  );
  al_and3 _600_ (
    .a(G24),
    .b(_196_),
    .c(_244_),
    .y(_252_)
  );
  al_nand2ft _601_ (
    .a(_252_),
    .b(_251_),
    .y(G1347)
  );
  al_and3fft _602_ (
    .a(_158_),
    .b(_010_),
    .c(_159_),
    .y(_253_)
  );
  al_and3 _603_ (
    .a(_253_),
    .b(_181_),
    .c(_232_),
    .y(_254_)
  );
  al_ao21 _604_ (
    .a(_041_),
    .b(_254_),
    .c(G25),
    .y(_255_)
  );
  al_and3 _605_ (
    .a(G25),
    .b(_041_),
    .c(_254_),
    .y(_256_)
  );
  al_nand2ft _606_ (
    .a(_256_),
    .b(_255_),
    .y(G1348)
  );
  al_ao21 _607_ (
    .a(_208_),
    .b(_254_),
    .c(G26),
    .y(_257_)
  );
  al_and3 _608_ (
    .a(G26),
    .b(_208_),
    .c(_254_),
    .y(_258_)
  );
  al_nand2ft _609_ (
    .a(_258_),
    .b(_257_),
    .y(G1349)
  );
  al_ao21 _610_ (
    .a(_093_),
    .b(_254_),
    .c(G27),
    .y(_259_)
  );
  al_and3 _611_ (
    .a(G27),
    .b(_093_),
    .c(_254_),
    .y(_260_)
  );
  al_nand2ft _612_ (
    .a(_260_),
    .b(_259_),
    .y(G1350)
  );
  al_ao21 _613_ (
    .a(_196_),
    .b(_254_),
    .c(G28),
    .y(_261_)
  );
  al_and3 _614_ (
    .a(G28),
    .b(_196_),
    .c(_254_),
    .y(_262_)
  );
  al_nand2ft _615_ (
    .a(_262_),
    .b(_261_),
    .y(G1351)
  );
  al_or2 _616_ (
    .a(_180_),
    .b(_161_),
    .y(_263_)
  );
  al_aoi21 _617_ (
    .a(_242_),
    .b(_229_),
    .c(_263_),
    .y(_264_)
  );
  al_ao21 _618_ (
    .a(_041_),
    .b(_264_),
    .c(G29),
    .y(_265_)
  );
  al_and3 _619_ (
    .a(G29),
    .b(_041_),
    .c(_264_),
    .y(_266_)
  );
  al_nand2ft _620_ (
    .a(_266_),
    .b(_265_),
    .y(G1352)
  );
  al_ao21 _621_ (
    .a(_208_),
    .b(_264_),
    .c(G30),
    .y(_267_)
  );
  al_and3 _622_ (
    .a(G30),
    .b(_208_),
    .c(_264_),
    .y(_268_)
  );
  al_nand2ft _623_ (
    .a(_268_),
    .b(_267_),
    .y(G1353)
  );
  al_ao21 _624_ (
    .a(_093_),
    .b(_264_),
    .c(G31),
    .y(_269_)
  );
  al_and3 _625_ (
    .a(G31),
    .b(_093_),
    .c(_264_),
    .y(_270_)
  );
  al_nand2ft _626_ (
    .a(_270_),
    .b(_269_),
    .y(G1354)
  );
  al_ao21 _627_ (
    .a(_196_),
    .b(_264_),
    .c(G32),
    .y(_271_)
  );
  al_and3 _628_ (
    .a(G32),
    .b(_196_),
    .c(_264_),
    .y(_272_)
  );
  al_nand2ft _629_ (
    .a(_272_),
    .b(_271_),
    .y(G1355)
  );
endmodule
