
module s15850(GND, VDD, CK, g100, g101, g102, g103, g10377, g10379, g104, g10455, g10457, g10459, g10461, g10463, g10465, g10628, g10801, g109, g11163, g11206, g11489, g1170, g1173, g1176, g1179, g1182, g1185, g1188, g1191, g1194, g1197, g1200, g1203, g1696, g1700, g1712, g18, g1957, g1960, g1961, g23, g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612, g2648, g27, g28, g29, g2986, g30, g3007, g3069, g31, g3327, g41, g4171, g4172, g4173, g4174, g4175, g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194, g4195, g4196, g4197, g4198, g4199, g42, g4200, g4201, g4202, g4203, g4204, g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, g4214, g4215, g4216, g43, g44, g45, g46, g47, g48, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6253, g6254, g6255, g6256, g6257, g6258, g6259, g6260, g6261, g6262, g6263, g6264, g6265, g6266, g6267, g6268, g6269, g6270, g6271, g6272, g6273, g6274, g6275, g6276, g6277, g6278, g6279, g6280, g6281, g6282, g6283, g6284, g6285, g6842, g6920, g6926, g6932, g6942, g6949, g6955, g741, g742, g743, g744, g750, g7744, g8061, g8062, g82, g8271, g83, g8313, g8316, g8318, g8323, g8328, g8331, g8335, g8340, g8347, g8349, g8352, g84, g85, g8561, g8562, g8563, g8564, g8565, g8566, g86, g87, g872, g873, g877, g88, g881, g886, g889, g89, g892, g895, g8976, g8977, g8978, g8979, g898, g8980, g8981, g8982, g8983, g8984, g8985, g8986, g90, g901, g904, g907, g91, g910, g913, g916, g919, g92, g922, g925, g93, g94, g9451, g95, g96, g99, g9961);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  input CK;
  wire \DFF_0.CK ;
  wire \DFF_0.D ;
  wire \DFF_0.Q ;
  wire \DFF_1.CK ;
  wire \DFF_1.D ;
  wire \DFF_1.Q ;
  wire \DFF_10.CK ;
  wire \DFF_10.D ;
  wire \DFF_10.Q ;
  wire \DFF_100.CK ;
  wire \DFF_100.D ;
  wire \DFF_100.Q ;
  wire \DFF_101.CK ;
  wire \DFF_101.D ;
  wire \DFF_101.Q ;
  wire \DFF_102.CK ;
  wire \DFF_102.D ;
  wire \DFF_102.Q ;
  wire \DFF_103.CK ;
  wire \DFF_103.D ;
  wire \DFF_103.Q ;
  wire \DFF_104.CK ;
  wire \DFF_104.D ;
  wire \DFF_104.Q ;
  wire \DFF_105.CK ;
  wire \DFF_105.D ;
  wire \DFF_105.Q ;
  wire \DFF_106.CK ;
  wire \DFF_106.D ;
  wire \DFF_106.Q ;
  wire \DFF_107.CK ;
  wire \DFF_108.CK ;
  wire \DFF_108.D ;
  wire \DFF_108.Q ;
  wire \DFF_109.CK ;
  wire \DFF_109.D ;
  wire \DFF_109.Q ;
  wire \DFF_11.CK ;
  wire \DFF_11.D ;
  wire \DFF_11.Q ;
  wire \DFF_110.CK ;
  wire \DFF_110.D ;
  wire \DFF_110.Q ;
  wire \DFF_111.CK ;
  wire \DFF_111.D ;
  wire \DFF_111.Q ;
  wire \DFF_112.CK ;
  wire \DFF_112.D ;
  wire \DFF_112.Q ;
  wire \DFF_113.CK ;
  wire \DFF_113.D ;
  wire \DFF_113.Q ;
  wire \DFF_114.CK ;
  wire \DFF_114.D ;
  wire \DFF_114.Q ;
  wire \DFF_115.CK ;
  wire \DFF_115.D ;
  wire \DFF_115.Q ;
  wire \DFF_116.CK ;
  wire \DFF_116.D ;
  wire \DFF_116.Q ;
  wire \DFF_117.CK ;
  wire \DFF_117.D ;
  wire \DFF_117.Q ;
  wire \DFF_118.CK ;
  wire \DFF_118.D ;
  wire \DFF_118.Q ;
  wire \DFF_119.CK ;
  wire \DFF_119.D ;
  wire \DFF_119.Q ;
  wire \DFF_12.CK ;
  wire \DFF_12.D ;
  wire \DFF_12.Q ;
  wire \DFF_120.CK ;
  wire \DFF_120.D ;
  wire \DFF_120.Q ;
  wire \DFF_121.CK ;
  wire \DFF_121.D ;
  wire \DFF_121.Q ;
  wire \DFF_122.CK ;
  wire \DFF_122.D ;
  wire \DFF_122.Q ;
  wire \DFF_123.CK ;
  wire \DFF_123.D ;
  wire \DFF_123.Q ;
  wire \DFF_124.CK ;
  wire \DFF_124.D ;
  wire \DFF_124.Q ;
  wire \DFF_125.CK ;
  wire \DFF_125.D ;
  wire \DFF_125.Q ;
  wire \DFF_126.CK ;
  wire \DFF_126.D ;
  wire \DFF_126.Q ;
  wire \DFF_127.CK ;
  wire \DFF_127.D ;
  wire \DFF_127.Q ;
  wire \DFF_128.CK ;
  wire \DFF_128.D ;
  wire \DFF_128.Q ;
  wire \DFF_129.CK ;
  wire \DFF_129.D ;
  wire \DFF_129.Q ;
  wire \DFF_13.CK ;
  wire \DFF_13.D ;
  wire \DFF_13.Q ;
  wire \DFF_130.CK ;
  wire \DFF_130.D ;
  wire \DFF_130.Q ;
  wire \DFF_131.CK ;
  wire \DFF_131.D ;
  wire \DFF_131.Q ;
  wire \DFF_132.CK ;
  wire \DFF_132.D ;
  wire \DFF_132.Q ;
  wire \DFF_133.CK ;
  wire \DFF_133.D ;
  wire \DFF_133.Q ;
  wire \DFF_134.CK ;
  wire \DFF_134.D ;
  wire \DFF_134.Q ;
  wire \DFF_135.CK ;
  wire \DFF_135.D ;
  wire \DFF_135.Q ;
  wire \DFF_136.CK ;
  wire \DFF_136.D ;
  wire \DFF_136.Q ;
  wire \DFF_137.CK ;
  wire \DFF_137.D ;
  wire \DFF_137.Q ;
  wire \DFF_138.CK ;
  wire \DFF_138.D ;
  wire \DFF_138.Q ;
  wire \DFF_139.CK ;
  wire \DFF_139.D ;
  wire \DFF_139.Q ;
  wire \DFF_14.CK ;
  wire \DFF_14.D ;
  wire \DFF_14.Q ;
  wire \DFF_140.CK ;
  wire \DFF_140.D ;
  wire \DFF_140.Q ;
  wire \DFF_141.CK ;
  wire \DFF_141.D ;
  wire \DFF_141.Q ;
  wire \DFF_142.CK ;
  wire \DFF_142.D ;
  wire \DFF_142.Q ;
  wire \DFF_143.CK ;
  wire \DFF_143.D ;
  wire \DFF_143.Q ;
  wire \DFF_144.CK ;
  wire \DFF_145.CK ;
  wire \DFF_145.D ;
  wire \DFF_145.Q ;
  wire \DFF_146.CK ;
  wire \DFF_146.D ;
  wire \DFF_146.Q ;
  wire \DFF_147.CK ;
  wire \DFF_147.D ;
  wire \DFF_147.Q ;
  wire \DFF_148.CK ;
  wire \DFF_148.D ;
  wire \DFF_148.Q ;
  wire \DFF_149.CK ;
  wire \DFF_149.D ;
  wire \DFF_149.Q ;
  wire \DFF_15.CK ;
  wire \DFF_15.D ;
  wire \DFF_15.Q ;
  wire \DFF_150.CK ;
  wire \DFF_150.D ;
  wire \DFF_150.Q ;
  wire \DFF_151.CK ;
  wire \DFF_151.D ;
  wire \DFF_151.Q ;
  wire \DFF_152.CK ;
  wire \DFF_152.D ;
  wire \DFF_152.Q ;
  wire \DFF_153.CK ;
  wire \DFF_153.D ;
  wire \DFF_153.Q ;
  wire \DFF_154.CK ;
  wire \DFF_154.D ;
  wire \DFF_154.Q ;
  wire \DFF_155.CK ;
  wire \DFF_155.D ;
  wire \DFF_155.Q ;
  wire \DFF_156.CK ;
  wire \DFF_156.D ;
  wire \DFF_156.Q ;
  wire \DFF_157.CK ;
  wire \DFF_157.D ;
  wire \DFF_157.Q ;
  wire \DFF_158.CK ;
  wire \DFF_158.D ;
  wire \DFF_158.Q ;
  wire \DFF_159.CK ;
  wire \DFF_159.D ;
  wire \DFF_159.Q ;
  wire \DFF_16.CK ;
  wire \DFF_16.D ;
  wire \DFF_16.Q ;
  wire \DFF_160.CK ;
  wire \DFF_160.D ;
  wire \DFF_160.Q ;
  wire \DFF_161.CK ;
  wire \DFF_161.D ;
  wire \DFF_161.Q ;
  wire \DFF_162.CK ;
  wire \DFF_162.D ;
  wire \DFF_162.Q ;
  wire \DFF_163.CK ;
  wire \DFF_163.D ;
  wire \DFF_163.Q ;
  wire \DFF_164.CK ;
  wire \DFF_164.D ;
  wire \DFF_164.Q ;
  wire \DFF_165.CK ;
  wire \DFF_165.D ;
  wire \DFF_165.Q ;
  wire \DFF_166.CK ;
  wire \DFF_166.D ;
  wire \DFF_166.Q ;
  wire \DFF_167.CK ;
  wire \DFF_167.D ;
  wire \DFF_167.Q ;
  wire \DFF_168.CK ;
  wire \DFF_168.D ;
  wire \DFF_168.Q ;
  wire \DFF_169.CK ;
  wire \DFF_169.D ;
  wire \DFF_169.Q ;
  wire \DFF_17.CK ;
  wire \DFF_17.D ;
  wire \DFF_17.Q ;
  wire \DFF_170.CK ;
  wire \DFF_170.D ;
  wire \DFF_170.Q ;
  wire \DFF_171.CK ;
  wire \DFF_171.D ;
  wire \DFF_171.Q ;
  wire \DFF_172.CK ;
  wire \DFF_172.D ;
  wire \DFF_172.Q ;
  wire \DFF_173.CK ;
  wire \DFF_173.D ;
  wire \DFF_173.Q ;
  wire \DFF_174.CK ;
  wire \DFF_174.D ;
  wire \DFF_174.Q ;
  wire \DFF_175.CK ;
  wire \DFF_175.D ;
  wire \DFF_175.Q ;
  wire \DFF_176.CK ;
  wire \DFF_176.D ;
  wire \DFF_176.Q ;
  wire \DFF_177.CK ;
  wire \DFF_177.D ;
  wire \DFF_177.Q ;
  wire \DFF_178.CK ;
  wire \DFF_178.D ;
  wire \DFF_178.Q ;
  wire \DFF_179.CK ;
  wire \DFF_179.D ;
  wire \DFF_179.Q ;
  wire \DFF_18.CK ;
  wire \DFF_18.D ;
  wire \DFF_18.Q ;
  wire \DFF_180.CK ;
  wire \DFF_180.D ;
  wire \DFF_180.Q ;
  wire \DFF_181.CK ;
  wire \DFF_181.D ;
  wire \DFF_181.Q ;
  wire \DFF_182.CK ;
  wire \DFF_182.D ;
  wire \DFF_182.Q ;
  wire \DFF_183.CK ;
  wire \DFF_183.D ;
  wire \DFF_183.Q ;
  wire \DFF_184.CK ;
  wire \DFF_184.D ;
  wire \DFF_184.Q ;
  wire \DFF_185.CK ;
  wire \DFF_185.D ;
  wire \DFF_185.Q ;
  wire \DFF_186.CK ;
  wire \DFF_186.D ;
  wire \DFF_186.Q ;
  wire \DFF_187.CK ;
  wire \DFF_187.D ;
  wire \DFF_187.Q ;
  wire \DFF_188.CK ;
  wire \DFF_188.D ;
  wire \DFF_188.Q ;
  wire \DFF_189.CK ;
  wire \DFF_189.D ;
  wire \DFF_189.Q ;
  wire \DFF_19.CK ;
  wire \DFF_19.D ;
  wire \DFF_19.Q ;
  wire \DFF_190.CK ;
  wire \DFF_190.D ;
  wire \DFF_190.Q ;
  wire \DFF_191.CK ;
  wire \DFF_191.D ;
  wire \DFF_191.Q ;
  wire \DFF_192.CK ;
  wire \DFF_192.D ;
  wire \DFF_192.Q ;
  wire \DFF_193.CK ;
  wire \DFF_193.D ;
  wire \DFF_193.Q ;
  wire \DFF_194.CK ;
  wire \DFF_194.D ;
  wire \DFF_194.Q ;
  wire \DFF_195.CK ;
  wire \DFF_195.D ;
  wire \DFF_195.Q ;
  wire \DFF_196.CK ;
  wire \DFF_196.D ;
  wire \DFF_196.Q ;
  wire \DFF_197.CK ;
  wire \DFF_197.D ;
  wire \DFF_197.Q ;
  wire \DFF_198.CK ;
  wire \DFF_198.D ;
  wire \DFF_198.Q ;
  wire \DFF_199.CK ;
  wire \DFF_199.D ;
  wire \DFF_199.Q ;
  wire \DFF_2.CK ;
  wire \DFF_2.D ;
  wire \DFF_2.Q ;
  wire \DFF_20.CK ;
  wire \DFF_20.D ;
  wire \DFF_20.Q ;
  wire \DFF_200.CK ;
  wire \DFF_200.D ;
  wire \DFF_200.Q ;
  wire \DFF_201.CK ;
  wire \DFF_201.D ;
  wire \DFF_201.Q ;
  wire \DFF_202.CK ;
  wire \DFF_202.D ;
  wire \DFF_202.Q ;
  wire \DFF_203.CK ;
  wire \DFF_203.D ;
  wire \DFF_203.Q ;
  wire \DFF_204.CK ;
  wire \DFF_204.D ;
  wire \DFF_204.Q ;
  wire \DFF_205.CK ;
  wire \DFF_205.D ;
  wire \DFF_205.Q ;
  wire \DFF_206.CK ;
  wire \DFF_206.D ;
  wire \DFF_206.Q ;
  wire \DFF_207.CK ;
  wire \DFF_207.D ;
  wire \DFF_207.Q ;
  wire \DFF_208.CK ;
  wire \DFF_208.D ;
  wire \DFF_208.Q ;
  wire \DFF_209.CK ;
  wire \DFF_209.D ;
  wire \DFF_209.Q ;
  wire \DFF_21.CK ;
  wire \DFF_21.D ;
  wire \DFF_21.Q ;
  wire \DFF_210.CK ;
  wire \DFF_210.D ;
  wire \DFF_210.Q ;
  wire \DFF_211.CK ;
  wire \DFF_211.D ;
  wire \DFF_211.Q ;
  wire \DFF_212.CK ;
  wire \DFF_212.D ;
  wire \DFF_212.Q ;
  wire \DFF_213.CK ;
  wire \DFF_213.D ;
  wire \DFF_213.Q ;
  wire \DFF_214.CK ;
  wire \DFF_214.D ;
  wire \DFF_214.Q ;
  wire \DFF_215.CK ;
  wire \DFF_215.D ;
  wire \DFF_215.Q ;
  wire \DFF_216.CK ;
  wire \DFF_216.D ;
  wire \DFF_216.Q ;
  wire \DFF_217.CK ;
  wire \DFF_217.D ;
  wire \DFF_217.Q ;
  wire \DFF_218.CK ;
  wire \DFF_218.D ;
  wire \DFF_218.Q ;
  wire \DFF_219.CK ;
  wire \DFF_22.CK ;
  wire \DFF_22.D ;
  wire \DFF_22.Q ;
  wire \DFF_220.CK ;
  wire \DFF_220.D ;
  wire \DFF_220.Q ;
  wire \DFF_221.CK ;
  wire \DFF_221.D ;
  wire \DFF_221.Q ;
  wire \DFF_222.CK ;
  wire \DFF_222.D ;
  wire \DFF_222.Q ;
  wire \DFF_223.CK ;
  wire \DFF_223.D ;
  wire \DFF_223.Q ;
  wire \DFF_224.CK ;
  wire \DFF_224.D ;
  wire \DFF_224.Q ;
  wire \DFF_225.CK ;
  wire \DFF_225.D ;
  wire \DFF_225.Q ;
  wire \DFF_226.CK ;
  wire \DFF_226.D ;
  wire \DFF_226.Q ;
  wire \DFF_227.CK ;
  wire \DFF_227.D ;
  wire \DFF_227.Q ;
  wire \DFF_228.CK ;
  wire \DFF_228.D ;
  wire \DFF_228.Q ;
  wire \DFF_229.CK ;
  wire \DFF_229.D ;
  wire \DFF_229.Q ;
  wire \DFF_23.CK ;
  wire \DFF_23.D ;
  wire \DFF_23.Q ;
  wire \DFF_230.CK ;
  wire \DFF_230.D ;
  wire \DFF_230.Q ;
  wire \DFF_231.CK ;
  wire \DFF_231.D ;
  wire \DFF_231.Q ;
  wire \DFF_232.CK ;
  wire \DFF_232.D ;
  wire \DFF_232.Q ;
  wire \DFF_233.CK ;
  wire \DFF_233.D ;
  wire \DFF_233.Q ;
  wire \DFF_234.CK ;
  wire \DFF_234.D ;
  wire \DFF_234.Q ;
  wire \DFF_235.CK ;
  wire \DFF_235.D ;
  wire \DFF_235.Q ;
  wire \DFF_236.CK ;
  wire \DFF_236.D ;
  wire \DFF_236.Q ;
  wire \DFF_237.CK ;
  wire \DFF_237.D ;
  wire \DFF_237.Q ;
  wire \DFF_238.CK ;
  wire \DFF_238.D ;
  wire \DFF_238.Q ;
  wire \DFF_239.CK ;
  wire \DFF_239.D ;
  wire \DFF_239.Q ;
  wire \DFF_24.CK ;
  wire \DFF_24.D ;
  wire \DFF_24.Q ;
  wire \DFF_240.CK ;
  wire \DFF_240.D ;
  wire \DFF_240.Q ;
  wire \DFF_241.CK ;
  wire \DFF_241.D ;
  wire \DFF_241.Q ;
  wire \DFF_242.CK ;
  wire \DFF_242.D ;
  wire \DFF_242.Q ;
  wire \DFF_243.CK ;
  wire \DFF_243.D ;
  wire \DFF_243.Q ;
  wire \DFF_244.CK ;
  wire \DFF_244.D ;
  wire \DFF_244.Q ;
  wire \DFF_245.CK ;
  wire \DFF_245.D ;
  wire \DFF_245.Q ;
  wire \DFF_246.CK ;
  wire \DFF_246.D ;
  wire \DFF_246.Q ;
  wire \DFF_247.CK ;
  wire \DFF_247.D ;
  wire \DFF_247.Q ;
  wire \DFF_248.CK ;
  wire \DFF_248.D ;
  wire \DFF_248.Q ;
  wire \DFF_249.CK ;
  wire \DFF_249.D ;
  wire \DFF_249.Q ;
  wire \DFF_25.CK ;
  wire \DFF_25.D ;
  wire \DFF_25.Q ;
  wire \DFF_250.CK ;
  wire \DFF_250.D ;
  wire \DFF_250.Q ;
  wire \DFF_251.CK ;
  wire \DFF_251.D ;
  wire \DFF_251.Q ;
  wire \DFF_252.CK ;
  wire \DFF_252.D ;
  wire \DFF_252.Q ;
  wire \DFF_253.CK ;
  wire \DFF_253.D ;
  wire \DFF_253.Q ;
  wire \DFF_254.CK ;
  wire \DFF_254.D ;
  wire \DFF_254.Q ;
  wire \DFF_255.CK ;
  wire \DFF_255.D ;
  wire \DFF_255.Q ;
  wire \DFF_256.CK ;
  wire \DFF_256.D ;
  wire \DFF_256.Q ;
  wire \DFF_257.CK ;
  wire \DFF_258.CK ;
  wire \DFF_258.D ;
  wire \DFF_258.Q ;
  wire \DFF_259.CK ;
  wire \DFF_259.D ;
  wire \DFF_259.Q ;
  wire \DFF_26.CK ;
  wire \DFF_26.D ;
  wire \DFF_26.Q ;
  wire \DFF_260.CK ;
  wire \DFF_260.D ;
  wire \DFF_260.Q ;
  wire \DFF_261.CK ;
  wire \DFF_261.D ;
  wire \DFF_261.Q ;
  wire \DFF_262.CK ;
  wire \DFF_262.D ;
  wire \DFF_262.Q ;
  wire \DFF_263.CK ;
  wire \DFF_263.D ;
  wire \DFF_263.Q ;
  wire \DFF_264.CK ;
  wire \DFF_264.D ;
  wire \DFF_264.Q ;
  wire \DFF_265.CK ;
  wire \DFF_265.D ;
  wire \DFF_265.Q ;
  wire \DFF_266.CK ;
  wire \DFF_266.D ;
  wire \DFF_266.Q ;
  wire \DFF_267.CK ;
  wire \DFF_267.D ;
  wire \DFF_267.Q ;
  wire \DFF_268.CK ;
  wire \DFF_268.D ;
  wire \DFF_268.Q ;
  wire \DFF_269.CK ;
  wire \DFF_269.D ;
  wire \DFF_269.Q ;
  wire \DFF_27.CK ;
  wire \DFF_27.D ;
  wire \DFF_27.Q ;
  wire \DFF_270.CK ;
  wire \DFF_270.D ;
  wire \DFF_270.Q ;
  wire \DFF_271.CK ;
  wire \DFF_271.D ;
  wire \DFF_271.Q ;
  wire \DFF_272.CK ;
  wire \DFF_272.D ;
  wire \DFF_272.Q ;
  wire \DFF_273.CK ;
  wire \DFF_273.D ;
  wire \DFF_273.Q ;
  wire \DFF_274.CK ;
  wire \DFF_274.D ;
  wire \DFF_274.Q ;
  wire \DFF_275.CK ;
  wire \DFF_275.D ;
  wire \DFF_275.Q ;
  wire \DFF_276.CK ;
  wire \DFF_276.D ;
  wire \DFF_276.Q ;
  wire \DFF_277.CK ;
  wire \DFF_277.D ;
  wire \DFF_277.Q ;
  wire \DFF_278.CK ;
  wire \DFF_278.D ;
  wire \DFF_278.Q ;
  wire \DFF_279.CK ;
  wire \DFF_279.D ;
  wire \DFF_279.Q ;
  wire \DFF_28.CK ;
  wire \DFF_28.D ;
  wire \DFF_28.Q ;
  wire \DFF_280.CK ;
  wire \DFF_280.D ;
  wire \DFF_280.Q ;
  wire \DFF_281.CK ;
  wire \DFF_281.D ;
  wire \DFF_281.Q ;
  wire \DFF_282.CK ;
  wire \DFF_282.D ;
  wire \DFF_282.Q ;
  wire \DFF_283.CK ;
  wire \DFF_283.D ;
  wire \DFF_283.Q ;
  wire \DFF_284.CK ;
  wire \DFF_284.D ;
  wire \DFF_284.Q ;
  wire \DFF_285.CK ;
  wire \DFF_285.D ;
  wire \DFF_285.Q ;
  wire \DFF_286.CK ;
  wire \DFF_286.D ;
  wire \DFF_286.Q ;
  wire \DFF_287.CK ;
  wire \DFF_287.D ;
  wire \DFF_287.Q ;
  wire \DFF_288.CK ;
  wire \DFF_288.D ;
  wire \DFF_288.Q ;
  wire \DFF_289.CK ;
  wire \DFF_289.D ;
  wire \DFF_289.Q ;
  wire \DFF_29.CK ;
  wire \DFF_29.D ;
  wire \DFF_29.Q ;
  wire \DFF_290.CK ;
  wire \DFF_290.D ;
  wire \DFF_290.Q ;
  wire \DFF_291.CK ;
  wire \DFF_291.D ;
  wire \DFF_291.Q ;
  wire \DFF_292.CK ;
  wire \DFF_292.D ;
  wire \DFF_292.Q ;
  wire \DFF_293.CK ;
  wire \DFF_293.D ;
  wire \DFF_293.Q ;
  wire \DFF_294.CK ;
  wire \DFF_294.D ;
  wire \DFF_294.Q ;
  wire \DFF_295.CK ;
  wire \DFF_295.D ;
  wire \DFF_295.Q ;
  wire \DFF_296.CK ;
  wire \DFF_296.D ;
  wire \DFF_296.Q ;
  wire \DFF_297.CK ;
  wire \DFF_297.D ;
  wire \DFF_297.Q ;
  wire \DFF_298.CK ;
  wire \DFF_298.D ;
  wire \DFF_298.Q ;
  wire \DFF_299.CK ;
  wire \DFF_299.D ;
  wire \DFF_299.Q ;
  wire \DFF_3.CK ;
  wire \DFF_3.D ;
  wire \DFF_3.Q ;
  wire \DFF_30.CK ;
  wire \DFF_30.D ;
  wire \DFF_30.Q ;
  wire \DFF_300.CK ;
  wire \DFF_300.D ;
  wire \DFF_300.Q ;
  wire \DFF_301.CK ;
  wire \DFF_301.D ;
  wire \DFF_301.Q ;
  wire \DFF_302.CK ;
  wire \DFF_302.D ;
  wire \DFF_302.Q ;
  wire \DFF_303.CK ;
  wire \DFF_303.D ;
  wire \DFF_303.Q ;
  wire \DFF_304.CK ;
  wire \DFF_304.D ;
  wire \DFF_304.Q ;
  wire \DFF_305.CK ;
  wire \DFF_305.D ;
  wire \DFF_305.Q ;
  wire \DFF_306.CK ;
  wire \DFF_306.D ;
  wire \DFF_306.Q ;
  wire \DFF_307.CK ;
  wire \DFF_307.D ;
  wire \DFF_307.Q ;
  wire \DFF_308.CK ;
  wire \DFF_308.D ;
  wire \DFF_308.Q ;
  wire \DFF_309.CK ;
  wire \DFF_309.D ;
  wire \DFF_309.Q ;
  wire \DFF_31.CK ;
  wire \DFF_31.D ;
  wire \DFF_31.Q ;
  wire \DFF_310.CK ;
  wire \DFF_310.D ;
  wire \DFF_310.Q ;
  wire \DFF_311.CK ;
  wire \DFF_311.D ;
  wire \DFF_311.Q ;
  wire \DFF_312.CK ;
  wire \DFF_312.D ;
  wire \DFF_312.Q ;
  wire \DFF_313.CK ;
  wire \DFF_313.D ;
  wire \DFF_313.Q ;
  wire \DFF_314.CK ;
  wire \DFF_314.D ;
  wire \DFF_314.Q ;
  wire \DFF_315.CK ;
  wire \DFF_315.D ;
  wire \DFF_315.Q ;
  wire \DFF_316.CK ;
  wire \DFF_316.D ;
  wire \DFF_316.Q ;
  wire \DFF_317.CK ;
  wire \DFF_317.D ;
  wire \DFF_317.Q ;
  wire \DFF_318.CK ;
  wire \DFF_318.D ;
  wire \DFF_318.Q ;
  wire \DFF_319.CK ;
  wire \DFF_319.D ;
  wire \DFF_319.Q ;
  wire \DFF_32.CK ;
  wire \DFF_32.D ;
  wire \DFF_32.Q ;
  wire \DFF_320.CK ;
  wire \DFF_320.D ;
  wire \DFF_320.Q ;
  wire \DFF_321.CK ;
  wire \DFF_321.D ;
  wire \DFF_321.Q ;
  wire \DFF_322.CK ;
  wire \DFF_322.D ;
  wire \DFF_322.Q ;
  wire \DFF_323.CK ;
  wire \DFF_323.D ;
  wire \DFF_323.Q ;
  wire \DFF_324.CK ;
  wire \DFF_324.D ;
  wire \DFF_324.Q ;
  wire \DFF_325.CK ;
  wire \DFF_325.D ;
  wire \DFF_325.Q ;
  wire \DFF_326.CK ;
  wire \DFF_326.D ;
  wire \DFF_326.Q ;
  wire \DFF_327.CK ;
  wire \DFF_327.D ;
  wire \DFF_327.Q ;
  wire \DFF_328.CK ;
  wire \DFF_328.D ;
  wire \DFF_328.Q ;
  wire \DFF_329.CK ;
  wire \DFF_329.D ;
  wire \DFF_329.Q ;
  wire \DFF_33.CK ;
  wire \DFF_33.D ;
  wire \DFF_33.Q ;
  wire \DFF_330.CK ;
  wire \DFF_330.D ;
  wire \DFF_330.Q ;
  wire \DFF_331.CK ;
  wire \DFF_331.D ;
  wire \DFF_331.Q ;
  wire \DFF_332.CK ;
  wire \DFF_332.D ;
  wire \DFF_332.Q ;
  wire \DFF_333.CK ;
  wire \DFF_333.D ;
  wire \DFF_333.Q ;
  wire \DFF_334.CK ;
  wire \DFF_334.D ;
  wire \DFF_334.Q ;
  wire \DFF_335.CK ;
  wire \DFF_335.D ;
  wire \DFF_335.Q ;
  wire \DFF_336.CK ;
  wire \DFF_336.D ;
  wire \DFF_336.Q ;
  wire \DFF_337.CK ;
  wire \DFF_337.D ;
  wire \DFF_337.Q ;
  wire \DFF_338.CK ;
  wire \DFF_338.D ;
  wire \DFF_338.Q ;
  wire \DFF_339.CK ;
  wire \DFF_339.D ;
  wire \DFF_339.Q ;
  wire \DFF_34.CK ;
  wire \DFF_34.D ;
  wire \DFF_34.Q ;
  wire \DFF_340.CK ;
  wire \DFF_340.D ;
  wire \DFF_340.Q ;
  wire \DFF_341.CK ;
  wire \DFF_342.CK ;
  wire \DFF_342.D ;
  wire \DFF_342.Q ;
  wire \DFF_343.CK ;
  wire \DFF_343.D ;
  wire \DFF_343.Q ;
  wire \DFF_344.CK ;
  wire \DFF_344.D ;
  wire \DFF_344.Q ;
  wire \DFF_345.CK ;
  wire \DFF_345.D ;
  wire \DFF_345.Q ;
  wire \DFF_346.CK ;
  wire \DFF_346.D ;
  wire \DFF_346.Q ;
  wire \DFF_347.CK ;
  wire \DFF_347.D ;
  wire \DFF_347.Q ;
  wire \DFF_348.CK ;
  wire \DFF_348.D ;
  wire \DFF_348.Q ;
  wire \DFF_349.CK ;
  wire \DFF_349.D ;
  wire \DFF_349.Q ;
  wire \DFF_35.CK ;
  wire \DFF_35.D ;
  wire \DFF_35.Q ;
  wire \DFF_350.CK ;
  wire \DFF_350.D ;
  wire \DFF_350.Q ;
  wire \DFF_351.CK ;
  wire \DFF_351.D ;
  wire \DFF_351.Q ;
  wire \DFF_352.CK ;
  wire \DFF_352.D ;
  wire \DFF_352.Q ;
  wire \DFF_353.CK ;
  wire \DFF_353.D ;
  wire \DFF_353.Q ;
  wire \DFF_354.CK ;
  wire \DFF_354.D ;
  wire \DFF_354.Q ;
  wire \DFF_355.CK ;
  wire \DFF_355.D ;
  wire \DFF_355.Q ;
  wire \DFF_356.CK ;
  wire \DFF_356.D ;
  wire \DFF_356.Q ;
  wire \DFF_357.CK ;
  wire \DFF_357.D ;
  wire \DFF_357.Q ;
  wire \DFF_358.CK ;
  wire \DFF_358.D ;
  wire \DFF_358.Q ;
  wire \DFF_359.CK ;
  wire \DFF_359.D ;
  wire \DFF_359.Q ;
  wire \DFF_36.CK ;
  wire \DFF_36.D ;
  wire \DFF_36.Q ;
  wire \DFF_360.CK ;
  wire \DFF_360.D ;
  wire \DFF_360.Q ;
  wire \DFF_361.CK ;
  wire \DFF_361.D ;
  wire \DFF_361.Q ;
  wire \DFF_362.CK ;
  wire \DFF_362.D ;
  wire \DFF_362.Q ;
  wire \DFF_363.CK ;
  wire \DFF_363.D ;
  wire \DFF_363.Q ;
  wire \DFF_364.CK ;
  wire \DFF_364.D ;
  wire \DFF_364.Q ;
  wire \DFF_365.CK ;
  wire \DFF_365.D ;
  wire \DFF_365.Q ;
  wire \DFF_366.CK ;
  wire \DFF_366.D ;
  wire \DFF_366.Q ;
  wire \DFF_367.CK ;
  wire \DFF_367.D ;
  wire \DFF_367.Q ;
  wire \DFF_368.CK ;
  wire \DFF_368.D ;
  wire \DFF_368.Q ;
  wire \DFF_369.CK ;
  wire \DFF_369.D ;
  wire \DFF_369.Q ;
  wire \DFF_37.CK ;
  wire \DFF_37.D ;
  wire \DFF_37.Q ;
  wire \DFF_370.CK ;
  wire \DFF_370.D ;
  wire \DFF_370.Q ;
  wire \DFF_371.CK ;
  wire \DFF_371.D ;
  wire \DFF_371.Q ;
  wire \DFF_372.CK ;
  wire \DFF_372.D ;
  wire \DFF_372.Q ;
  wire \DFF_373.CK ;
  wire \DFF_373.D ;
  wire \DFF_373.Q ;
  wire \DFF_374.CK ;
  wire \DFF_374.D ;
  wire \DFF_374.Q ;
  wire \DFF_375.CK ;
  wire \DFF_376.CK ;
  wire \DFF_376.D ;
  wire \DFF_376.Q ;
  wire \DFF_377.CK ;
  wire \DFF_377.D ;
  wire \DFF_377.Q ;
  wire \DFF_378.CK ;
  wire \DFF_378.D ;
  wire \DFF_378.Q ;
  wire \DFF_379.CK ;
  wire \DFF_379.D ;
  wire \DFF_379.Q ;
  wire \DFF_38.CK ;
  wire \DFF_38.D ;
  wire \DFF_38.Q ;
  wire \DFF_380.CK ;
  wire \DFF_380.D ;
  wire \DFF_380.Q ;
  wire \DFF_381.CK ;
  wire \DFF_381.D ;
  wire \DFF_381.Q ;
  wire \DFF_382.CK ;
  wire \DFF_382.D ;
  wire \DFF_382.Q ;
  wire \DFF_383.CK ;
  wire \DFF_383.D ;
  wire \DFF_383.Q ;
  wire \DFF_384.CK ;
  wire \DFF_384.D ;
  wire \DFF_384.Q ;
  wire \DFF_385.CK ;
  wire \DFF_385.D ;
  wire \DFF_385.Q ;
  wire \DFF_386.CK ;
  wire \DFF_386.D ;
  wire \DFF_386.Q ;
  wire \DFF_387.CK ;
  wire \DFF_387.D ;
  wire \DFF_387.Q ;
  wire \DFF_388.CK ;
  wire \DFF_388.D ;
  wire \DFF_388.Q ;
  wire \DFF_389.CK ;
  wire \DFF_389.D ;
  wire \DFF_389.Q ;
  wire \DFF_39.CK ;
  wire \DFF_39.D ;
  wire \DFF_39.Q ;
  wire \DFF_390.CK ;
  wire \DFF_390.D ;
  wire \DFF_390.Q ;
  wire \DFF_391.CK ;
  wire \DFF_391.D ;
  wire \DFF_391.Q ;
  wire \DFF_392.CK ;
  wire \DFF_392.D ;
  wire \DFF_392.Q ;
  wire \DFF_393.CK ;
  wire \DFF_393.D ;
  wire \DFF_393.Q ;
  wire \DFF_394.CK ;
  wire \DFF_394.D ;
  wire \DFF_394.Q ;
  wire \DFF_395.CK ;
  wire \DFF_395.D ;
  wire \DFF_395.Q ;
  wire \DFF_396.CK ;
  wire \DFF_396.D ;
  wire \DFF_396.Q ;
  wire \DFF_397.CK ;
  wire \DFF_397.D ;
  wire \DFF_397.Q ;
  wire \DFF_398.CK ;
  wire \DFF_398.D ;
  wire \DFF_398.Q ;
  wire \DFF_399.CK ;
  wire \DFF_399.D ;
  wire \DFF_399.Q ;
  wire \DFF_4.CK ;
  wire \DFF_4.D ;
  wire \DFF_4.Q ;
  wire \DFF_40.CK ;
  wire \DFF_400.CK ;
  wire \DFF_400.D ;
  wire \DFF_400.Q ;
  wire \DFF_401.CK ;
  wire \DFF_401.D ;
  wire \DFF_401.Q ;
  wire \DFF_402.CK ;
  wire \DFF_402.D ;
  wire \DFF_402.Q ;
  wire \DFF_403.CK ;
  wire \DFF_403.D ;
  wire \DFF_403.Q ;
  wire \DFF_404.CK ;
  wire \DFF_404.D ;
  wire \DFF_404.Q ;
  wire \DFF_405.CK ;
  wire \DFF_405.D ;
  wire \DFF_405.Q ;
  wire \DFF_406.CK ;
  wire \DFF_406.D ;
  wire \DFF_406.Q ;
  wire \DFF_407.CK ;
  wire \DFF_407.D ;
  wire \DFF_407.Q ;
  wire \DFF_408.CK ;
  wire \DFF_408.D ;
  wire \DFF_408.Q ;
  wire \DFF_409.CK ;
  wire \DFF_409.D ;
  wire \DFF_409.Q ;
  wire \DFF_41.CK ;
  wire \DFF_41.D ;
  wire \DFF_41.Q ;
  wire \DFF_410.CK ;
  wire \DFF_410.D ;
  wire \DFF_410.Q ;
  wire \DFF_411.CK ;
  wire \DFF_411.D ;
  wire \DFF_411.Q ;
  wire \DFF_412.CK ;
  wire \DFF_412.D ;
  wire \DFF_412.Q ;
  wire \DFF_413.CK ;
  wire \DFF_413.D ;
  wire \DFF_413.Q ;
  wire \DFF_414.CK ;
  wire \DFF_414.D ;
  wire \DFF_414.Q ;
  wire \DFF_415.CK ;
  wire \DFF_415.D ;
  wire \DFF_415.Q ;
  wire \DFF_416.CK ;
  wire \DFF_416.D ;
  wire \DFF_416.Q ;
  wire \DFF_417.CK ;
  wire \DFF_417.D ;
  wire \DFF_417.Q ;
  wire \DFF_418.CK ;
  wire \DFF_418.D ;
  wire \DFF_418.Q ;
  wire \DFF_419.CK ;
  wire \DFF_419.D ;
  wire \DFF_419.Q ;
  wire \DFF_42.CK ;
  wire \DFF_42.D ;
  wire \DFF_42.Q ;
  wire \DFF_420.CK ;
  wire \DFF_420.D ;
  wire \DFF_420.Q ;
  wire \DFF_421.CK ;
  wire \DFF_421.D ;
  wire \DFF_421.Q ;
  wire \DFF_422.CK ;
  wire \DFF_422.D ;
  wire \DFF_422.Q ;
  wire \DFF_423.CK ;
  wire \DFF_423.D ;
  wire \DFF_423.Q ;
  wire \DFF_424.CK ;
  wire \DFF_424.D ;
  wire \DFF_424.Q ;
  wire \DFF_425.CK ;
  wire \DFF_425.D ;
  wire \DFF_425.Q ;
  wire \DFF_426.CK ;
  wire \DFF_426.D ;
  wire \DFF_426.Q ;
  wire \DFF_427.CK ;
  wire \DFF_427.D ;
  wire \DFF_427.Q ;
  wire \DFF_428.CK ;
  wire \DFF_428.D ;
  wire \DFF_428.Q ;
  wire \DFF_429.CK ;
  wire \DFF_429.D ;
  wire \DFF_429.Q ;
  wire \DFF_43.CK ;
  wire \DFF_43.D ;
  wire \DFF_43.Q ;
  wire \DFF_430.CK ;
  wire \DFF_430.D ;
  wire \DFF_430.Q ;
  wire \DFF_431.CK ;
  wire \DFF_431.D ;
  wire \DFF_431.Q ;
  wire \DFF_432.CK ;
  wire \DFF_432.D ;
  wire \DFF_432.Q ;
  wire \DFF_433.CK ;
  wire \DFF_433.D ;
  wire \DFF_433.Q ;
  wire \DFF_434.CK ;
  wire \DFF_434.D ;
  wire \DFF_434.Q ;
  wire \DFF_435.CK ;
  wire \DFF_435.D ;
  wire \DFF_435.Q ;
  wire \DFF_436.CK ;
  wire \DFF_436.D ;
  wire \DFF_436.Q ;
  wire \DFF_437.CK ;
  wire \DFF_437.D ;
  wire \DFF_437.Q ;
  wire \DFF_438.CK ;
  wire \DFF_438.D ;
  wire \DFF_438.Q ;
  wire \DFF_439.CK ;
  wire \DFF_439.D ;
  wire \DFF_439.Q ;
  wire \DFF_44.CK ;
  wire \DFF_44.D ;
  wire \DFF_44.Q ;
  wire \DFF_440.CK ;
  wire \DFF_440.D ;
  wire \DFF_440.Q ;
  wire \DFF_441.CK ;
  wire \DFF_441.D ;
  wire \DFF_441.Q ;
  wire \DFF_442.CK ;
  wire \DFF_442.D ;
  wire \DFF_442.Q ;
  wire \DFF_443.CK ;
  wire \DFF_443.D ;
  wire \DFF_443.Q ;
  wire \DFF_444.CK ;
  wire \DFF_444.D ;
  wire \DFF_444.Q ;
  wire \DFF_445.CK ;
  wire \DFF_445.D ;
  wire \DFF_445.Q ;
  wire \DFF_446.CK ;
  wire \DFF_446.D ;
  wire \DFF_446.Q ;
  wire \DFF_447.CK ;
  wire \DFF_447.D ;
  wire \DFF_447.Q ;
  wire \DFF_448.CK ;
  wire \DFF_448.D ;
  wire \DFF_448.Q ;
  wire \DFF_449.CK ;
  wire \DFF_449.D ;
  wire \DFF_449.Q ;
  wire \DFF_45.CK ;
  wire \DFF_45.D ;
  wire \DFF_45.Q ;
  wire \DFF_450.CK ;
  wire \DFF_450.D ;
  wire \DFF_450.Q ;
  wire \DFF_451.CK ;
  wire \DFF_451.D ;
  wire \DFF_451.Q ;
  wire \DFF_452.CK ;
  wire \DFF_452.D ;
  wire \DFF_452.Q ;
  wire \DFF_453.CK ;
  wire \DFF_453.D ;
  wire \DFF_453.Q ;
  wire \DFF_454.CK ;
  wire \DFF_454.D ;
  wire \DFF_454.Q ;
  wire \DFF_455.CK ;
  wire \DFF_455.D ;
  wire \DFF_455.Q ;
  wire \DFF_456.CK ;
  wire \DFF_456.D ;
  wire \DFF_456.Q ;
  wire \DFF_457.CK ;
  wire \DFF_457.D ;
  wire \DFF_457.Q ;
  wire \DFF_458.CK ;
  wire \DFF_458.D ;
  wire \DFF_458.Q ;
  wire \DFF_459.CK ;
  wire \DFF_459.D ;
  wire \DFF_459.Q ;
  wire \DFF_46.CK ;
  wire \DFF_46.D ;
  wire \DFF_46.Q ;
  wire \DFF_460.CK ;
  wire \DFF_460.D ;
  wire \DFF_460.Q ;
  wire \DFF_461.CK ;
  wire \DFF_461.D ;
  wire \DFF_461.Q ;
  wire \DFF_462.CK ;
  wire \DFF_462.D ;
  wire \DFF_462.Q ;
  wire \DFF_463.CK ;
  wire \DFF_463.D ;
  wire \DFF_463.Q ;
  wire \DFF_464.CK ;
  wire \DFF_464.D ;
  wire \DFF_464.Q ;
  wire \DFF_465.CK ;
  wire \DFF_465.D ;
  wire \DFF_465.Q ;
  wire \DFF_466.CK ;
  wire \DFF_466.D ;
  wire \DFF_466.Q ;
  wire \DFF_467.CK ;
  wire \DFF_467.D ;
  wire \DFF_467.Q ;
  wire \DFF_468.CK ;
  wire \DFF_468.D ;
  wire \DFF_468.Q ;
  wire \DFF_469.CK ;
  wire \DFF_47.CK ;
  wire \DFF_47.D ;
  wire \DFF_47.Q ;
  wire \DFF_470.CK ;
  wire \DFF_470.D ;
  wire \DFF_470.Q ;
  wire \DFF_471.CK ;
  wire \DFF_471.D ;
  wire \DFF_471.Q ;
  wire \DFF_472.CK ;
  wire \DFF_472.D ;
  wire \DFF_472.Q ;
  wire \DFF_473.CK ;
  wire \DFF_473.D ;
  wire \DFF_473.Q ;
  wire \DFF_474.CK ;
  wire \DFF_474.D ;
  wire \DFF_474.Q ;
  wire \DFF_475.CK ;
  wire \DFF_475.D ;
  wire \DFF_475.Q ;
  wire \DFF_476.CK ;
  wire \DFF_476.D ;
  wire \DFF_476.Q ;
  wire \DFF_477.CK ;
  wire \DFF_477.D ;
  wire \DFF_477.Q ;
  wire \DFF_478.CK ;
  wire \DFF_478.D ;
  wire \DFF_478.Q ;
  wire \DFF_479.CK ;
  wire \DFF_479.D ;
  wire \DFF_479.Q ;
  wire \DFF_48.CK ;
  wire \DFF_48.D ;
  wire \DFF_48.Q ;
  wire \DFF_480.CK ;
  wire \DFF_480.D ;
  wire \DFF_480.Q ;
  wire \DFF_481.CK ;
  wire \DFF_481.D ;
  wire \DFF_481.Q ;
  wire \DFF_482.CK ;
  wire \DFF_482.D ;
  wire \DFF_482.Q ;
  wire \DFF_483.CK ;
  wire \DFF_483.D ;
  wire \DFF_483.Q ;
  wire \DFF_484.CK ;
  wire \DFF_484.D ;
  wire \DFF_484.Q ;
  wire \DFF_485.CK ;
  wire \DFF_485.D ;
  wire \DFF_485.Q ;
  wire \DFF_486.CK ;
  wire \DFF_486.D ;
  wire \DFF_486.Q ;
  wire \DFF_487.CK ;
  wire \DFF_487.D ;
  wire \DFF_487.Q ;
  wire \DFF_488.CK ;
  wire \DFF_488.D ;
  wire \DFF_488.Q ;
  wire \DFF_489.CK ;
  wire \DFF_489.D ;
  wire \DFF_489.Q ;
  wire \DFF_49.CK ;
  wire \DFF_49.D ;
  wire \DFF_49.Q ;
  wire \DFF_490.CK ;
  wire \DFF_490.D ;
  wire \DFF_490.Q ;
  wire \DFF_491.CK ;
  wire \DFF_491.D ;
  wire \DFF_491.Q ;
  wire \DFF_492.CK ;
  wire \DFF_492.D ;
  wire \DFF_492.Q ;
  wire \DFF_493.CK ;
  wire \DFF_493.D ;
  wire \DFF_493.Q ;
  wire \DFF_494.CK ;
  wire \DFF_494.D ;
  wire \DFF_494.Q ;
  wire \DFF_495.CK ;
  wire \DFF_495.D ;
  wire \DFF_495.Q ;
  wire \DFF_496.CK ;
  wire \DFF_496.D ;
  wire \DFF_496.Q ;
  wire \DFF_497.CK ;
  wire \DFF_497.D ;
  wire \DFF_497.Q ;
  wire \DFF_498.CK ;
  wire \DFF_498.D ;
  wire \DFF_498.Q ;
  wire \DFF_499.CK ;
  wire \DFF_499.D ;
  wire \DFF_499.Q ;
  wire \DFF_5.CK ;
  wire \DFF_5.D ;
  wire \DFF_5.Q ;
  wire \DFF_50.CK ;
  wire \DFF_50.D ;
  wire \DFF_50.Q ;
  wire \DFF_500.CK ;
  wire \DFF_500.D ;
  wire \DFF_500.Q ;
  wire \DFF_501.CK ;
  wire \DFF_501.D ;
  wire \DFF_501.Q ;
  wire \DFF_502.CK ;
  wire \DFF_502.D ;
  wire \DFF_502.Q ;
  wire \DFF_503.CK ;
  wire \DFF_503.D ;
  wire \DFF_503.Q ;
  wire \DFF_504.CK ;
  wire \DFF_504.D ;
  wire \DFF_504.Q ;
  wire \DFF_505.CK ;
  wire \DFF_505.D ;
  wire \DFF_505.Q ;
  wire \DFF_506.CK ;
  wire \DFF_506.D ;
  wire \DFF_506.Q ;
  wire \DFF_507.CK ;
  wire \DFF_507.D ;
  wire \DFF_507.Q ;
  wire \DFF_508.CK ;
  wire \DFF_508.D ;
  wire \DFF_508.Q ;
  wire \DFF_509.CK ;
  wire \DFF_509.D ;
  wire \DFF_509.Q ;
  wire \DFF_51.CK ;
  wire \DFF_51.D ;
  wire \DFF_51.Q ;
  wire \DFF_510.CK ;
  wire \DFF_510.D ;
  wire \DFF_510.Q ;
  wire \DFF_511.CK ;
  wire \DFF_511.D ;
  wire \DFF_511.Q ;
  wire \DFF_512.CK ;
  wire \DFF_512.D ;
  wire \DFF_512.Q ;
  wire \DFF_513.CK ;
  wire \DFF_513.D ;
  wire \DFF_513.Q ;
  wire \DFF_514.CK ;
  wire \DFF_514.D ;
  wire \DFF_514.Q ;
  wire \DFF_515.CK ;
  wire \DFF_515.D ;
  wire \DFF_515.Q ;
  wire \DFF_516.CK ;
  wire \DFF_516.D ;
  wire \DFF_516.Q ;
  wire \DFF_517.CK ;
  wire \DFF_517.D ;
  wire \DFF_517.Q ;
  wire \DFF_518.CK ;
  wire \DFF_518.D ;
  wire \DFF_518.Q ;
  wire \DFF_519.CK ;
  wire \DFF_519.D ;
  wire \DFF_519.Q ;
  wire \DFF_52.CK ;
  wire \DFF_52.D ;
  wire \DFF_52.Q ;
  wire \DFF_520.CK ;
  wire \DFF_520.D ;
  wire \DFF_520.Q ;
  wire \DFF_521.CK ;
  wire \DFF_521.D ;
  wire \DFF_521.Q ;
  wire \DFF_522.CK ;
  wire \DFF_522.D ;
  wire \DFF_522.Q ;
  wire \DFF_523.CK ;
  wire \DFF_523.D ;
  wire \DFF_523.Q ;
  wire \DFF_524.CK ;
  wire \DFF_524.D ;
  wire \DFF_524.Q ;
  wire \DFF_525.CK ;
  wire \DFF_525.D ;
  wire \DFF_525.Q ;
  wire \DFF_526.CK ;
  wire \DFF_526.D ;
  wire \DFF_526.Q ;
  wire \DFF_527.CK ;
  wire \DFF_527.D ;
  wire \DFF_527.Q ;
  wire \DFF_528.CK ;
  wire \DFF_528.D ;
  wire \DFF_528.Q ;
  wire \DFF_529.CK ;
  wire \DFF_529.D ;
  wire \DFF_529.Q ;
  wire \DFF_53.CK ;
  wire \DFF_53.D ;
  wire \DFF_53.Q ;
  wire \DFF_530.CK ;
  wire \DFF_530.D ;
  wire \DFF_530.Q ;
  wire \DFF_531.CK ;
  wire \DFF_531.D ;
  wire \DFF_531.Q ;
  wire \DFF_532.CK ;
  wire \DFF_532.D ;
  wire \DFF_532.Q ;
  wire \DFF_533.CK ;
  wire \DFF_533.D ;
  wire \DFF_533.Q ;
  wire \DFF_54.CK ;
  wire \DFF_54.D ;
  wire \DFF_54.Q ;
  wire \DFF_55.CK ;
  wire \DFF_55.D ;
  wire \DFF_55.Q ;
  wire \DFF_56.CK ;
  wire \DFF_56.D ;
  wire \DFF_56.Q ;
  wire \DFF_57.CK ;
  wire \DFF_57.D ;
  wire \DFF_57.Q ;
  wire \DFF_58.CK ;
  wire \DFF_58.D ;
  wire \DFF_58.Q ;
  wire \DFF_59.CK ;
  wire \DFF_59.D ;
  wire \DFF_59.Q ;
  wire \DFF_6.CK ;
  wire \DFF_6.D ;
  wire \DFF_6.Q ;
  wire \DFF_60.CK ;
  wire \DFF_60.D ;
  wire \DFF_60.Q ;
  wire \DFF_61.CK ;
  wire \DFF_61.D ;
  wire \DFF_61.Q ;
  wire \DFF_62.CK ;
  wire \DFF_62.D ;
  wire \DFF_62.Q ;
  wire \DFF_63.CK ;
  wire \DFF_63.D ;
  wire \DFF_63.Q ;
  wire \DFF_64.CK ;
  wire \DFF_64.D ;
  wire \DFF_64.Q ;
  wire \DFF_65.CK ;
  wire \DFF_65.D ;
  wire \DFF_65.Q ;
  wire \DFF_66.CK ;
  wire \DFF_66.D ;
  wire \DFF_66.Q ;
  wire \DFF_67.CK ;
  wire \DFF_67.D ;
  wire \DFF_67.Q ;
  wire \DFF_68.CK ;
  wire \DFF_68.D ;
  wire \DFF_68.Q ;
  wire \DFF_69.CK ;
  wire \DFF_69.D ;
  wire \DFF_69.Q ;
  wire \DFF_7.CK ;
  wire \DFF_7.D ;
  wire \DFF_7.Q ;
  wire \DFF_70.CK ;
  wire \DFF_70.D ;
  wire \DFF_70.Q ;
  wire \DFF_71.CK ;
  wire \DFF_71.D ;
  wire \DFF_71.Q ;
  wire \DFF_72.CK ;
  wire \DFF_72.D ;
  wire \DFF_72.Q ;
  wire \DFF_73.CK ;
  wire \DFF_73.D ;
  wire \DFF_73.Q ;
  wire \DFF_74.CK ;
  wire \DFF_74.D ;
  wire \DFF_74.Q ;
  wire \DFF_75.CK ;
  wire \DFF_75.D ;
  wire \DFF_75.Q ;
  wire \DFF_76.CK ;
  wire \DFF_76.D ;
  wire \DFF_76.Q ;
  wire \DFF_77.CK ;
  wire \DFF_77.D ;
  wire \DFF_77.Q ;
  wire \DFF_78.CK ;
  wire \DFF_78.D ;
  wire \DFF_78.Q ;
  wire \DFF_79.CK ;
  wire \DFF_79.D ;
  wire \DFF_79.Q ;
  wire \DFF_8.CK ;
  wire \DFF_80.CK ;
  wire \DFF_80.D ;
  wire \DFF_80.Q ;
  wire \DFF_81.CK ;
  wire \DFF_81.D ;
  wire \DFF_81.Q ;
  wire \DFF_82.CK ;
  wire \DFF_82.D ;
  wire \DFF_82.Q ;
  wire \DFF_83.CK ;
  wire \DFF_83.D ;
  wire \DFF_83.Q ;
  wire \DFF_84.CK ;
  wire \DFF_85.CK ;
  wire \DFF_85.D ;
  wire \DFF_85.Q ;
  wire \DFF_86.CK ;
  wire \DFF_86.D ;
  wire \DFF_86.Q ;
  wire \DFF_87.CK ;
  wire \DFF_87.D ;
  wire \DFF_87.Q ;
  wire \DFF_88.CK ;
  wire \DFF_88.D ;
  wire \DFF_88.Q ;
  wire \DFF_89.CK ;
  wire \DFF_89.D ;
  wire \DFF_89.Q ;
  wire \DFF_9.CK ;
  wire \DFF_9.D ;
  wire \DFF_9.Q ;
  wire \DFF_90.CK ;
  wire \DFF_90.D ;
  wire \DFF_90.Q ;
  wire \DFF_91.CK ;
  wire \DFF_91.D ;
  wire \DFF_91.Q ;
  wire \DFF_92.CK ;
  wire \DFF_92.D ;
  wire \DFF_92.Q ;
  wire \DFF_93.CK ;
  wire \DFF_93.D ;
  wire \DFF_93.Q ;
  wire \DFF_94.CK ;
  wire \DFF_94.D ;
  wire \DFF_94.Q ;
  wire \DFF_95.CK ;
  wire \DFF_95.D ;
  wire \DFF_95.Q ;
  wire \DFF_96.CK ;
  wire \DFF_96.D ;
  wire \DFF_96.Q ;
  wire \DFF_97.CK ;
  wire \DFF_97.D ;
  wire \DFF_97.Q ;
  wire \DFF_98.CK ;
  wire \DFF_98.D ;
  wire \DFF_98.Q ;
  wire \DFF_99.CK ;
  wire \DFF_99.D ;
  wire \DFF_99.Q ;
  input GND;
  wire I10015;
  wire I10698;
  wire I11397;
  wire I11989;
  wire I12655;
  wire I12690;
  wire I13117;
  wire I13185;
  wire I16387;
  wire I5254;
  wire I5336;
  wire I5801;
  wire I5815;
  wire I5827;
  wire I5830;
  wire I5847;
  wire I5850;
  wire I5913;
  wire I5922;
  wire I5926;
  wire I5935;
  wire I5940;
  wire I5946;
  wire I5952;
  wire I5957;
  wire I5963;
  wire I5970;
  wire I5976;
  wire I5986;
  wire I5992;
  wire I5995;
  wire I5998;
  wire I6007;
  wire I6013;
  wire I6016;
  wire I6028;
  wire I6031;
  wire I6034;
  wire I6040;
  wire I6046;
  wire I6049;
  wire I6052;
  wire I6061;
  wire I6065;
  wire I6068;
  wire I6074;
  wire I6085;
  wire I6088;
  wire I6102;
  wire I6118;
  wire I6133;
  wire I6163;
  wire I6217;
  wire I6233;
  wire I6260;
  wire I6264;
  wire I6343;
  wire I6360;
  wire I6367;
  wire I6373;
  wire I6461;
  wire I6474;
  wire I6498;
  wire I6507;
  wire I6513;
  wire I6520;
  wire I6523;
  wire I6531;
  wire I6535;
  wire I6538;
  wire I6543;
  wire I6549;
  wire I6553;
  wire I6560;
  wire I6569;
  wire I6572;
  wire I6580;
  wire I6590;
  wire I6601;
  wire I6616;
  wire I6679;
  wire I6690;
  wire I6694;
  wire I6738;
  wire I6812;
  wire I6856;
  wire I6894;
  wire I6901;
  wire I6904;
  wire I6911;
  wire I6914;
  wire I6917;
  wire I6921;
  wire I6924;
  wire I6929;
  wire I6932;
  wire I6938;
  wire I6941;
  wire I6944;
  wire I6947;
  wire I6952;
  wire I6955;
  wire I6958;
  wire I6965;
  wire I6968;
  wire I6971;
  wire I6976;
  wire I6979;
  wire I6982;
  wire I6985;
  wire I6996;
  wire I6999;
  wire I7002;
  wire I7006;
  wire I7009;
  wire I7014;
  wire I7022;
  wire I7029;
  wire I7061;
  wire I7076;
  wire I7086;
  wire I7096;
  wire I7104;
  wire I7112;
  wire I7311;
  wire I7468;
  wire I7478;
  wire I7509;
  wire I7625;
  wire I7633;
  wire I7636;
  wire I7639;
  wire I7648;
  wire I7651;
  wire I7654;
  wire I7659;
  wire I7662;
  wire I7665;
  wire I7668;
  wire I7671;
  wire I7674;
  wire I7677;
  wire I7680;
  wire I7691;
  wire I7694;
  wire I7697;
  wire I7707;
  wire I7710;
  wire I7713;
  wire I7716;
  wire I7719;
  wire I7726;
  wire I7729;
  wire I7732;
  wire I7735;
  wire I7743;
  wire I7746;
  wire I7749;
  wire I7757;
  wire I7760;
  wire I7763;
  wire I7766;
  wire I7776;
  wire I7779;
  wire I7782;
  wire I7790;
  wire I7793;
  wire I7800;
  wire I7810;
  wire I7820;
  wire I7906;
  wire I8031;
  wire I8164;
  wire I8192;
  wire I8211;
  wire I8231;
  wire I8311;
  wire I8324;
  wire I8337;
  wire I8351;
  wire I8358;
  wire I8418;
  wire I9040;
  wire I9084;
  wire I9424;
  wire I9427;
  input VDD;
  wire g1;
  input g100;
  wire g1003;
  wire g1007;
  input g101;
  wire g1011;
  wire g1015;
  wire g1019;
  input g102;
  wire g1023;
  wire g1027;
  input g103;
  wire g1032;
  wire g10336;
  wire g10339;
  wire g1035;
  output g10377;
  wire g10378;
  output g10379;
  wire g1038;
  wire g10380;
  input g104;
  wire g10402;
  wire g10405;
  wire g10408;
  wire g1041;
  wire g10411;
  wire g10414;
  wire g10417;
  wire g1044;
  output g10455;
  wire g10456;
  output g10457;
  wire g10458;
  output g10459;
  wire g10460;
  output g10461;
  wire g10462;
  output g10463;
  wire g10464;
  output g10465;
  wire g10466;
  wire g1047;
  wire g105;
  wire g1050;
  wire g10515;
  wire g1053;
  wire g10531;
  wire g10532;
  wire g1056;
  wire g10575;
  wire g10576;
  wire g10577;
  wire g10578;
  wire g10579;
  wire g10580;
  wire g10583;
  wire g10589;
  wire g1059;
  wire g1062;
  output g10628;
  wire g1065;
  wire g10663;
  wire g10664;
  wire g1068;
  wire g10707;
  wire g1071;
  wire g10711;
  wire g10712;
  wire g10717;
  wire g10718;
  wire g10719;
  wire g10720;
  wire g10721;
  wire g10722;
  wire g10724;
  wire g10726;
  wire g10734;
  wire g10735;
  wire g1074;
  wire g10765;
  wire g10767;
  wire g1077;
  wire g10770;
  wire g10771;
  wire g10773;
  wire g10774;
  wire g10775;
  wire g10776;
  wire g10779;
  wire g10780;
  wire g10781;
  wire g10782;
  wire g10783;
  wire g10784;
  wire g10785;
  wire g10786;
  wire g10787;
  wire g10788;
  wire g10791;
  wire g10792;
  wire g10793;
  wire g10794;
  wire g10795;
  wire g10796;
  wire g10797;
  wire g10798;
  wire g10799;
  wire g108;
  wire g1080;
  wire g10800;
  output g10801;
  wire g10802;
  wire g10803;
  wire g10804;
  wire g10806;
  wire g10819;
  wire g10821;
  wire g10825;
  wire g10826;
  wire g1083;
  wire g10848;
  wire g10850;
  wire g10854;
  wire g10855;
  wire g10858;
  wire g10859;
  wire g1086;
  wire g10860;
  wire g10861;
  wire g10862;
  wire g10863;
  wire g10864;
  wire g10865;
  wire g10866;
  wire g10867;
  wire g10868;
  wire g10869;
  wire g10870;
  wire g10871;
  wire g10872;
  wire g10874;
  wire g10875;
  wire g10876;
  wire g10877;
  wire g10878;
  wire g10879;
  wire g10880;
  wire g10881;
  wire g10882;
  wire g10887;
  wire g10888;
  wire g10889;
  wire g1089;
  wire g10890;
  wire g10891;
  wire g10892;
  wire g10893;
  wire g10894;
  wire g10895;
  wire g10896;
  wire g10898;
  input g109;
  wire g10900;
  wire g10902;
  wire g10904;
  wire g10905;
  wire g10906;
  wire g10907;
  wire g10908;
  wire g10909;
  wire g10910;
  wire g10911;
  wire g10912;
  wire g10913;
  wire g1092;
  wire g10936;
  wire g1095;
  wire g10972;
  wire g10973;
  wire g1098;
  wire g110;
  wire g1101;
  wire g11014;
  wire g11033;
  wire g11034;
  wire g11035;
  wire g11036;
  wire g11037;
  wire g11038;
  wire g11039;
  wire g1104;
  wire g11040;
  wire g11041;
  wire g11042;
  wire g11043;
  wire g11044;
  wire g11047;
  wire g11048;
  wire g11049;
  wire g11050;
  wire g11051;
  wire g11052;
  wire g1107;
  wire g11074;
  wire g11076;
  wire g11079;
  wire g11080;
  wire g11081;
  wire g11082;
  wire g11084;
  wire g11086;
  wire g11088;
  wire g11096;
  wire g1110;
  wire g1113;
  output g11163;
  wire g1117;
  wire g11179;
  wire g11180;
  wire g11181;
  wire g11182;
  wire g11183;
  wire g11184;
  wire g11185;
  output g11206;
  wire g11207;
  wire g1121;
  wire g1125;
  wire g11256;
  wire g11257;
  wire g11258;
  wire g11259;
  wire g11260;
  wire g11261;
  wire g11262;
  wire g11263;
  wire g11264;
  wire g11265;
  wire g11266;
  wire g11267;
  wire g11268;
  wire g11269;
  wire g11270;
  wire g11286;
  wire g1129;
  wire g11290;
  wire g11291;
  wire g11292;
  wire g11293;
  wire g11294;
  wire g11298;
  wire g113;
  wire g11300;
  wire g11303;
  wire g11305;
  wire g11306;
  wire g11308;
  wire g11310;
  wire g11312;
  wire g11314;
  wire g11320;
  wire g11324;
  wire g11325;
  wire g11326;
  wire g11327;
  wire g11328;
  wire g11329;
  wire g1133;
  wire g11330;
  wire g11331;
  wire g11332;
  wire g11333;
  wire g11334;
  wire g11335;
  wire g11336;
  wire g11337;
  wire g11338;
  wire g11340;
  wire g11341;
  wire g11342;
  wire g11343;
  wire g11344;
  wire g11345;
  wire g11346;
  wire g11347;
  wire g11349;
  wire g11350;
  wire g11351;
  wire g11352;
  wire g11353;
  wire g1137;
  wire g11372;
  wire g11376;
  wire g11380;
  wire g11388;
  wire g11389;
  wire g11390;
  wire g11391;
  wire g11392;
  wire g11393;
  wire g11394;
  wire g11395;
  wire g11396;
  wire g11397;
  wire g11398;
  wire g11399;
  wire g114;
  wire g11400;
  wire g11401;
  wire g11402;
  wire g11403;
  wire g11404;
  wire g11405;
  wire g11406;
  wire g11408;
  wire g11409;
  wire g1141;
  wire g11410;
  wire g11411;
  wire g11412;
  wire g11417;
  wire g11419;
  wire g11420;
  wire g11421;
  wire g11423;
  wire g11424;
  wire g11436;
  wire g11437;
  wire g11438;
  wire g11439;
  wire g11440;
  wire g11441;
  wire g11442;
  wire g11443;
  wire g11444;
  wire g11445;
  wire g11446;
  wire g1145;
  wire g11450;
  wire g11451;
  wire g11453;
  wire g11454;
  wire g11457;
  wire g11466;
  wire g11467;
  wire g11468;
  wire g11469;
  wire g11470;
  wire g11471;
  wire g11472;
  wire g11473;
  wire g11478;
  wire g11481;
  wire g11482;
  wire g11483;
  wire g11484;
  wire g11485;
  wire g11486;
  wire g11487;
  wire g11488;
  output g11489;
  wire g1149;
  wire g11495;
  wire g11497;
  wire g11498;
  wire g11499;
  wire g115;
  wire g11500;
  wire g11501;
  wire g11502;
  wire g11503;
  wire g11504;
  wire g11505;
  wire g11506;
  wire g11507;
  wire g11508;
  wire g11509;
  wire g11510;
  wire g11511;
  wire g11512;
  wire g11513;
  wire g11514;
  wire g1153;
  wire g11550;
  wire g11561;
  wire g1157;
  wire g11577;
  wire g11578;
  wire g11579;
  wire g11593;
  wire g11594;
  wire g11598;
  wire g1160;
  wire g11602;
  wire g11603;
  wire g11604;
  wire g11605;
  wire g11606;
  wire g11607;
  wire g11608;
  wire g11609;
  wire g11610;
  wire g11611;
  wire g11614;
  wire g11616;
  wire g11617;
  wire g11618;
  wire g11619;
  wire g11620;
  wire g11621;
  wire g11622;
  wire g11623;
  wire g11625;
  wire g11627;
  wire g11628;
  wire g11629;
  wire g1163;
  wire g11630;
  wire g11631;
  wire g11632;
  wire g11633;
  wire g11634;
  wire g11635;
  wire g11636;
  wire g11638;
  wire g11639;
  wire g11640;
  wire g11641;
  wire g11642;
  wire g11643;
  wire g11644;
  wire g11645;
  wire g11646;
  wire g11647;
  wire g11648;
  wire g11649;
  wire g11650;
  wire g11651;
  wire g11652;
  wire g11653;
  wire g11654;
  wire g11655;
  wire g11656;
  wire g11657;
  wire g1166;
  input g1170;
  input g1173;
  input g1176;
  input g1179;
  input g1182;
  input g1185;
  input g1188;
  wire g119;
  input g1191;
  input g1194;
  input g1197;
  wire g12;
  input g1200;
  input g1203;
  wire g1206;
  wire g1212;
  wire g1216;
  wire g1217;
  wire g1218;
  wire g1223;
  wire g1227;
  wire g123;
  wire g1231;
  wire g1235;
  wire g1240;
  wire g1245;
  wire g1250;
  wire g1255;
  wire g1260;
  wire g1265;
  wire g127;
  wire g1270;
  wire g1275;
  wire g1280;
  wire g1284;
  wire g1289;
  wire g1292;
  wire g1296;
  wire g1300;
  wire g1304;
  wire g1308;
  wire g131;
  wire g1311;
  wire g1314;
  wire g1317;
  wire g1318;
  wire g1321;
  wire g1324;
  wire g1327;
  wire g1330;
  wire g1333;
  wire g1336;
  wire g1341;
  wire g1346;
  wire g135;
  wire g1351;
  wire g1356;
  wire g1357;
  wire g1360;
  wire g1361;
  wire g1362;
  wire g1365;
  wire g1368;
  wire g1371;
  wire g1374;
  wire g1377;
  wire g1380;
  wire g1383;
  wire g1386;
  wire g1389;
  wire g139;
  wire g1393;
  wire g1394;
  wire g1397;
  wire g1400;
  wire g1403;
  wire g1407;
  wire g1411;
  wire g1415;
  wire g1419;
  wire g1424;
  wire g1428;
  wire g143;
  wire g1432;
  wire g1436;
  wire g1440;
  wire g1444;
  wire g1448;
  wire g1453;
  wire g1458;
  wire g1462;
  wire g1466;
  wire g1470;
  wire g1474;
  wire g1478;
  wire g148;
  wire g1482;
  wire g1486;
  wire g1490;
  wire g1494;
  wire g1499;
  wire g1504;
  wire g1508;
  wire g1512;
  wire g1515;
  wire g1520;
  wire g1524;
  wire g1528;
  wire g153;
  wire g1531;
  wire g1534;
  wire g1537;
  wire g1540;
  wire g1543;
  wire g1546;
  wire g1549;
  wire g1552;
  wire g1555;
  wire g1558;
  wire g1561;
  wire g1564;
  wire g1567;
  wire g1571;
  wire g1574;
  wire g1577;
  wire g158;
  wire g1580;
  wire g1583;
  wire g1586;
  wire g1589;
  wire g1592;
  wire g1595;
  wire g1598;
  wire g16;
  wire g1601;
  wire g1604;
  wire g1607;
  wire g1610;
  wire g1615;
  wire g1618;
  wire g162;
  wire g1621;
  wire g1624;
  wire g1627;
  wire g1630;
  wire g1633;
  wire g1636;
  wire g1639;
  wire g1642;
  wire g1645;
  wire g1648;
  wire g1651;
  wire g1654;
  wire g1657;
  wire g166;
  wire g1660;
  wire g1663;
  wire g1666;
  wire g1669;
  wire g1672;
  wire g1675;
  wire g1678;
  wire g1681;
  wire g1684;
  wire g1687;
  wire g1690;
  input g1696;
  wire g17;
  wire g170;
  input g1700;
  wire g1703;
  wire g1707;
  wire g1710;
  input g1712;
  wire g1713;
  wire g1718;
  wire g1721;
  wire g1724;
  wire g1727;
  wire g1730;
  wire g1733;
  wire g1736;
  wire g1737;
  wire g1738;
  wire g174;
  wire g1741;
  wire g1744;
  wire g1747;
  wire g1750;
  wire g1753;
  wire g1756;
  wire g1759;
  wire g1762;
  wire g1765;
  wire g1766;
  wire g1771;
  wire g1776;
  wire g178;
  wire g1781;
  wire g1786;
  wire g1791;
  wire g1796;
  input g18;
  wire g1801;
  wire g1806;
  wire g1810;
  wire g1811;
  wire g1814;
  wire g182;
  wire g1822;
  wire g1828;
  wire g1834;
  wire g1840;
  wire g1845;
  wire g1848;
  wire g1849;
  wire g1850;
  wire g1853;
  wire g1854;
  wire g1857;
  wire g186;
  wire g1861;
  wire g1864;
  wire g1868;
  wire g1872;
  wire g1878;
  wire g1882;
  wire g1887;
  wire g1891;
  wire g1896;
  wire g1900;
  wire g1905;
  wire g1909;
  wire g1914;
  wire g1918;
  wire g192;
  wire g1923;
  wire g1927;
  wire g1932;
  wire g1936;
  wire g1941;
  wire g1945;
  wire g1950;
  wire g1955;
  wire g1956;
  output g1957;
  wire g1958;
  wire g1959;
  input g1960;
  input g1961;
  wire g197;
  wire g2004;
  wire g201;
  wire g2044;
  wire g2056;
  wire g2068;
  wire g2069;
  wire g207;
  wire g2071;
  wire g2072;
  wire g2073;
  wire g2075;
  wire g2076;
  wire g2079;
  wire g2080;
  wire g2084;
  wire g2085;
  wire g2086;
  wire g2089;
  wire g2090;
  wire g2094;
  wire g2097;
  wire g2098;
  wire g2100;
  wire g2101;
  wire g2103;
  wire g2108;
  wire g2110;
  wire g2116;
  wire g2119;
  wire g2121;
  wire g2122;
  wire g2123;
  wire g2124;
  wire g2125;
  wire g213;
  wire g2130;
  wire g2131;
  wire g2135;
  wire g2154;
  wire g2155;
  wire g2156;
  wire g2158;
  wire g2159;
  wire g2162;
  wire g2163;
  wire g2164;
  wire g2165;
  wire g2166;
  wire g2168;
  wire g2171;
  wire g2173;
  wire g2181;
  wire g219;
  wire g2190;
  wire g22;
  wire g2206;
  wire g2207;
  wire g2217;
  wire g2221;
  wire g2225;
  wire g2231;
  wire g2232;
  wire g2233;
  wire g2238;
  wire g2239;
  wire g2242;
  wire g2243;
  wire g2244;
  wire g2245;
  wire g2246;
  wire g2247;
  wire g225;
  wire g2252;
  wire g2255;
  wire g2256;
  wire g2258;
  wire g2259;
  wire g2267;
  wire g2269;
  wire g2270;
  wire g2296;
  wire g2298;
  input g23;
  wire g2304;
  wire g231;
  wire g2322;
  wire g2329;
  wire g2334;
  wire g2335;
  wire g2337;
  wire g2339;
  wire g2341;
  wire g2342;
  wire g2344;
  wire g2346;
  wire g2348;
  wire g2349;
  wire g2350;
  wire g2351;
  wire g2352;
  output g2355;
  wire g2356;
  wire g2363;
  wire g2368;
  wire g237;
  wire g2390;
  wire g2391;
  wire g2411;
  wire g2418;
  wire g243;
  wire g2431;
  wire g2432;
  wire g2436;
  wire g2454;
  wire g2462;
  wire g2478;
  wire g248;
  wire g2480;
  wire g2482;
  wire g2502;
  wire g2507;
  wire g2509;
  wire g2523;
  wire g2529;
  wire g253;
  wire g2530;
  wire g2537;
  wire g2539;
  wire g254;
  wire g2540;
  wire g2541;
  wire g2543;
  wire g2547;
  wire g2548;
  wire g255;
  wire g2554;
  wire g256;
  wire g2560;
  wire g2569;
  wire g257;
  wire g2578;
  wire g2579;
  wire g258;
  wire g2586;
  wire g259;
  wire g2593;
  wire g260;
  output g2601;
  output g2602;
  output g2603;
  output g2604;
  output g2605;
  output g2606;
  output g2607;
  output g2608;
  output g2609;
  wire g261;
  output g2610;
  output g2611;
  output g2612;
  wire g2613;
  wire g2614;
  wire g2617;
  wire g262;
  wire g2620;
  wire g2623;
  wire g2626;
  wire g2629;
  wire g263;
  wire g2632;
  wire g2635;
  wire g2638;
  wire g2639;
  wire g2640;
  wire g2641;
  wire g2642;
  wire g2643;
  wire g2644;
  wire g2645;
  wire g2646;
  wire g2647;
  output g2648;
  wire g2649;
  wire g2650;
  wire g2651;
  wire g2652;
  wire g2653;
  wire g2654;
  wire g2655;
  wire g266;
  wire g2662;
  wire g2669;
  wire g2677;
  wire g2683;
  wire g2689;
  wire g269;
  wire g2695;
  input g27;
  wire g2701;
  wire g2707;
  wire g2713;
  wire g2719;
  wire g272;
  wire g2725;
  wire g2726;
  wire g2727;
  wire g2728;
  wire g2731;
  wire g2732;
  wire g2733;
  wire g2742;
  wire g2745;
  wire g2748;
  wire g275;
  wire g2750;
  wire g2751;
  wire g2752;
  wire g2755;
  wire g2757;
  wire g2758;
  wire g2759;
  wire g2765;
  wire g2771;
  wire g2772;
  wire g2773;
  wire g2775;
  wire g2779;
  wire g278;
  wire g2791;
  wire g2797;
  wire g2798;
  input g28;
  wire g2809;
  wire g281;
  wire g2814;
  wire g2817;
  wire g2821;
  wire g2824;
  wire g2829;
  wire g2833;
  wire g284;
  wire g2840;
  wire g2844;
  wire g2847;
  wire g2851;
  wire g2855;
  wire g2861;
  wire g2864;
  wire g2868;
  wire g287;
  wire g2873;
  wire g2874;
  wire g2877;
  wire g2883;
  wire g2885;
  wire g2891;
  input g29;
  wire g290;
  wire g2902;
  wire g2906;
  wire g2908;
  wire g2909;
  wire g2914;
  wire g2915;
  wire g2916;
  wire g293;
  wire g2937;
  wire g2942;
  wire g2949;
  wire g2952;
  wire g2955;
  wire g2956;
  wire g2958;
  wire g296;
  wire g2960;
  wire g2962;
  wire g2964;
  wire g2965;
  wire g2971;
  wire g2980;
  output g2986;
  wire g299;
  wire g2994;
  input g30;
  output g3007;
  wire g3012;
  wire g302;
  wire g3038;
  wire g3044;
  wire g305;
  wire g3067;
  output g3069;
  wire g3076;
  wire g3077;
  wire g3088;
  wire g309;
  wire g3093;
  wire g3094;
  input g31;
  wire g3119;
  wire g312;
  wire g315;
  wire g3164;
  wire g318;
  wire g32;
  wire g3206;
  wire g321;
  wire g3213;
  wire g3214;
  wire g3219;
  wire g3220;
  wire g3226;
  wire g3227;
  wire g3228;
  wire g324;
  wire g3252;
  wire g3253;
  wire g3255;
  wire g3256;
  wire g3260;
  wire g3262;
  wire g3266;
  wire g3267;
  wire g327;
  wire g3271;
  wire g3272;
  wire g3274;
  wire g3292;
  wire g33;
  wire g330;
  wire g3306;
  wire g3307;
  wire g3318;
  wire g3321;
  wire g3323;
  wire g3326;
  output g3327;
  wire g3328;
  wire g3329;
  wire g333;
  wire g3331;
  wire g3334;
  wire g3344;
  wire g3353;
  wire g336;
  wire g3364;
  wire g3371;
  wire g3372;
  wire g3373;
  wire g3379;
  wire g3380;
  wire g3381;
  wire g3385;
  wire g3386;
  wire g3387;
  wire g339;
  wire g3390;
  wire g3391;
  wire g3392;
  wire g3393;
  wire g3394;
  wire g3397;
  wire g3398;
  wire g3399;
  wire g34;
  wire g3404;
  wire g3405;
  wire g3406;
  wire g3407;
  wire g3413;
  wire g3414;
  wire g3415;
  wire g3416;
  wire g3417;
  wire g3418;
  wire g342;
  wire g3424;
  wire g3425;
  wire g3426;
  wire g3427;
  wire g3428;
  wire g3431;
  wire g3432;
  wire g3433;
  wire g3435;
  wire g3436;
  wire g3437;
  wire g3438;
  wire g3439;
  wire g345;
  wire g3458;
  wire g3459;
  wire g3461;
  wire g3462;
  wire g3473;
  wire g3474;
  wire g348;
  wire g35;
  wire g3506;
  wire g351;
  wire g3524;
  wire g3538;
  wire g354;
  wire g3545;
  wire g357;
  wire g3583;
  wire g36;
  wire g360;
  wire g3621;
  wire g3622;
  wire g3624;
  wire g3627;
  wire g363;
  wire g3630;
  wire g3632;
  wire g3633;
  wire g3636;
  wire g3637;
  wire g366;
  wire g3663;
  wire g3682;
  wire g3683;
  wire g369;
  wire g3693;
  wire g3694;
  wire g3697;
  wire g37;
  wire g3703;
  wire g3704;
  wire g3705;
  wire g3707;
  wire g3708;
  wire g3715;
  wire g3716;
  wire g3719;
  wire g3720;
  wire g3721;
  wire g3726;
  wire g3729;
  wire g3737;
  wire g374;
  wire g3761;
  wire g378;
  wire g38;
  wire g3817;
  wire g382;
  wire g3828;
  wire g386;
  wire g3861;
  wire g3862;
  wire g3874;
  wire g3878;
  wire g39;
  wire g3905;
  wire g3909;
  wire g391;
  wire g3913;
  wire g3938;
  wire g3940;
  wire g3944;
  wire g3946;
  wire g396;
  wire g3975;
  wire g3980;
  wire g3982;
  wire g3988;
  wire g3990;
  wire g3995;
  wire g3996;
  wire g3997;
  wire g4;
  wire g40;
  wire g4002;
  wire g4003;
  wire g4004;
  wire g4005;
  wire g401;
  wire g4010;
  wire g4011;
  wire g4012;
  wire g4049;
  wire g4050;
  wire g4051;
  wire g4055;
  wire g4056;
  wire g4057;
  wire g406;
  wire g4060;
  wire g4061;
  wire g4062;
  wire g4066;
  wire g4067;
  wire g4076;
  wire g4077;
  wire g4078;
  wire g4080;
  wire g4081;
  wire g4082;
  wire g4083;
  wire g4087;
  wire g4089;
  wire g4095;
  wire g4096;
  wire g4098;
  input g41;
  wire g4102;
  wire g4105;
  wire g411;
  wire g4113;
  wire g4114;
  wire g4116;
  wire g4117;
  wire g4121;
  wire g4124;
  wire g4125;
  wire g4127;
  wire g4140;
  wire g4142;
  wire g4156;
  wire g4159;
  wire g416;
  wire g4160;
  wire g4166;
  wire g4167;
  output g4171;
  output g4172;
  output g4173;
  output g4174;
  output g4175;
  output g4176;
  output g4177;
  output g4178;
  output g4179;
  output g4180;
  output g4181;
  wire g4182;
  wire g4183;
  wire g4184;
  wire g4185;
  wire g4186;
  wire g4187;
  wire g4188;
  wire g4189;
  wire g4190;
  output g4191;
  output g4192;
  output g4193;
  output g4194;
  output g4195;
  output g4196;
  output g4197;
  output g4198;
  output g4199;
  input g42;
  output g4200;
  output g4201;
  output g4202;
  output g4203;
  output g4204;
  output g4205;
  output g4206;
  output g4207;
  output g4208;
  output g4209;
  wire g421;
  output g4210;
  output g4211;
  output g4212;
  output g4213;
  output g4214;
  output g4215;
  output g4216;
  wire g4217;
  wire g4219;
  wire g4231;
  wire g4232;
  wire g4238;
  wire g4239;
  wire g4255;
  wire g426;
  wire g4264;
  wire g4268;
  wire g4271;
  wire g4274;
  wire g4279;
  wire g4283;
  wire g4287;
  wire g4293;
  wire g4295;
  wire g4296;
  input g43;
  wire g4309;
  wire g431;
  wire g4310;
  wire g4317;
  wire g4322;
  wire g4325;
  wire g4327;
  wire g4330;
  wire g4331;
  wire g4334;
  wire g4335;
  wire g4338;
  wire g4340;
  wire g4342;
  wire g435;
  wire g4351;
  wire g4352;
  input g44;
  wire g440;
  wire g4414;
  wire g4425;
  wire g4437;
  wire g444;
  wire g4443;
  wire g4452;
  wire g4456;
  wire g4458;
  wire g4462;
  wire g4464;
  wire g4465;
  wire g4469;
  wire g4471;
  wire g4472;
  wire g4473;
  wire g4475;
  wire g4477;
  wire g448;
  wire g4480;
  wire g4484;
  wire g4485;
  wire g4490;
  wire g4491;
  wire g4495;
  wire g4496;
  wire g4498;
  wire g4499;
  input g45;
  wire g4500;
  wire g4504;
  wire g4506;
  wire g4507;
  wire g4510;
  wire g4513;
  wire g452;
  wire g4520;
  wire g4523;
  wire g4526;
  wire g4533;
  wire g4541;
  wire g4549;
  wire g4555;
  wire g4556;
  wire g456;
  wire g4562;
  wire g4577;
  wire g4589;
  wire g4590;
  input g46;
  wire g461;
  wire g4615;
  wire g4637;
  wire g466;
  wire g4674;
  wire g4678;
  wire g4681;
  input g47;
  wire g471;
  wire g4711;
  wire g4713;
  wire g4716;
  wire g4721;
  wire g4726;
  wire g4728;
  wire g4730;
  wire g4733;
  wire g4735;
  wire g4746;
  wire g4748;
  wire g4757;
  wire g476;
  wire g4762;
  wire g4767;
  wire g4773;
  wire g4781;
  wire g4785;
  wire g4786;
  wire g4789;
  wire g4790;
  wire g4791;
  input g48;
  wire g4802;
  wire g4805;
  wire g481;
  wire g486;
  output g4887;
  output g4888;
  wire g4890;
  wire g4891;
  wire g4892;
  wire g4893;
  wire g4894;
  wire g4895;
  wire g4896;
  wire g4897;
  wire g4898;
  wire g49;
  wire g4901;
  wire g4902;
  wire g4903;
  wire g4904;
  wire g4905;
  wire g4906;
  wire g4907;
  wire g4908;
  wire g491;
  wire g4915;
  wire g4933;
  wire g4934;
  wire g4935;
  wire g4940;
  wire g4942;
  wire g4944;
  wire g4951;
  wire g4954;
  wire g496;
  wire g4961;
  wire g4963;
  wire g4970;
  wire g5007;
  wire g501;
  wire g5011;
  wire g5012;
  wire g5027;
  wire g5032;
  wire g5033;
  wire g5035;
  wire g5037;
  wire g5040;
  wire g5047;
  wire g5050;
  wire g5052;
  wire g506;
  wire g5063;
  wire g5066;
  wire g5069;
  wire g5072;
  wire g5075;
  wire g5078;
  wire g5081;
  wire g5083;
  wire g5085;
  wire g5088;
  wire g5091;
  wire g5094;
  output g5101;
  wire g5102;
  output g5105;
  wire g5106;
  wire g5107;
  wire g5109;
  wire g511;
  wire g5111;
  wire g5114;
  wire g5120;
  wire g5126;
  wire g5127;
  wire g5128;
  wire g5148;
  wire g5149;
  wire g5151;
  wire g516;
  wire g5173;
  wire g5194;
  wire g5195;
  wire g5197;
  wire g5198;
  wire g52;
  wire g5205;
  wire g521;
  wire g5210;
  wire g5218;
  wire g5236;
  wire g5241;
  wire g5245;
  wire g525;
  wire g5253;
  wire g5262;
  wire g5265;
  wire g5270;
  wire g5272;
  wire g5275;
  wire g5281;
  wire g5284;
  wire g5287;
  wire g5288;
  wire g5291;
  wire g5296;
  wire g5299;
  wire g530;
  wire g5301;
  wire g5305;
  wire g5314;
  wire g5320;
  wire g534;
  wire g5344;
  wire g5348;
  wire g5353;
  wire g5354;
  wire g538;
  wire g5390;
  wire g5391;
  wire g5392;
  wire g5395;
  wire g5396;
  wire g5397;
  wire g5401;
  wire g5402;
  wire g5404;
  wire g5415;
  wire g5416;
  wire g5417;
  wire g5419;
  wire g542;
  wire g5421;
  wire g5445;
  wire g546;
  wire g5471;
  wire g5486;
  wire g549;
  wire g5494;
  wire g55;
  wire g5504;
  wire g5509;
  wire g5511;
  wire g5515;
  wire g5529;
  wire g5536;
  wire g554;
  wire g5543;
  wire g5556;
  wire g5567;
  wire g5568;
  wire g557;
  wire g5572;
  wire g5586;
  wire g5589;
  wire g5593;
  wire g5596;
  wire g560;
  wire g5603;
  wire g5615;
  wire g5620;
  wire g563;
  wire g5633;
  wire g5643;
  wire g5644;
  wire g5645;
  wire g5646;
  wire g5647;
  wire g5648;
  wire g5649;
  wire g5650;
  wire g5651;
  wire g5652;
  wire g5653;
  wire g5654;
  wire g5655;
  wire g5656;
  wire g5657;
  output g5658;
  output g5659;
  wire g566;
  wire g5660;
  wire g5661;
  wire g5662;
  wire g5663;
  wire g5664;
  wire g5665;
  wire g5666;
  wire g5667;
  wire g5668;
  wire g5669;
  wire g5670;
  wire g5671;
  wire g5672;
  wire g5673;
  wire g5676;
  wire g5677;
  wire g5679;
  wire g5682;
  wire g5683;
  wire g5685;
  wire g5688;
  wire g5689;
  wire g569;
  wire g5692;
  wire g5693;
  wire g5696;
  wire g5697;
  wire g5700;
  wire g5701;
  wire g5702;
  wire g5705;
  wire g5708;
  wire g5718;
  wire g5719;
  wire g572;
  wire g5723;
  wire g5724;
  wire g5727;
  wire g5728;
  wire g5729;
  wire g5730;
  wire g5734;
  wire g5735;
  wire g5736;
  wire g5741;
  wire g5742;
  wire g5743;
  wire g575;
  wire g5751;
  wire g5752;
  wire g5753;
  wire g5754;
  wire g5755;
  wire g5763;
  wire g5766;
  wire g5767;
  wire g5768;
  wire g5770;
  wire g5777;
  wire g5778;
  wire g5779;
  wire g578;
  wire g5787;
  wire g579;
  wire g5794;
  wire g58;
  wire g580;
  wire g5800;
  wire g581;
  wire g5811;
  wire g5815;
  output g5816;
  wire g5817;
  wire g582;
  wire g5821;
  wire g5826;
  wire g583;
  wire g5830;
  wire g5839;
  wire g584;
  wire g5843;
  wire g5844;
  wire g5849;
  wire g585;
  wire g5858;
  wire g586;
  wire g5862;
  wire g5864;
  wire g5865;
  wire g587;
  wire g5874;
  wire g5879;
  wire g588;
  wire g5884;
  wire g5887;
  wire g5889;
  wire g589;
  wire g590;
  wire g5904;
  wire g591;
  wire g5910;
  wire g5914;
  wire g5918;
  wire g5919;
  wire g5936;
  wire g5937;
  wire g5941;
  wire g5943;
  wire g5947;
  wire g5948;
  wire g5980;
  wire g5982;
  wire g5987;
  wire g599;
  wire g5992;
  wire g5994;
  wire g5996;
  wire g6000;
  wire g6002;
  wire g6015;
  wire g6026;
  wire g6030;
  wire g6035;
  wire g6036;
  wire g6038;
  wire g6040;
  wire g6042;
  wire g6045;
  wire g6049;
  wire g605;
  wire g6051;
  wire g6054;
  wire g6059;
  wire g6068;
  wire g6071;
  wire g6080;
  wire g6088;
  wire g6093;
  wire g6096;
  wire g6099;
  wire g61;
  wire g6100;
  wire g6103;
  wire g6104;
  wire g6106;
  wire g6107;
  wire g6108;
  wire g611;
  wire g6110;
  wire g6111;
  wire g6112;
  wire g6114;
  wire g6115;
  wire g6116;
  wire g6117;
  wire g6118;
  wire g6120;
  wire g6123;
  wire g6126;
  wire g6127;
  wire g6132;
  wire g6155;
  wire g6163;
  wire g617;
  wire g6179;
  wire g6180;
  wire g6193;
  wire g6198;
  wire g6205;
  wire g6215;
  wire g6216;
  wire g622;
  wire g6224;
  wire g6234;
  wire g6237;
  wire g6241;
  wire g6242;
  wire g6243;
  wire g6244;
  wire g6248;
  wire g6249;
  wire g6251;
  output g6253;
  output g6254;
  output g6255;
  output g6256;
  output g6257;
  output g6258;
  output g6259;
  output g6260;
  output g6261;
  output g6262;
  output g6263;
  output g6264;
  output g6265;
  output g6266;
  output g6267;
  output g6268;
  output g6269;
  wire g627;
  output g6270;
  output g6271;
  output g6272;
  output g6273;
  output g6274;
  output g6275;
  output g6276;
  output g6277;
  output g6278;
  output g6279;
  output g6280;
  output g6281;
  output g6282;
  output g6283;
  output g6284;
  output g6285;
  wire g6286;
  wire g6287;
  wire g6288;
  wire g6289;
  wire g6290;
  wire g6291;
  wire g6292;
  wire g6293;
  wire g6294;
  wire g6295;
  wire g6296;
  wire g6297;
  wire g6298;
  wire g6299;
  wire g630;
  wire g6300;
  wire g6301;
  wire g6302;
  wire g6303;
  wire g6304;
  wire g6305;
  wire g6306;
  wire g6307;
  wire g6308;
  wire g6309;
  wire g631;
  wire g6310;
  wire g6311;
  wire g6312;
  wire g6313;
  wire g632;
  wire g6330;
  wire g6331;
  wire g6332;
  wire g6333;
  wire g6334;
  wire g6336;
  wire g6337;
  wire g6338;
  wire g6339;
  wire g6340;
  wire g6344;
  wire g635;
  wire g636;
  wire g6365;
  wire g6382;
  wire g6386;
  wire g6388;
  wire g639;
  wire g6392;
  wire g6396;
  wire g6397;
  wire g6398;
  wire g6399;
  wire g64;
  wire g6406;
  wire g6412;
  wire g6419;
  wire g6426;
  wire g643;
  wire g6433;
  wire g6434;
  wire g6439;
  wire g6442;
  wire g6445;
  wire g6450;
  wire g6453;
  wire g6454;
  wire g646;
  wire g6468;
  wire g6469;
  wire g6470;
  wire g6471;
  wire g6478;
  wire g6479;
  wire g6480;
  wire g6481;
  wire g6482;
  wire g650;
  wire g6500;
  wire g6501;
  wire g6502;
  wire g6503;
  wire g6506;
  wire g6507;
  wire g6508;
  wire g6509;
  wire g6513;
  wire g6514;
  wire g6515;
  wire g6516;
  wire g6517;
  wire g6521;
  wire g6522;
  wire g6523;
  wire g6524;
  wire g6525;
  wire g6526;
  wire g6527;
  wire g6528;
  wire g6529;
  wire g6531;
  wire g6533;
  wire g6534;
  wire g6536;
  wire g6537;
  wire g6538;
  wire g6539;
  wire g654;
  wire g6541;
  wire g6542;
  wire g6543;
  wire g6545;
  wire g6546;
  wire g6547;
  wire g6551;
  wire g6553;
  wire g6558;
  wire g6571;
  wire g658;
  wire g6584;
  wire g6588;
  wire g6594;
  wire g6596;
  wire g6620;
  wire g6621;
  wire g6627;
  wire g6629;
  wire g6634;
  wire g6635;
  wire g6638;
  wire g664;
  wire g6641;
  wire g6644;
  wire g6648;
  wire g6649;
  wire g6652;
  wire g6653;
  wire g6656;
  wire g6657;
  wire g6660;
  wire g6667;
  wire g6670;
  wire g6672;
  wire g6674;
  wire g6679;
  wire g668;
  wire g6680;
  wire g6685;
  wire g6686;
  wire g6688;
  wire g6692;
  wire g6694;
  wire g6695;
  wire g6698;
  wire g67;
  wire g6703;
  wire g6705;
  wire g6706;
  wire g6708;
  wire g6710;
  wire g6715;
  wire g6717;
  wire g6719;
  wire g6723;
  wire g6728;
  wire g6729;
  wire g673;
  wire g6733;
  wire g6734;
  wire g6735;
  wire g6747;
  wire g6751;
  wire g6755;
  wire g6757;
  wire g6759;
  wire g677;
  wire g6786;
  wire g6793;
  wire g6795;
  wire g6796;
  wire g6797;
  wire g6798;
  wire g6799;
  wire g6800;
  wire g6801;
  wire g6802;
  wire g6803;
  wire g6804;
  wire g6805;
  wire g6806;
  wire g6807;
  wire g6808;
  wire g6809;
  wire g6810;
  wire g6811;
  wire g6812;
  wire g6813;
  wire g6814;
  wire g6815;
  wire g6816;
  wire g6817;
  wire g6818;
  wire g6819;
  wire g682;
  wire g6820;
  wire g6821;
  wire g6822;
  wire g6823;
  wire g6824;
  wire g6825;
  wire g6826;
  wire g6827;
  wire g6828;
  wire g6829;
  wire g6830;
  wire g6831;
  wire g6832;
  wire g6833;
  wire g6834;
  wire g6835;
  wire g6836;
  wire g6837;
  wire g6838;
  wire g6839;
  wire g6840;
  wire g6841;
  output g6842;
  wire g6843;
  wire g6844;
  wire g6845;
  wire g6846;
  wire g6852;
  wire g6854;
  wire g6857;
  wire g686;
  wire g6860;
  wire g6869;
  wire g6877;
  wire g6881;
  wire g6888;
  wire g6893;
  wire g6894;
  wire g6895;
  wire g6896;
  wire g6897;
  wire g6898;
  wire g6900;
  wire g6901;
  wire g6902;
  wire g6903;
  wire g6904;
  wire g6905;
  wire g6906;
  wire g6907;
  wire g6908;
  wire g6909;
  wire g691;
  wire g6910;
  wire g6911;
  wire g6912;
  wire g6913;
  wire g6914;
  wire g6915;
  wire g6916;
  wire g6918;
  wire g6919;
  output g6920;
  wire g6921;
  wire g6922;
  wire g6923;
  wire g6924;
  wire g6925;
  output g6926;
  wire g6927;
  wire g6928;
  wire g6929;
  wire g6930;
  wire g6931;
  output g6932;
  wire g6933;
  wire g6934;
  wire g6938;
  wire g6939;
  output g6942;
  wire g6943;
  wire g6947;
  wire g6948;
  output g6949;
  wire g695;
  wire g6950;
  wire g6954;
  output g6955;
  wire g6956;
  wire g6960;
  wire g6970;
  wire g6983;
  wire g6993;
  wire g7;
  wire g70;
  wire g700;
  wire g7007;
  wire g7008;
  wire g7009;
  wire g7010;
  wire g7020;
  wire g7021;
  wire g7023;
  wire g7024;
  wire g7026;
  wire g7027;
  wire g7029;
  wire g7030;
  wire g7032;
  wire g7033;
  wire g7034;
  wire g7035;
  wire g7037;
  wire g7038;
  wire g7039;
  wire g704;
  wire g7040;
  wire g7042;
  wire g7043;
  wire g7044;
  wire g7047;
  wire g7048;
  wire g7049;
  wire g7051;
  wire g7052;
  wire g7053;
  wire g7056;
  wire g7057;
  wire g7058;
  wire g7064;
  wire g7065;
  wire g7066;
  wire g7069;
  wire g7070;
  wire g7072;
  wire g7073;
  wire g7076;
  wire g7078;
  wire g7082;
  wire g7089;
  wire g709;
  wire g7093;
  wire g7097;
  wire g7098;
  wire g7103;
  wire g7106;
  wire g7107;
  wire g7110;
  wire g7113;
  wire g7116;
  wire g7119;
  wire g7122;
  wire g7126;
  wire g713;
  wire g7133;
  wire g7134;
  wire g7137;
  wire g7143;
  wire g7144;
  wire g7147;
  wire g718;
  wire g7183;
  wire g7187;
  wire g7189;
  wire g7191;
  wire g7192;
  wire g7195;
  wire g7202;
  wire g7203;
  wire g7204;
  wire g7211;
  wire g7212;
  wire g7218;
  wire g7219;
  wire g722;
  wire g7225;
  wire g7231;
  wire g7236;
  wire g7240;
  wire g7242;
  wire g7244;
  wire g7245;
  wire g7257;
  wire g7258;
  wire g727;
  wire g7284;
  wire g7285;
  wire g7287;
  wire g7288;
  wire g7289;
  wire g7290;
  wire g7291;
  wire g7292;
  wire g7293;
  wire g7294;
  wire g7295;
  wire g7296;
  wire g7297;
  wire g7298;
  wire g7299;
  wire g73;
  wire g7300;
  wire g7301;
  wire g7302;
  wire g7303;
  wire g7304;
  wire g7305;
  wire g7306;
  wire g7307;
  wire g7308;
  wire g7309;
  wire g731;
  wire g7310;
  wire g7311;
  wire g7312;
  wire g7313;
  wire g7314;
  wire g7315;
  wire g7316;
  wire g7317;
  wire g7318;
  wire g7319;
  wire g7320;
  wire g7321;
  wire g7322;
  wire g7323;
  wire g7324;
  wire g7325;
  wire g7326;
  wire g7327;
  wire g7328;
  wire g7329;
  wire g7330;
  wire g7331;
  wire g7332;
  wire g7333;
  wire g7334;
  wire g7335;
  wire g7336;
  wire g7337;
  wire g7338;
  wire g7339;
  wire g7340;
  wire g7341;
  wire g7342;
  wire g7343;
  wire g7344;
  wire g7345;
  wire g7346;
  wire g7347;
  wire g7348;
  wire g7349;
  wire g7350;
  wire g7351;
  wire g7352;
  wire g7353;
  wire g7354;
  wire g7355;
  wire g7356;
  wire g7357;
  wire g7358;
  wire g7359;
  wire g736;
  wire g7360;
  wire g7361;
  wire g7362;
  wire g7363;
  wire g7364;
  wire g7365;
  wire g7366;
  wire g7369;
  wire g7374;
  wire g7376;
  wire g7377;
  wire g7380;
  wire g7387;
  wire g7388;
  wire g7390;
  wire g7395;
  input g741;
  wire g7415;
  input g742;
  wire g7421;
  input g743;
  input g744;
  wire g7441;
  wire g7445;
  wire g7446;
  wire g745;
  wire g7450;
  wire g7454;
  wire g746;
  wire g7460;
  wire g7464;
  wire g7467;
  wire g7473;
  wire g7477;
  wire g7497;
  input g750;
  wire g7501;
  wire g7502;
  wire g7505;
  wire g7509;
  wire g7512;
  wire g7516;
  wire g7520;
  wire g7521;
  wire g7522;
  wire g7525;
  wire g7527;
  wire g7530;
  wire g7531;
  wire g7532;
  wire g7534;
  wire g7537;
  wire g7538;
  wire g7539;
  wire g754;
  wire g7540;
  wire g7541;
  wire g7543;
  wire g7544;
  wire g7545;
  wire g7546;
  wire g755;
  wire g7550;
  wire g7555;
  wire g7556;
  wire g7559;
  wire g756;
  wire g7560;
  wire g7561;
  wire g7562;
  wire g7568;
  wire g7569;
  wire g757;
  wire g7570;
  wire g7571;
  wire g7574;
  wire g7579;
  wire g758;
  wire g7580;
  wire g7581;
  wire g7585;
  wire g7586;
  wire g7589;
  wire g7590;
  wire g7594;
  wire g76;
  wire g7608;
  wire g7611;
  wire g7618;
  wire g7619;
  wire g762;
  wire g7626;
  wire g7627;
  wire g7628;
  wire g7629;
  wire g7630;
  wire g7631;
  wire g7632;
  wire g7633;
  wire g7634;
  wire g7635;
  wire g7636;
  wire g7637;
  wire g7648;
  wire g7649;
  wire g7650;
  wire g7656;
  wire g7657;
  wire g7658;
  wire g7659;
  wire g766;
  wire g7660;
  wire g7662;
  wire g7663;
  wire g7669;
  wire g7672;
  wire g7673;
  wire g7675;
  wire g7676;
  wire g7677;
  wire g7678;
  wire g7680;
  wire g7681;
  wire g7682;
  wire g7683;
  wire g7684;
  wire g7685;
  wire g7686;
  wire g7688;
  wire g7692;
  wire g7696;
  wire g770;
  wire g7705;
  wire g7706;
  wire g7709;
  wire g7723;
  wire g7724;
  wire g7725;
  wire g7726;
  wire g7727;
  wire g7728;
  wire g7729;
  wire g7731;
  wire g7733;
  wire g7735;
  wire g7737;
  wire g774;
  output g7744;
  wire g7745;
  wire g7746;
  wire g7747;
  wire g7748;
  wire g7749;
  wire g7750;
  wire g7751;
  wire g7752;
  wire g7753;
  wire g7754;
  wire g7755;
  wire g7756;
  wire g7757;
  wire g7758;
  wire g7759;
  wire g7760;
  wire g7761;
  wire g7762;
  wire g7763;
  wire g7764;
  wire g7765;
  wire g7766;
  wire g7767;
  wire g7768;
  wire g7769;
  wire g7770;
  wire g7771;
  wire g7772;
  wire g7773;
  wire g7774;
  wire g7775;
  wire g7776;
  wire g7777;
  wire g7778;
  wire g7779;
  wire g778;
  wire g7780;
  wire g7781;
  wire g7782;
  wire g7783;
  wire g7784;
  wire g7785;
  wire g7786;
  wire g7787;
  wire g7788;
  wire g7789;
  wire g7790;
  wire g7791;
  wire g7792;
  wire g7793;
  wire g7794;
  wire g7795;
  wire g7796;
  wire g7797;
  wire g7798;
  wire g7799;
  wire g7800;
  wire g7801;
  wire g7802;
  wire g7803;
  wire g7804;
  wire g7805;
  wire g7806;
  wire g7807;
  wire g7808;
  wire g7809;
  wire g7810;
  wire g7811;
  wire g7812;
  wire g7813;
  wire g7814;
  wire g7815;
  wire g7816;
  wire g7817;
  wire g782;
  wire g7843;
  wire g7844;
  wire g7845;
  wire g7848;
  wire g7849;
  wire g786;
  wire g7896;
  wire g7899;
  wire g79;
  wire g790;
  wire g7904;
  wire g7906;
  wire g7921;
  wire g7922;
  wire g7924;
  wire g7925;
  wire g7927;
  wire g7928;
  wire g7929;
  wire g7930;
  wire g794;
  wire g7959;
  wire g7966;
  wire g7975;
  wire g7976;
  wire g7977;
  wire g7979;
  wire g798;
  wire g7981;
  wire g7982;
  wire g7983;
  wire g7984;
  wire g7985;
  wire g7989;
  wire g7991;
  wire g7993;
  wire g7995;
  wire g7998;
  wire g7999;
  wire g8;
  wire g8001;
  wire g8002;
  wire g8003;
  wire g8004;
  wire g8007;
  wire g8008;
  wire g8009;
  wire g8019;
  wire g802;
  wire g8024;
  wire g8039;
  wire g8040;
  wire g8041;
  wire g8042;
  wire g8043;
  wire g8044;
  wire g8045;
  wire g8046;
  wire g8047;
  wire g8048;
  wire g8049;
  wire g8050;
  wire g8051;
  wire g8052;
  wire g8053;
  wire g8054;
  wire g8055;
  wire g8059;
  wire g806;
  wire g8060;
  output g8061;
  output g8062;
  wire g8063;
  wire g8064;
  wire g8065;
  wire g8066;
  wire g8067;
  wire g8076;
  wire g8077;
  wire g8078;
  wire g8079;
  wire g8080;
  wire g8093;
  wire g8096;
  wire g810;
  wire g8116;
  wire g8121;
  wire g8122;
  wire g8125;
  wire g8126;
  wire g8128;
  wire g8132;
  wire g8133;
  wire g8134;
  wire g8137;
  wire g8138;
  wire g814;
  wire g8140;
  wire g8141;
  wire g8142;
  wire g8144;
  wire g8145;
  wire g8147;
  wire g8149;
  wire g8150;
  wire g8152;
  wire g8155;
  wire g8156;
  wire g8160;
  wire g8164;
  wire g8171;
  wire g8173;
  wire g8178;
  wire g8179;
  wire g818;
  wire g8181;
  wire g8182;
  wire g8183;
  wire g8184;
  wire g8186;
  wire g8187;
  wire g8191;
  wire g8192;
  wire g8193;
  wire g8194;
  wire g8195;
  wire g8196;
  wire g8197;
  wire g8198;
  input g82;
  wire g8200;
  wire g8203;
  wire g8206;
  wire g8210;
  wire g8214;
  wire g822;
  wire g8221;
  wire g8226;
  wire g8230;
  wire g8233;
  wire g8236;
  wire g8241;
  wire g8244;
  wire g8245;
  wire g8250;
  wire g8251;
  wire g8254;
  wire g826;
  wire g8260;
  output g8271;
  wire g8272;
  wire g8273;
  wire g8274;
  wire g8275;
  wire g8276;
  wire g8277;
  wire g8278;
  wire g8279;
  wire g8280;
  wire g8281;
  wire g8282;
  wire g8283;
  wire g8284;
  wire g8285;
  wire g8286;
  wire g8287;
  wire g8288;
  wire g829;
  wire g8292;
  wire g8294;
  input g83;
  wire g8304;
  wire g8306;
  wire g8310;
  wire g8311;
  wire g8312;
  output g8313;
  wire g8314;
  wire g8315;
  output g8316;
  wire g8317;
  output g8318;
  wire g8319;
  wire g8320;
  wire g8321;
  output g8323;
  wire g8324;
  wire g8325;
  wire g8326;
  output g8328;
  wire g8329;
  wire g833;
  wire g8330;
  output g8331;
  wire g8332;
  wire g8333;
  wire g8334;
  output g8335;
  wire g8336;
  wire g8337;
  wire g8338;
  wire g8339;
  output g8340;
  wire g8341;
  wire g8342;
  wire g8343;
  wire g8344;
  wire g8345;
  wire g8346;
  output g8347;
  wire g8348;
  output g8349;
  wire g8350;
  wire g8351;
  output g8352;
  wire g8353;
  wire g8354;
  wire g8355;
  wire g8356;
  wire g8357;
  wire g8358;
  wire g8359;
  wire g8360;
  wire g8361;
  wire g8362;
  wire g8363;
  wire g837;
  wire g8375;
  wire g8376;
  wire g8378;
  wire g8379;
  wire g8381;
  wire g8384;
  input g84;
  wire g841;
  wire g8418;
  wire g8419;
  wire g8420;
  wire g8421;
  wire g8422;
  wire g8423;
  wire g8424;
  wire g8425;
  wire g8426;
  wire g8427;
  wire g8428;
  wire g8429;
  wire g8430;
  wire g8431;
  wire g8432;
  wire g8433;
  wire g8434;
  wire g8435;
  wire g8436;
  wire g8437;
  wire g8438;
  wire g8439;
  wire g8440;
  wire g8441;
  wire g8442;
  wire g8443;
  wire g8444;
  wire g8445;
  wire g8446;
  wire g8447;
  wire g8448;
  wire g8449;
  wire g845;
  wire g8450;
  wire g8472;
  wire g8473;
  wire g8476;
  wire g8478;
  wire g8480;
  wire g849;
  input g85;
  wire g8500;
  wire g8505;
  wire g8513;
  wire g8514;
  wire g8515;
  wire g8516;
  wire g8517;
  wire g8518;
  wire g8519;
  wire g853;
  wire g8559;
  wire g8560;
  output g8561;
  output g8562;
  output g8563;
  output g8564;
  output g8565;
  output g8566;
  wire g8567;
  wire g8568;
  wire g8569;
  wire g857;
  wire g8570;
  wire g8571;
  wire g8572;
  wire g8573;
  wire g8575;
  wire g8588;
  input g86;
  wire g8600;
  wire g8601;
  wire g8604;
  wire g8606;
  wire g8608;
  wire g861;
  wire g8610;
  wire g8613;
  wire g8622;
  wire g8624;
  wire g8625;
  wire g8626;
  wire g8631;
  wire g8649;
  wire g865;
  wire g8650;
  wire g868;
  wire g869;
  wire g8694;
  wire g8695;
  input g87;
  wire g8714;
  input g872;
  input g873;
  wire g874;
  wire g8747;
  wire g875;
  wire g8758;
  wire g876;
  wire g8765;
  wire g8766;
  wire g8767;
  wire g8768;
  wire g8769;
  input g877;
  wire g8770;
  wire g8771;
  wire g8772;
  wire g8773;
  wire g8774;
  wire g8775;
  wire g8776;
  wire g8777;
  wire g8779;
  wire g878;
  wire g8780;
  wire g8781;
  wire g8782;
  wire g8784;
  wire g8785;
  wire g8788;
  wire g8790;
  wire g8792;
  wire g8794;
  wire g8795;
  wire g8797;
  wire g8798;
  input g88;
  wire g8800;
  wire g8802;
  wire g8803;
  wire g8804;
  wire g8805;
  wire g8806;
  input g881;
  wire g8810;
  wire g8811;
  wire g8812;
  wire g8813;
  wire g8814;
  wire g8815;
  wire g8816;
  wire g8817;
  wire g8818;
  wire g8819;
  wire g882;
  wire g8820;
  wire g883;
  input g886;
  wire g8868;
  wire g8869;
  wire g8870;
  wire g8871;
  wire g8872;
  wire g8873;
  wire g8874;
  wire g8883;
  wire g8884;
  wire g8885;
  wire g8886;
  wire g8887;
  wire g8888;
  wire g8889;
  input g889;
  wire g8890;
  wire g8891;
  input g89;
  input g892;
  wire g8920;
  wire g8921;
  wire g8922;
  wire g8923;
  wire g8924;
  wire g8926;
  wire g8928;
  wire g8937;
  wire g8938;
  wire g8939;
  wire g8940;
  wire g8941;
  wire g8943;
  wire g8944;
  wire g8945;
  wire g8946;
  wire g8948;
  input g895;
  wire g8950;
  wire g8951;
  wire g8952;
  wire g8953;
  wire g8954;
  wire g8956;
  wire g8958;
  wire g8959;
  wire g8961;
  wire g8969;
  wire g8973;
  output g8976;
  output g8977;
  output g8978;
  output g8979;
  input g898;
  output g8980;
  output g8981;
  output g8982;
  output g8983;
  output g8984;
  output g8985;
  output g8986;
  wire g8987;
  wire g8988;
  wire g8989;
  wire g8990;
  wire g8991;
  wire g8992;
  wire g8993;
  wire g9;
  input g90;
  wire g9009;
  input g901;
  wire g9024;
  wire g9025;
  wire g9026;
  wire g9027;
  wire g9028;
  wire g9029;
  input g904;
  input g907;
  wire g9088;
  input g91;
  input g910;
  wire g9106;
  wire g9108;
  wire g9109;
  wire g9110;
  wire g9124;
  input g913;
  wire g9150;
  input g916;
  input g919;
  input g92;
  input g922;
  input g925;
  wire g9262;
  wire g9264;
  wire g9266;
  wire g9269;
  wire g9270;
  wire g9272;
  wire g9273;
  wire g928;
  wire g9290;
  input g93;
  wire g9308;
  wire g9310;
  wire g9311;
  wire g9312;
  wire g932;
  wire g9338;
  wire g9339;
  wire g9340;
  wire g9341;
  wire g9342;
  wire g9343;
  wire g9344;
  wire g9345;
  wire g9346;
  wire g9347;
  wire g9348;
  wire g9349;
  wire g9350;
  wire g9351;
  wire g9352;
  wire g9353;
  wire g9354;
  wire g9355;
  wire g9356;
  wire g936;
  wire g9360;
  input g94;
  wire g940;
  wire g944;
  output g9451;
  wire g9452;
  wire g947;
  input g95;
  wire g950;
  wire g9507;
  wire g9508;
  wire g9525;
  wire g9526;
  wire g953;
  wire g9532;
  wire g9533;
  wire g9535;
  wire g9555;
  wire g956;
  wire g959;
  input g96;
  wire g962;
  wire g965;
  wire g9661;
  wire g9666;
  wire g9670;
  wire g9671;
  wire g9672;
  wire g968;
  wire g97;
  wire g971;
  wire g9721;
  wire g9732;
  wire g9733;
  wire g976;
  wire g9762;
  wire g9763;
  wire g9765;
  wire g9767;
  wire g9769;
  wire g98;
  wire g981;
  wire g9813;
  wire g9818;
  wire g9819;
  wire g9820;
  wire g9821;
  wire g9822;
  wire g9823;
  wire g9824;
  wire g9825;
  wire g9826;
  wire g9827;
  wire g9832;
  wire g9845;
  wire g986;
  wire g9875;
  wire g9895;
  input g99;
  wire g991;
  wire g9919;
  wire g9930;
  wire g9931;
  wire g995;
  wire g9958;
  output g9961;
  wire g999;
  al_and3ftt _1417_ (
    .a(\DFF_194.Q ),
    .b(g109),
    .c(\DFF_328.Q ),
    .y(_0000_)
  );
  al_aoi21 _1418_ (
    .a(\DFF_335.Q ),
    .b(g109),
    .c(_0000_),
    .y(\DFF_226.D )
  );
  al_inv _1419_ (
    .a(g23),
    .y(g3327)
  );
  al_and3ftt _1420_ (
    .a(\DFF_332.Q ),
    .b(\DFF_346.Q ),
    .c(\DFF_523.Q ),
    .y(_0001_)
  );
  al_and2 _1421_ (
    .a(\DFF_103.Q ),
    .b(\DFF_268.Q ),
    .y(_0002_)
  );
  al_nand3 _1422_ (
    .a(\DFF_75.Q ),
    .b(\DFF_59.Q ),
    .c(_0002_),
    .y(_0003_)
  );
  al_and2 _1423_ (
    .a(\DFF_77.Q ),
    .b(\DFF_276.Q ),
    .y(_0004_)
  );
  al_nand3 _1424_ (
    .a(\DFF_324.Q ),
    .b(\DFF_104.Q ),
    .c(_0004_),
    .y(_0005_)
  );
  al_nor3ftt _1425_ (
    .a(_0001_),
    .b(_0003_),
    .c(_0005_),
    .y(\DFF_318.D )
  );
  al_and2ft _1426_ (
    .a(\DFF_77.Q ),
    .b(g1700),
    .y(\DFF_77.D )
  );
  al_and2ft _1427_ (
    .a(\DFF_431.Q ),
    .b(g750),
    .y(_0006_)
  );
  al_and2ft _1428_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .y(_0007_)
  );
  al_mux2h _1429_ (
    .a(_0006_),
    .b(_0007_),
    .s(\DFF_304.Q ),
    .y(\DFF_431.D )
  );
  al_inv _1430_ (
    .a(g1700),
    .y(\DFF_275.D )
  );
  al_inv _1431_ (
    .a(g47),
    .y(_0008_)
  );
  al_nand3fft _1432_ (
    .a(g41),
    .b(g31),
    .c(g48),
    .y(_0009_)
  );
  al_or3 _1433_ (
    .a(g41),
    .b(g30),
    .c(g48),
    .y(_0010_)
  );
  al_ao21 _1434_ (
    .a(_0009_),
    .b(_0010_),
    .c(_0008_),
    .y(_0011_)
  );
  al_inv _1435_ (
    .a(g41),
    .y(_0012_)
  );
  al_nor2 _1436_ (
    .a(g45),
    .b(g44),
    .y(_0013_)
  );
  al_nand3fft _1437_ (
    .a(g43),
    .b(g48),
    .c(_0013_),
    .y(_0014_)
  );
  al_or3fft _1438_ (
    .a(_0012_),
    .b(g42),
    .c(_0014_),
    .y(_0015_)
  );
  al_or3 _1439_ (
    .a(g46),
    .b(_0011_),
    .c(_0015_),
    .y(\DFF_137.D )
  );
  al_inv _1440_ (
    .a(\DFF_297.Q ),
    .y(_0016_)
  );
  al_or2 _1441_ (
    .a(\DFF_369.Q ),
    .b(\DFF_302.Q ),
    .y(_0017_)
  );
  al_aoi21ftf _1442_ (
    .a(\DFF_455.Q ),
    .b(_0017_),
    .c(_0016_),
    .y(\DFF_122.D )
  );
  al_ao21 _1443_ (
    .a(_0009_),
    .b(_0010_),
    .c(g47),
    .y(_0018_)
  );
  al_nand3ftt _1444_ (
    .a(g41),
    .b(g42),
    .c(g48),
    .y(_0019_)
  );
  al_and2 _1445_ (
    .a(g45),
    .b(g44),
    .y(_0020_)
  );
  al_nand3fft _1446_ (
    .a(g43),
    .b(_0019_),
    .c(_0020_),
    .y(_0021_)
  );
  al_nor3ftt _1447_ (
    .a(g46),
    .b(_0021_),
    .c(_0018_),
    .y(_0022_)
  );
  al_nand2ft _1448_ (
    .a(g44),
    .b(g45),
    .y(_0023_)
  );
  al_nor3ftt _1449_ (
    .a(g43),
    .b(_0019_),
    .c(_0023_),
    .y(_0024_)
  );
  al_or3fft _1450_ (
    .a(g46),
    .b(_0024_),
    .c(_0018_),
    .y(_0025_)
  );
  al_inv _1451_ (
    .a(g46),
    .y(_0026_)
  );
  al_and3ftt _1452_ (
    .a(g45),
    .b(g43),
    .c(g44),
    .y(_0027_)
  );
  al_nand2ft _1453_ (
    .a(_0019_),
    .b(_0027_),
    .y(_0028_)
  );
  al_or3 _1454_ (
    .a(_0026_),
    .b(_0028_),
    .c(_0018_),
    .y(_0029_)
  );
  al_and3ftt _1455_ (
    .a(_0022_),
    .b(_0025_),
    .c(_0029_),
    .y(_0030_)
  );
  al_and2ft _1456_ (
    .a(g31),
    .b(g48),
    .y(_0031_)
  );
  al_nand3fft _1457_ (
    .a(g41),
    .b(g42),
    .c(g48),
    .y(_0032_)
  );
  al_or3 _1458_ (
    .a(g43),
    .b(_0032_),
    .c(_0023_),
    .y(_0033_)
  );
  al_or3 _1459_ (
    .a(_0026_),
    .b(_0033_),
    .c(_0018_),
    .y(_0034_)
  );
  al_nand3ftt _1460_ (
    .a(g45),
    .b(g43),
    .c(g44),
    .y(_0035_)
  );
  al_nor3ftt _1461_ (
    .a(g46),
    .b(_0032_),
    .c(_0035_),
    .y(_0036_)
  );
  al_ao21ttf _1462_ (
    .a(_0009_),
    .b(_0010_),
    .c(_0036_),
    .y(_0037_)
  );
  al_and3 _1463_ (
    .a(_0031_),
    .b(_0037_),
    .c(_0034_),
    .y(_0038_)
  );
  al_ao21ftf _1464_ (
    .a(g41),
    .b(_0031_),
    .c(_0010_),
    .y(_0039_)
  );
  al_and3 _1465_ (
    .a(_0008_),
    .b(g46),
    .c(_0039_),
    .y(_0040_)
  );
  al_nand3fft _1466_ (
    .a(g45),
    .b(g43),
    .c(g44),
    .y(_0041_)
  );
  al_and3fft _1467_ (
    .a(g41),
    .b(_0041_),
    .c(g48),
    .y(_0042_)
  );
  al_and3fft _1468_ (
    .a(g46),
    .b(_0018_),
    .c(_0042_),
    .y(_0043_)
  );
  al_and3fft _1469_ (
    .a(g43),
    .b(g44),
    .c(g45),
    .y(_0044_)
  );
  al_and2ft _1470_ (
    .a(_0019_),
    .b(_0044_),
    .y(_0045_)
  );
  al_ao21 _1471_ (
    .a(_0045_),
    .b(_0040_),
    .c(_0043_),
    .y(_0046_)
  );
  al_and3ftt _1472_ (
    .a(_0046_),
    .b(_0038_),
    .c(_0030_),
    .y(_0047_)
  );
  al_nand3fft _1473_ (
    .a(g46),
    .b(_0018_),
    .c(_0045_),
    .y(_0048_)
  );
  al_or3 _1474_ (
    .a(g46),
    .b(_0033_),
    .c(_0018_),
    .y(_0049_)
  );
  al_and2ft _1475_ (
    .a(_0019_),
    .b(_0027_),
    .y(_0050_)
  );
  al_nand2ft _1476_ (
    .a(_0032_),
    .b(_0027_),
    .y(_0051_)
  );
  al_and3 _1477_ (
    .a(_0008_),
    .b(_0026_),
    .c(_0039_),
    .y(_0052_)
  );
  al_ao21ftf _1478_ (
    .a(_0050_),
    .b(_0051_),
    .c(_0052_),
    .y(_0053_)
  );
  al_and3 _1479_ (
    .a(_0048_),
    .b(_0049_),
    .c(_0053_),
    .y(_0054_)
  );
  al_and3 _1480_ (
    .a(g47),
    .b(_0026_),
    .c(_0039_),
    .y(_0055_)
  );
  al_and2ft _1481_ (
    .a(_0032_),
    .b(_0044_),
    .y(_0056_)
  );
  al_ao21ftf _1482_ (
    .a(_0056_),
    .b(_0028_),
    .c(_0055_),
    .y(_0057_)
  );
  al_and3 _1483_ (
    .a(g45),
    .b(g43),
    .c(g44),
    .y(_0058_)
  );
  al_and3fft _1484_ (
    .a(g46),
    .b(_0011_),
    .c(_0058_),
    .y(_0059_)
  );
  al_nand3 _1485_ (
    .a(_0012_),
    .b(g48),
    .c(_0059_),
    .y(_0060_)
  );
  al_and3 _1486_ (
    .a(_0057_),
    .b(_0060_),
    .c(_0054_),
    .y(_0061_)
  );
  al_and3fft _1487_ (
    .a(_0032_),
    .b(_0018_),
    .c(_0026_),
    .y(_0062_)
  );
  al_and3fft _1488_ (
    .a(g45),
    .b(g44),
    .c(g43),
    .y(_0063_)
  );
  al_nor3fft _1489_ (
    .a(g43),
    .b(_0013_),
    .c(_0019_),
    .y(_0064_)
  );
  al_nor3fft _1490_ (
    .a(_0026_),
    .b(_0064_),
    .c(_0018_),
    .y(_0065_)
  );
  al_aoi21 _1491_ (
    .a(_0063_),
    .b(_0062_),
    .c(_0065_),
    .y(_0066_)
  );
  al_nand3 _1492_ (
    .a(_0066_),
    .b(_0047_),
    .c(_0061_),
    .y(_0067_)
  );
  al_or3 _1493_ (
    .a(g46),
    .b(_0032_),
    .c(_0018_),
    .y(_0068_)
  );
  al_mux2l _1494_ (
    .a(_0041_),
    .b(_0068_),
    .s(\DFF_390.Q ),
    .y(_0069_)
  );
  al_nand3fft _1495_ (
    .a(\DFF_511.Q ),
    .b(_0041_),
    .c(_0062_),
    .y(_0070_)
  );
  al_or3fft _1496_ (
    .a(_0043_),
    .b(_0070_),
    .c(_0069_),
    .y(_0071_)
  );
  al_and3ftt _1497_ (
    .a(_0032_),
    .b(_0058_),
    .c(_0055_),
    .y(_0072_)
  );
  al_and3ftt _1498_ (
    .a(_0019_),
    .b(\DFF_321.Q ),
    .c(_0059_),
    .y(_0073_)
  );
  al_aoi21 _1499_ (
    .a(\DFF_410.Q ),
    .b(_0072_),
    .c(_0073_),
    .y(_0074_)
  );
  al_or3 _1500_ (
    .a(g46),
    .b(_0051_),
    .c(_0018_),
    .y(_0075_)
  );
  al_nand3 _1501_ (
    .a(\DFF_122.Q ),
    .b(_0063_),
    .c(_0062_),
    .y(_0076_)
  );
  al_ao21ftf _1502_ (
    .a(_0075_),
    .b(\DFF_256.Q ),
    .c(_0076_),
    .y(_0077_)
  );
  al_nand3ftt _1503_ (
    .a(_0077_),
    .b(_0071_),
    .c(_0074_),
    .y(_0078_)
  );
  al_nand3 _1504_ (
    .a(g1182),
    .b(_0050_),
    .c(_0055_),
    .y(_0079_)
  );
  al_aoi21ftf _1505_ (
    .a(_0029_),
    .b(g910),
    .c(_0079_),
    .y(_0080_)
  );
  al_nand3 _1506_ (
    .a(\DFF_445.Q ),
    .b(_0064_),
    .c(_0052_),
    .y(_0081_)
  );
  al_nand3 _1507_ (
    .a(\DFF_426.Q ),
    .b(_0050_),
    .c(_0052_),
    .y(_0082_)
  );
  al_nand3 _1508_ (
    .a(\DFF_20.Q ),
    .b(_0045_),
    .c(_0052_),
    .y(_0083_)
  );
  al_nand3 _1509_ (
    .a(_0081_),
    .b(_0082_),
    .c(_0083_),
    .y(_0084_)
  );
  al_and3 _1510_ (
    .a(\DFF_195.Q ),
    .b(_0056_),
    .c(_0055_),
    .y(_0085_)
  );
  al_and3 _1511_ (
    .a(\DFF_148.Q ),
    .b(_0056_),
    .c(_0040_),
    .y(_0086_)
  );
  al_oa21ftt _1512_ (
    .a(g48),
    .b(g31),
    .c(\DFF_350.Q ),
    .y(_0087_)
  );
  al_oa21ftf _1513_ (
    .a(\DFF_81.Q ),
    .b(_0049_),
    .c(_0087_),
    .y(_0088_)
  );
  al_nand3fft _1514_ (
    .a(_0085_),
    .b(_0086_),
    .c(_0088_),
    .y(_0089_)
  );
  al_nor3ftt _1515_ (
    .a(_0080_),
    .b(_0084_),
    .c(_0089_),
    .y(_0090_)
  );
  al_nand3ftt _1516_ (
    .a(_0078_),
    .b(_0090_),
    .c(_0067_),
    .y(\DFF_350.D )
  );
  al_ao21ftf _1517_ (
    .a(_0045_),
    .b(_0033_),
    .c(_0052_),
    .y(_0091_)
  );
  al_and3ftt _1518_ (
    .a(_0019_),
    .b(_0058_),
    .c(_0055_),
    .y(_0092_)
  );
  al_and3ftt _1519_ (
    .a(_0092_),
    .b(_0091_),
    .c(_0053_),
    .y(_0093_)
  );
  al_ao21ftf _1520_ (
    .a(_0045_),
    .b(_0028_),
    .c(_0055_),
    .y(_0094_)
  );
  al_nand3 _1521_ (
    .a(_0094_),
    .b(_0093_),
    .c(_0047_),
    .y(_0095_)
  );
  al_nand3 _1522_ (
    .a(\DFF_481.Q ),
    .b(_0045_),
    .c(_0055_),
    .y(_0096_)
  );
  al_nand3 _1523_ (
    .a(g1191),
    .b(_0050_),
    .c(_0055_),
    .y(_0097_)
  );
  al_and2 _1524_ (
    .a(\DFF_123.Q ),
    .b(_0032_),
    .y(_0098_)
  );
  al_nand3 _1525_ (
    .a(_0042_),
    .b(_0098_),
    .c(_0052_),
    .y(_0099_)
  );
  al_aoi21ftf _1526_ (
    .a(_0048_),
    .b(\DFF_138.Q ),
    .c(_0099_),
    .y(_0100_)
  );
  al_and3 _1527_ (
    .a(_0096_),
    .b(_0097_),
    .c(_0100_),
    .y(_0101_)
  );
  al_nand3ftt _1528_ (
    .a(_0019_),
    .b(\DFF_131.Q ),
    .c(_0059_),
    .y(_0102_)
  );
  al_nand3fft _1529_ (
    .a(_0026_),
    .b(_0018_),
    .c(_0045_),
    .y(_0103_)
  );
  al_oa21ftt _1530_ (
    .a(g48),
    .b(g31),
    .c(\DFF_319.Q ),
    .y(_0104_)
  );
  al_oa21ftf _1531_ (
    .a(\DFF_454.Q ),
    .b(_0103_),
    .c(_0104_),
    .y(_0105_)
  );
  al_or3 _1532_ (
    .a(g46),
    .b(_0028_),
    .c(_0018_),
    .y(_0106_)
  );
  al_nand3 _1533_ (
    .a(g919),
    .b(_0050_),
    .c(_0040_),
    .y(_0107_)
  );
  al_mux2h _1534_ (
    .a(_0032_),
    .b(_0035_),
    .s(\DFF_258.Q ),
    .y(_0108_)
  );
  al_aoi21ftf _1535_ (
    .a(_0106_),
    .b(_0108_),
    .c(_0107_),
    .y(_0109_)
  );
  al_and3 _1536_ (
    .a(_0102_),
    .b(_0105_),
    .c(_0109_),
    .y(_0110_)
  );
  al_nand3 _1537_ (
    .a(_0101_),
    .b(_0110_),
    .c(_0095_),
    .y(\DFF_319.D )
  );
  al_nand3 _1538_ (
    .a(\DFF_269.Q ),
    .b(g109),
    .c(\DFF_319.D ),
    .y(_0111_)
  );
  al_aoi21ttf _1539_ (
    .a(_0000_),
    .b(\DFF_350.D ),
    .c(_0111_),
    .y(_0112_)
  );
  al_and2 _1540_ (
    .a(\DFF_335.Q ),
    .b(g109),
    .y(_0113_)
  );
  al_and3 _1541_ (
    .a(_0053_),
    .b(_0091_),
    .c(_0060_),
    .y(_0114_)
  );
  al_and3ftt _1542_ (
    .a(_0043_),
    .b(_0103_),
    .c(_0038_),
    .y(_0115_)
  );
  al_and3 _1543_ (
    .a(_0066_),
    .b(_0030_),
    .c(_0115_),
    .y(_0116_)
  );
  al_or3 _1544_ (
    .a(g46),
    .b(_0033_),
    .c(_0011_),
    .y(_0117_)
  );
  al_or3 _1545_ (
    .a(g46),
    .b(_0051_),
    .c(_0011_),
    .y(_0118_)
  );
  al_and3 _1546_ (
    .a(_0117_),
    .b(_0118_),
    .c(_0094_),
    .y(_0119_)
  );
  al_nand3 _1547_ (
    .a(_0114_),
    .b(_0119_),
    .c(_0116_),
    .y(_0120_)
  );
  al_nand3 _1548_ (
    .a(\DFF_267.Q ),
    .b(_0064_),
    .c(_0052_),
    .y(_0121_)
  );
  al_aoi21ttf _1549_ (
    .a(\DFF_13.Q ),
    .b(_0022_),
    .c(_0121_),
    .y(_0122_)
  );
  al_and2ft _1550_ (
    .a(_0032_),
    .b(_0027_),
    .y(_0123_)
  );
  al_nand3 _1551_ (
    .a(g1203),
    .b(_0123_),
    .c(_0055_),
    .y(_0124_)
  );
  al_ao21ftf _1552_ (
    .a(_0103_),
    .b(\DFF_293.Q ),
    .c(_0124_),
    .y(_0125_)
  );
  al_nor3fft _1553_ (
    .a(_0026_),
    .b(_0045_),
    .c(_0018_),
    .y(_0126_)
  );
  al_nand3 _1554_ (
    .a(\DFF_392.Q ),
    .b(_0049_),
    .c(_0126_),
    .y(_0127_)
  );
  al_oai21ftt _1555_ (
    .a(g48),
    .b(g31),
    .c(\DFF_228.Q ),
    .y(_0128_)
  );
  al_nand3 _1556_ (
    .a(\DFF_106.Q ),
    .b(_0056_),
    .c(_0040_),
    .y(_0129_)
  );
  al_and3 _1557_ (
    .a(_0128_),
    .b(_0129_),
    .c(_0127_),
    .y(_0130_)
  );
  al_and3ftt _1558_ (
    .a(_0125_),
    .b(_0122_),
    .c(_0130_),
    .y(_0131_)
  );
  al_nand3 _1559_ (
    .a(\DFF_325.Q ),
    .b(_0056_),
    .c(_0055_),
    .y(_0132_)
  );
  al_nand3 _1560_ (
    .a(g1179),
    .b(_0050_),
    .c(_0055_),
    .y(_0133_)
  );
  al_and3 _1561_ (
    .a(\DFF_506.Q ),
    .b(_0045_),
    .c(_0055_),
    .y(_0134_)
  );
  al_and3ftt _1562_ (
    .a(_0134_),
    .b(_0132_),
    .c(_0133_),
    .y(_0135_)
  );
  al_nand3 _1563_ (
    .a(g907),
    .b(_0050_),
    .c(_0040_),
    .y(_0136_)
  );
  al_nand3 _1564_ (
    .a(g895),
    .b(_0024_),
    .c(_0040_),
    .y(_0137_)
  );
  al_nand3 _1565_ (
    .a(\DFF_218.Q ),
    .b(_0056_),
    .c(_0052_),
    .y(_0138_)
  );
  al_aoi21ftf _1566_ (
    .a(_0075_),
    .b(\DFF_10.Q ),
    .c(_0138_),
    .y(_0139_)
  );
  al_and3 _1567_ (
    .a(_0136_),
    .b(_0137_),
    .c(_0139_),
    .y(_0140_)
  );
  al_and3 _1568_ (
    .a(_0135_),
    .b(_0140_),
    .c(_0131_),
    .y(_0141_)
  );
  al_mux2l _1569_ (
    .a(_0041_),
    .b(_0068_),
    .s(\DFF_345.Q ),
    .y(_0142_)
  );
  al_nand3fft _1570_ (
    .a(\DFF_279.Q ),
    .b(_0041_),
    .c(_0062_),
    .y(_0143_)
  );
  al_or3fft _1571_ (
    .a(_0043_),
    .b(_0143_),
    .c(_0142_),
    .y(_0144_)
  );
  al_nand3ftt _1572_ (
    .a(_0019_),
    .b(\DFF_96.Q ),
    .c(_0059_),
    .y(_0145_)
  );
  al_ao21ftf _1573_ (
    .a(_0106_),
    .b(\DFF_42.Q ),
    .c(_0145_),
    .y(_0146_)
  );
  al_and3 _1574_ (
    .a(\DFF_262.Q ),
    .b(_0063_),
    .c(_0062_),
    .y(_0147_)
  );
  al_aoi21 _1575_ (
    .a(\DFF_200.Q ),
    .b(_0072_),
    .c(_0147_),
    .y(_0148_)
  );
  al_and3ftt _1576_ (
    .a(_0146_),
    .b(_0144_),
    .c(_0148_),
    .y(_0149_)
  );
  al_nand3 _1577_ (
    .a(_0149_),
    .b(_0120_),
    .c(_0141_),
    .y(\DFF_228.D )
  );
  al_and2 _1578_ (
    .a(_0113_),
    .b(\DFF_228.D ),
    .y(_0150_)
  );
  al_inv _1579_ (
    .a(g109),
    .y(_0151_)
  );
  al_nand3 _1580_ (
    .a(_0057_),
    .b(_0114_),
    .c(_0047_),
    .y(_0152_)
  );
  al_nand3ftt _1581_ (
    .a(_0032_),
    .b(\DFF_78.Q ),
    .c(_0059_),
    .y(_0153_)
  );
  al_nand3 _1582_ (
    .a(g1185),
    .b(_0050_),
    .c(_0055_),
    .y(_0154_)
  );
  al_oai21ftt _1583_ (
    .a(g48),
    .b(g31),
    .c(\DFF_116.Q ),
    .y(_0155_)
  );
  al_nand3 _1584_ (
    .a(_0155_),
    .b(_0154_),
    .c(_0153_),
    .y(_0156_)
  );
  al_nand3 _1585_ (
    .a(\DFF_181.Q ),
    .b(_0056_),
    .c(_0040_),
    .y(_0157_)
  );
  al_ao21ftf _1586_ (
    .a(_0029_),
    .b(g913),
    .c(_0157_),
    .y(_0158_)
  );
  al_nand3 _1587_ (
    .a(\DFF_477.Q ),
    .b(_0044_),
    .c(_0062_),
    .y(_0159_)
  );
  al_or3ftt _1588_ (
    .a(_0159_),
    .b(_0158_),
    .c(_0156_),
    .y(_0160_)
  );
  al_nand3fft _1589_ (
    .a(\DFF_229.Q ),
    .b(_0041_),
    .c(_0062_),
    .y(_0161_)
  );
  al_mux2l _1590_ (
    .a(_0041_),
    .b(_0068_),
    .s(\DFF_46.Q ),
    .y(_0162_)
  );
  al_or3fft _1591_ (
    .a(_0043_),
    .b(_0161_),
    .c(_0162_),
    .y(_0163_)
  );
  al_inv _1592_ (
    .a(\DFF_326.Q ),
    .y(_0164_)
  );
  al_nand3fft _1593_ (
    .a(_0019_),
    .b(_0035_),
    .c(_0052_),
    .y(_0165_)
  );
  al_nand3 _1594_ (
    .a(\DFF_254.Q ),
    .b(_0045_),
    .c(_0052_),
    .y(_0166_)
  );
  al_mux2h _1595_ (
    .a(_0164_),
    .b(_0165_),
    .s(_0166_),
    .y(_0167_)
  );
  al_nand3 _1596_ (
    .a(\DFF_432.Q ),
    .b(_0056_),
    .c(_0055_),
    .y(_0168_)
  );
  al_ao21ftf _1597_ (
    .a(_0075_),
    .b(\DFF_130.Q ),
    .c(_0168_),
    .y(_0169_)
  );
  al_and3ftt _1598_ (
    .a(_0169_),
    .b(_0167_),
    .c(_0163_),
    .y(_0170_)
  );
  al_nand3ftt _1599_ (
    .a(_0160_),
    .b(_0170_),
    .c(_0152_),
    .y(\DFF_116.D )
  );
  al_nand3fft _1600_ (
    .a(_0151_),
    .b(\DFF_161.Q ),
    .c(\DFF_116.D ),
    .y(_0171_)
  );
  al_nand3fft _1601_ (
    .a(g46),
    .b(_0011_),
    .c(_0045_),
    .y(_0172_)
  );
  al_nand3 _1602_ (
    .a(_0172_),
    .b(_0047_),
    .c(_0061_),
    .y(_0173_)
  );
  al_and3 _1603_ (
    .a(\DFF_466.Q ),
    .b(_0045_),
    .c(_0052_),
    .y(_0174_)
  );
  al_nor3ftt _1604_ (
    .a(_0026_),
    .b(_0028_),
    .c(_0011_),
    .y(_0175_)
  );
  al_oai21ftt _1605_ (
    .a(g48),
    .b(g31),
    .c(\DFF_22.Q ),
    .y(_0176_)
  );
  al_oa21ftt _1606_ (
    .a(_0036_),
    .b(_0011_),
    .c(_0176_),
    .y(_0177_)
  );
  al_ao21ttf _1607_ (
    .a(g1188),
    .b(_0175_),
    .c(_0177_),
    .y(_0178_)
  );
  al_and3ftt _1608_ (
    .a(_0032_),
    .b(\DFF_282.Q ),
    .c(_0059_),
    .y(_0179_)
  );
  al_aoi21 _1609_ (
    .a(\DFF_272.Q ),
    .b(_0092_),
    .c(_0179_),
    .y(_0180_)
  );
  al_nand3fft _1610_ (
    .a(_0174_),
    .b(_0178_),
    .c(_0180_),
    .y(_0181_)
  );
  al_nand3 _1611_ (
    .a(g916),
    .b(_0050_),
    .c(_0040_),
    .y(_0182_)
  );
  al_nand3 _1612_ (
    .a(\DFF_312.Q ),
    .b(_0045_),
    .c(_0040_),
    .y(_0183_)
  );
  al_and3 _1613_ (
    .a(\DFF_134.Q ),
    .b(_0045_),
    .c(_0055_),
    .y(_0184_)
  );
  al_and3ftt _1614_ (
    .a(_0184_),
    .b(_0182_),
    .c(_0183_),
    .y(_0185_)
  );
  al_nand3 _1615_ (
    .a(\DFF_351.Q ),
    .b(_0056_),
    .c(_0040_),
    .y(_0186_)
  );
  al_aoi21ftf _1616_ (
    .a(_0117_),
    .b(\DFF_146.Q ),
    .c(_0186_),
    .y(_0187_)
  );
  al_nand3 _1617_ (
    .a(\DFF_133.Q ),
    .b(_0032_),
    .c(_0043_),
    .y(_0188_)
  );
  al_aoi21ftf _1618_ (
    .a(_0106_),
    .b(\DFF_39.Q ),
    .c(_0188_),
    .y(_0189_)
  );
  al_and3 _1619_ (
    .a(_0187_),
    .b(_0189_),
    .c(_0185_),
    .y(_0190_)
  );
  al_nand3ftt _1620_ (
    .a(_0181_),
    .b(_0190_),
    .c(_0173_),
    .y(\DFF_22.D )
  );
  al_and3 _1621_ (
    .a(g109),
    .b(\DFF_323.Q ),
    .c(\DFF_320.Q ),
    .y(\DFF_21.D )
  );
  al_aoi21ttf _1622_ (
    .a(\DFF_22.D ),
    .b(\DFF_21.D ),
    .c(_0171_),
    .y(_0191_)
  );
  al_and3ftt _1623_ (
    .a(_0150_),
    .b(_0112_),
    .c(_0191_),
    .y(_0192_)
  );
  al_nand3 _1624_ (
    .a(\DFF_408.Q ),
    .b(_0056_),
    .c(_0040_),
    .y(_0193_)
  );
  al_nand3 _1625_ (
    .a(\DFF_52.Q ),
    .b(_0045_),
    .c(_0040_),
    .y(_0194_)
  );
  al_nand3 _1626_ (
    .a(g904),
    .b(_0050_),
    .c(_0040_),
    .y(_0195_)
  );
  al_aoi21ftf _1627_ (
    .a(_0025_),
    .b(g892),
    .c(_0195_),
    .y(_0196_)
  );
  al_and3 _1628_ (
    .a(_0193_),
    .b(_0194_),
    .c(_0196_),
    .y(_0197_)
  );
  al_nand3 _1629_ (
    .a(\DFF_198.Q ),
    .b(_0045_),
    .c(_0055_),
    .y(_0198_)
  );
  al_nand3 _1630_ (
    .a(\DFF_458.Q ),
    .b(_0056_),
    .c(_0055_),
    .y(_0199_)
  );
  al_nand3 _1631_ (
    .a(g1176),
    .b(_0050_),
    .c(_0055_),
    .y(_0200_)
  );
  al_aoi21ftf _1632_ (
    .a(_0118_),
    .b(g1200),
    .c(_0200_),
    .y(_0201_)
  );
  al_and3 _1633_ (
    .a(_0198_),
    .b(_0199_),
    .c(_0201_),
    .y(_0202_)
  );
  al_and3 _1634_ (
    .a(\DFF_528.Q ),
    .b(_0064_),
    .c(_0052_),
    .y(_0203_)
  );
  al_and3ftt _1635_ (
    .a(_0032_),
    .b(\DFF_501.Q ),
    .c(_0059_),
    .y(_0204_)
  );
  al_inv _1636_ (
    .a(\DFF_17.Q ),
    .y(_0205_)
  );
  al_inv _1637_ (
    .a(\DFF_164.Q ),
    .y(_0206_)
  );
  al_nand3fft _1638_ (
    .a(_0206_),
    .b(_0028_),
    .c(_0052_),
    .y(_0207_)
  );
  al_aoi21ftf _1639_ (
    .a(_0205_),
    .b(_0126_),
    .c(_0207_),
    .y(_0208_)
  );
  al_nand3fft _1640_ (
    .a(_0203_),
    .b(_0204_),
    .c(_0208_),
    .y(_0209_)
  );
  al_and3ftt _1641_ (
    .a(_0209_),
    .b(_0197_),
    .c(_0202_),
    .y(_0210_)
  );
  al_mux2l _1642_ (
    .a(_0041_),
    .b(_0068_),
    .s(\DFF_176.Q ),
    .y(_0211_)
  );
  al_nand3fft _1643_ (
    .a(\DFF_197.Q ),
    .b(_0041_),
    .c(_0062_),
    .y(_0212_)
  );
  al_or3fft _1644_ (
    .a(_0043_),
    .b(_0212_),
    .c(_0211_),
    .y(_0213_)
  );
  al_oai21ftt _1645_ (
    .a(g48),
    .b(g31),
    .c(\DFF_242.Q ),
    .y(_0214_)
  );
  al_nand3ftt _1646_ (
    .a(_0021_),
    .b(\DFF_340.Q ),
    .c(_0040_),
    .y(_0215_)
  );
  al_nand3ftt _1647_ (
    .a(_0019_),
    .b(\DFF_370.Q ),
    .c(_0059_),
    .y(_0216_)
  );
  al_nand3 _1648_ (
    .a(_0214_),
    .b(_0215_),
    .c(_0216_),
    .y(_0217_)
  );
  al_and3 _1649_ (
    .a(\DFF_514.Q ),
    .b(_0123_),
    .c(_0052_),
    .y(_0218_)
  );
  al_nand3 _1650_ (
    .a(\DFF_179.Q ),
    .b(_0063_),
    .c(_0062_),
    .y(_0219_)
  );
  al_nand3 _1651_ (
    .a(\DFF_456.Q ),
    .b(_0044_),
    .c(_0062_),
    .y(_0220_)
  );
  al_and3ftt _1652_ (
    .a(_0218_),
    .b(_0219_),
    .c(_0220_),
    .y(_0221_)
  );
  al_and3ftt _1653_ (
    .a(_0217_),
    .b(_0213_),
    .c(_0221_),
    .y(_0222_)
  );
  al_nand3 _1654_ (
    .a(_0222_),
    .b(_0120_),
    .c(_0210_),
    .y(\DFF_242.D )
  );
  al_or3fft _1655_ (
    .a(_0141_),
    .b(_0149_),
    .c(\DFF_242.D ),
    .y(_0223_)
  );
  al_ao21ttf _1656_ (
    .a(\DFF_228.D ),
    .b(\DFF_242.D ),
    .c(_0223_),
    .y(_0224_)
  );
  al_and3 _1657_ (
    .a(_0114_),
    .b(_0119_),
    .c(_0116_),
    .y(_0225_)
  );
  al_nand3 _1658_ (
    .a(g1197),
    .b(_0123_),
    .c(_0055_),
    .y(_0226_)
  );
  al_ao21ftf _1659_ (
    .a(_0029_),
    .b(g901),
    .c(_0226_),
    .y(_0227_)
  );
  al_nand3 _1660_ (
    .a(\DFF_425.Q ),
    .b(_0056_),
    .c(_0052_),
    .y(_0228_)
  );
  al_nand3 _1661_ (
    .a(\DFF_317.Q ),
    .b(_0056_),
    .c(_0040_),
    .y(_0229_)
  );
  al_or3fft _1662_ (
    .a(_0228_),
    .b(_0229_),
    .c(_0227_),
    .y(_0230_)
  );
  al_or3fft _1663_ (
    .a(g925),
    .b(_0036_),
    .c(_0018_),
    .y(_0231_)
  );
  al_aoi21ftf _1664_ (
    .a(_0031_),
    .b(\DFF_384.Q ),
    .c(_0231_),
    .y(_0232_)
  );
  al_aoi21ftf _1665_ (
    .a(_0172_),
    .b(\DFF_470.Q ),
    .c(_0232_),
    .y(_0233_)
  );
  al_aoi21ttf _1666_ (
    .a(\DFF_530.Q ),
    .b(_0092_),
    .c(_0233_),
    .y(_0234_)
  );
  al_nand3 _1667_ (
    .a(g889),
    .b(_0024_),
    .c(_0040_),
    .y(_0235_)
  );
  al_nand3 _1668_ (
    .a(g1173),
    .b(_0050_),
    .c(_0055_),
    .y(_0236_)
  );
  al_and3 _1669_ (
    .a(\DFF_14.Q ),
    .b(_0045_),
    .c(_0040_),
    .y(_0237_)
  );
  al_and3ftt _1670_ (
    .a(_0237_),
    .b(_0235_),
    .c(_0236_),
    .y(_0238_)
  );
  al_nand3 _1671_ (
    .a(\DFF_29.Q ),
    .b(_0064_),
    .c(_0052_),
    .y(_0239_)
  );
  al_aoi21ttf _1672_ (
    .a(\DFF_83.Q ),
    .b(_0022_),
    .c(_0239_),
    .y(_0240_)
  );
  al_nand3 _1673_ (
    .a(\DFF_448.Q ),
    .b(_0056_),
    .c(_0055_),
    .y(_0241_)
  );
  al_ao21ftf _1674_ (
    .a(_0075_),
    .b(\DFF_463.Q ),
    .c(_0241_),
    .y(_0242_)
  );
  al_and3ftt _1675_ (
    .a(_0242_),
    .b(_0240_),
    .c(_0238_),
    .y(_0243_)
  );
  al_and3ftt _1676_ (
    .a(_0230_),
    .b(_0234_),
    .c(_0243_),
    .y(_0244_)
  );
  al_mux2l _1677_ (
    .a(_0041_),
    .b(_0068_),
    .s(\DFF_485.Q ),
    .y(_0245_)
  );
  al_nand3fft _1678_ (
    .a(\DFF_251.Q ),
    .b(_0041_),
    .c(_0062_),
    .y(_0246_)
  );
  al_or3fft _1679_ (
    .a(_0043_),
    .b(_0246_),
    .c(_0245_),
    .y(_0247_)
  );
  al_and3ftt _1680_ (
    .a(_0032_),
    .b(_0063_),
    .c(_0052_),
    .y(_0248_)
  );
  al_nand3 _1681_ (
    .a(\DFF_140.Q ),
    .b(_0049_),
    .c(_0126_),
    .y(_0249_)
  );
  al_aoi21ttf _1682_ (
    .a(\DFF_531.Q ),
    .b(_0248_),
    .c(_0249_),
    .y(_0250_)
  );
  al_nand3ftt _1683_ (
    .a(_0032_),
    .b(\DFF_388.Q ),
    .c(_0059_),
    .y(_0251_)
  );
  al_ao21ftf _1684_ (
    .a(_0106_),
    .b(\DFF_505.Q ),
    .c(_0251_),
    .y(_0252_)
  );
  al_and3ftt _1685_ (
    .a(_0252_),
    .b(_0247_),
    .c(_0250_),
    .y(_0253_)
  );
  al_nand3 _1686_ (
    .a(_0253_),
    .b(_0120_),
    .c(_0244_),
    .y(\DFF_384.D )
  );
  al_nand3 _1687_ (
    .a(g1194),
    .b(_0123_),
    .c(_0055_),
    .y(_0254_)
  );
  al_ao21ttf _1688_ (
    .a(\DFF_243.Q ),
    .b(_0022_),
    .c(_0254_),
    .y(_0255_)
  );
  al_nand3 _1689_ (
    .a(g898),
    .b(_0050_),
    .c(_0040_),
    .y(_0256_)
  );
  al_ao21ftf _1690_ (
    .a(_0172_),
    .b(\DFF_344.Q ),
    .c(_0256_),
    .y(_0257_)
  );
  al_nand3 _1691_ (
    .a(\DFF_391.Q ),
    .b(_0050_),
    .c(_0052_),
    .y(_0258_)
  );
  al_nand3 _1692_ (
    .a(\DFF_453.Q ),
    .b(_0123_),
    .c(_0052_),
    .y(_0259_)
  );
  al_nor3fft _1693_ (
    .a(g922),
    .b(_0036_),
    .c(_0018_),
    .y(_0260_)
  );
  al_oa21ftt _1694_ (
    .a(g48),
    .b(g31),
    .c(\DFF_168.Q ),
    .y(_0261_)
  );
  al_oai21ftf _1695_ (
    .a(_0036_),
    .b(_0011_),
    .c(_0261_),
    .y(_0262_)
  );
  al_nor2 _1696_ (
    .a(_0260_),
    .b(_0262_),
    .y(_0263_)
  );
  al_and3 _1697_ (
    .a(_0258_),
    .b(_0259_),
    .c(_0263_),
    .y(_0264_)
  );
  al_nand3fft _1698_ (
    .a(_0255_),
    .b(_0257_),
    .c(_0264_),
    .y(_0265_)
  );
  al_nand3 _1699_ (
    .a(\DFF_342.Q ),
    .b(_0056_),
    .c(_0055_),
    .y(_0266_)
  );
  al_ao21ftf _1700_ (
    .a(_0103_),
    .b(\DFF_294.Q ),
    .c(_0266_),
    .y(_0267_)
  );
  al_nand3 _1701_ (
    .a(g1170),
    .b(_0050_),
    .c(_0055_),
    .y(_0268_)
  );
  al_ao21ftf _1702_ (
    .a(_0025_),
    .b(g886),
    .c(_0268_),
    .y(_0269_)
  );
  al_inv _1703_ (
    .a(\DFF_520.Q ),
    .y(_0270_)
  );
  al_nand3 _1704_ (
    .a(\DFF_371.Q ),
    .b(_0056_),
    .c(_0052_),
    .y(_0271_)
  );
  al_aoi21ftf _1705_ (
    .a(_0270_),
    .b(_0126_),
    .c(_0271_),
    .y(_0272_)
  );
  al_nand3 _1706_ (
    .a(\DFF_365.Q ),
    .b(_0056_),
    .c(_0040_),
    .y(_0273_)
  );
  al_nand3 _1707_ (
    .a(\DFF_4.Q ),
    .b(_0064_),
    .c(_0052_),
    .y(_0274_)
  );
  al_and3 _1708_ (
    .a(_0273_),
    .b(_0274_),
    .c(_0272_),
    .y(_0275_)
  );
  al_nand3fft _1709_ (
    .a(_0267_),
    .b(_0269_),
    .c(_0275_),
    .y(_0276_)
  );
  al_mux2l _1710_ (
    .a(_0041_),
    .b(_0068_),
    .s(\DFF_386.Q ),
    .y(_0277_)
  );
  al_nand3fft _1711_ (
    .a(\DFF_259.Q ),
    .b(_0041_),
    .c(_0062_),
    .y(_0278_)
  );
  al_or3fft _1712_ (
    .a(_0043_),
    .b(_0278_),
    .c(_0277_),
    .y(_0279_)
  );
  al_nand3ftt _1713_ (
    .a(_0019_),
    .b(\DFF_120.Q ),
    .c(_0059_),
    .y(_0280_)
  );
  al_and3 _1714_ (
    .a(\DFF_380.Q ),
    .b(_0063_),
    .c(_0062_),
    .y(_0281_)
  );
  al_aoi21 _1715_ (
    .a(\DFF_9.Q ),
    .b(_0072_),
    .c(_0281_),
    .y(_0282_)
  );
  al_nand3 _1716_ (
    .a(_0280_),
    .b(_0279_),
    .c(_0282_),
    .y(_0283_)
  );
  al_or3 _1717_ (
    .a(_0283_),
    .b(_0265_),
    .c(_0276_),
    .y(_0284_)
  );
  al_oai21 _1718_ (
    .a(_0225_),
    .b(_0284_),
    .c(\DFF_384.D ),
    .y(_0285_)
  );
  al_ao21ttf _1719_ (
    .a(_0123_),
    .b(_0052_),
    .c(\DFF_391.Q ),
    .y(_0286_)
  );
  al_ao21 _1720_ (
    .a(_0259_),
    .b(_0286_),
    .c(_0053_),
    .y(_0287_)
  );
  al_ao21ftf _1721_ (
    .a(_0270_),
    .b(_0126_),
    .c(_0280_),
    .y(_0288_)
  );
  al_aoi21 _1722_ (
    .a(\DFF_4.Q ),
    .b(_0065_),
    .c(_0281_),
    .y(_0289_)
  );
  al_nand3ftt _1723_ (
    .a(_0288_),
    .b(_0289_),
    .c(_0287_),
    .y(_0290_)
  );
  al_nand3ftt _1724_ (
    .a(_0021_),
    .b(\DFF_243.Q ),
    .c(_0040_),
    .y(_0291_)
  );
  al_and3 _1725_ (
    .a(\DFF_294.Q ),
    .b(_0045_),
    .c(_0040_),
    .y(_0292_)
  );
  al_and3ftt _1726_ (
    .a(_0292_),
    .b(_0291_),
    .c(_0256_),
    .y(_0293_)
  );
  al_aoi21ftf _1727_ (
    .a(_0172_),
    .b(\DFF_344.Q ),
    .c(_0254_),
    .y(_0294_)
  );
  al_ao21ftf _1728_ (
    .a(_0025_),
    .b(g886),
    .c(_0273_),
    .y(_0295_)
  );
  al_and3ftt _1729_ (
    .a(_0295_),
    .b(_0294_),
    .c(_0293_),
    .y(_0296_)
  );
  al_nand3ftt _1730_ (
    .a(_0032_),
    .b(\DFF_9.Q ),
    .c(_0059_),
    .y(_0297_)
  );
  al_ao21ftf _1731_ (
    .a(_0049_),
    .b(\DFF_371.Q ),
    .c(_0297_),
    .y(_0298_)
  );
  al_nand3fft _1732_ (
    .a(_0260_),
    .b(_0262_),
    .c(_0268_),
    .y(_0299_)
  );
  al_nor3ftt _1733_ (
    .a(_0266_),
    .b(_0299_),
    .c(_0298_),
    .y(_0300_)
  );
  al_and3 _1734_ (
    .a(_0279_),
    .b(_0300_),
    .c(_0296_),
    .y(_0301_)
  );
  al_nand3fft _1735_ (
    .a(_0290_),
    .b(_0225_),
    .c(_0301_),
    .y(\DFF_168.D )
  );
  al_or3fft _1736_ (
    .a(_0244_),
    .b(_0253_),
    .c(\DFF_168.D ),
    .y(_0302_)
  );
  al_or3fft _1737_ (
    .a(_0285_),
    .b(_0302_),
    .c(_0224_),
    .y(_0303_)
  );
  al_aoi21ttf _1738_ (
    .a(_0285_),
    .b(_0302_),
    .c(_0224_),
    .y(_0304_)
  );
  al_nand2ft _1739_ (
    .a(_0304_),
    .b(_0303_),
    .y(_0305_)
  );
  al_and2 _1740_ (
    .a(\DFF_116.D ),
    .b(\DFF_350.D ),
    .y(_0306_)
  );
  al_nor2 _1741_ (
    .a(\DFF_116.D ),
    .b(\DFF_350.D ),
    .y(_0307_)
  );
  al_or2 _1742_ (
    .a(_0307_),
    .b(_0306_),
    .y(_0308_)
  );
  al_or2 _1743_ (
    .a(\DFF_319.D ),
    .b(\DFF_22.D ),
    .y(_0309_)
  );
  al_and2 _1744_ (
    .a(\DFF_319.D ),
    .b(\DFF_22.D ),
    .y(_0310_)
  );
  al_ao21ftt _1745_ (
    .a(_0310_),
    .b(_0309_),
    .c(_0308_),
    .y(_0311_)
  );
  al_and3ftt _1746_ (
    .a(_0310_),
    .b(_0309_),
    .c(_0308_),
    .y(_0312_)
  );
  al_ao21ftt _1747_ (
    .a(_0312_),
    .b(_0311_),
    .c(_0305_),
    .y(_0313_)
  );
  al_nand3ftt _1748_ (
    .a(_0312_),
    .b(_0311_),
    .c(_0305_),
    .y(_0314_)
  );
  al_and2 _1749_ (
    .a(_0314_),
    .b(_0313_),
    .y(_0315_)
  );
  al_oa21ttf _1750_ (
    .a(\DFF_92.Q ),
    .b(_0031_),
    .c(_0315_),
    .y(_0316_)
  );
  al_nand3fft _1751_ (
    .a(\DFF_92.Q ),
    .b(_0031_),
    .c(_0315_),
    .y(_0317_)
  );
  al_nor3fft _1752_ (
    .a(_0192_),
    .b(_0317_),
    .c(_0316_),
    .y(_0318_)
  );
  al_oai21ftf _1753_ (
    .a(_0317_),
    .b(_0316_),
    .c(_0192_),
    .y(_0319_)
  );
  al_nand2ft _1754_ (
    .a(_0318_),
    .b(_0319_),
    .y(g11163)
  );
  al_and3 _1755_ (
    .a(\DFF_294.Q ),
    .b(\DFF_52.Q ),
    .c(\DFF_14.Q ),
    .y(_0320_)
  );
  al_and2 _1756_ (
    .a(\DFF_293.Q ),
    .b(_0320_),
    .y(\DFF_53.D )
  );
  al_inv _1757_ (
    .a(\DFF_233.Q ),
    .y(g5816)
  );
  al_or3 _1758_ (
    .a(g41),
    .b(g42),
    .c(_0014_),
    .y(_0321_)
  );
  al_or3 _1759_ (
    .a(_0026_),
    .b(_0018_),
    .c(_0321_),
    .y(\DFF_357.D )
  );
  al_nand3ftt _1760_ (
    .a(\DFF_121.Q ),
    .b(g109),
    .c(\DFF_291.Q ),
    .y(_0322_)
  );
  al_aoi21ttf _1761_ (
    .a(g881),
    .b(g109),
    .c(_0322_),
    .y(\DFF_71.D )
  );
  al_nor2 _1762_ (
    .a(\DFF_323.Q ),
    .b(\DFF_25.Q ),
    .y(\DFF_320.D )
  );
  al_and2ft _1763_ (
    .a(g750),
    .b(\DFF_304.Q ),
    .y(g4171)
  );
  al_or3 _1764_ (
    .a(_0026_),
    .b(_0018_),
    .c(_0015_),
    .y(\DFF_398.D )
  );
  al_nand3fft _1765_ (
    .a(_0151_),
    .b(\DFF_412.Q ),
    .c(\DFF_228.D ),
    .y(_0323_)
  );
  al_ao21ttf _1766_ (
    .a(g109),
    .b(\DFF_228.D ),
    .c(\DFF_412.Q ),
    .y(_0324_)
  );
  al_and2 _1767_ (
    .a(_0323_),
    .b(_0324_),
    .y(_0325_)
  );
  al_nand3fft _1768_ (
    .a(_0151_),
    .b(\DFF_338.Q ),
    .c(\DFF_384.D ),
    .y(_0326_)
  );
  al_ao21ttf _1769_ (
    .a(g109),
    .b(\DFF_384.D ),
    .c(\DFF_338.Q ),
    .y(_0327_)
  );
  al_inv _1770_ (
    .a(\DFF_343.Q ),
    .y(_0328_)
  );
  al_ao21 _1771_ (
    .a(g109),
    .b(\DFF_116.D ),
    .c(_0328_),
    .y(_0329_)
  );
  al_and3 _1772_ (
    .a(_0329_),
    .b(_0326_),
    .c(_0327_),
    .y(_0330_)
  );
  al_nor2 _1773_ (
    .a(\DFF_248.Q ),
    .b(\DFF_55.Q ),
    .y(_0331_)
  );
  al_ao21 _1774_ (
    .a(g109),
    .b(\DFF_168.D ),
    .c(_0331_),
    .y(_0332_)
  );
  al_and2 _1775_ (
    .a(\DFF_248.Q ),
    .b(\DFF_55.Q ),
    .y(_0333_)
  );
  al_nand3ftt _1776_ (
    .a(_0333_),
    .b(g109),
    .c(\DFF_168.D ),
    .y(_0334_)
  );
  al_nand3fft _1777_ (
    .a(_0151_),
    .b(\DFF_433.Q ),
    .c(\DFF_350.D ),
    .y(_0335_)
  );
  al_nand3 _1778_ (
    .a(_0335_),
    .b(_0334_),
    .c(_0332_),
    .y(_0336_)
  );
  al_and3ftt _1779_ (
    .a(_0336_),
    .b(_0325_),
    .c(_0330_),
    .y(_0337_)
  );
  al_and3 _1780_ (
    .a(g109),
    .b(\DFF_405.Q ),
    .c(\DFF_22.D ),
    .y(_0338_)
  );
  al_ao21 _1781_ (
    .a(g109),
    .b(\DFF_22.D ),
    .c(\DFF_405.Q ),
    .y(_0339_)
  );
  al_nand2ft _1782_ (
    .a(_0338_),
    .b(_0339_),
    .y(_0340_)
  );
  al_inv _1783_ (
    .a(\DFF_367.Q ),
    .y(_0341_)
  );
  al_and3 _1784_ (
    .a(g109),
    .b(_0341_),
    .c(\DFF_319.D ),
    .y(_0342_)
  );
  al_ao21 _1785_ (
    .a(g109),
    .b(\DFF_319.D ),
    .c(_0341_),
    .y(_0343_)
  );
  al_nand3fft _1786_ (
    .a(_0151_),
    .b(\DFF_343.Q ),
    .c(\DFF_116.D ),
    .y(_0344_)
  );
  al_and3ftt _1787_ (
    .a(_0342_),
    .b(_0343_),
    .c(_0344_),
    .y(_0345_)
  );
  al_ao21 _1788_ (
    .a(g109),
    .b(\DFF_242.D ),
    .c(\DFF_309.Q ),
    .y(_0346_)
  );
  al_and3 _1789_ (
    .a(g109),
    .b(\DFF_309.Q ),
    .c(\DFF_242.D ),
    .y(_0347_)
  );
  al_ao21ttf _1790_ (
    .a(g109),
    .b(\DFF_350.D ),
    .c(\DFF_433.Q ),
    .y(_0348_)
  );
  al_aoi21ftf _1791_ (
    .a(_0347_),
    .b(_0346_),
    .c(_0348_),
    .y(_0349_)
  );
  al_and3 _1792_ (
    .a(_0345_),
    .b(_0340_),
    .c(_0349_),
    .y(_0350_)
  );
  al_or3 _1793_ (
    .a(\DFF_309.Q ),
    .b(\DFF_405.Q ),
    .c(\DFF_343.Q ),
    .y(_0351_)
  );
  al_nor2 _1794_ (
    .a(\DFF_433.Q ),
    .b(\DFF_338.Q ),
    .y(_0352_)
  );
  al_nand3fft _1795_ (
    .a(\DFF_412.Q ),
    .b(\DFF_367.Q ),
    .c(_0352_),
    .y(_0353_)
  );
  al_and3fft _1796_ (
    .a(_0351_),
    .b(_0353_),
    .c(_0331_),
    .y(_0354_)
  );
  al_ao21ttf _1797_ (
    .a(_0350_),
    .b(_0337_),
    .c(_0354_),
    .y(_0355_)
  );
  al_and3 _1798_ (
    .a(\DFF_19.Q ),
    .b(\DFF_207.Q ),
    .c(\DFF_409.Q ),
    .y(_0356_)
  );
  al_and2 _1799_ (
    .a(\DFF_483.Q ),
    .b(_0356_),
    .y(_0357_)
  );
  al_inv _1800_ (
    .a(\DFF_265.Q ),
    .y(_0358_)
  );
  al_inv _1801_ (
    .a(\DFF_492.Q ),
    .y(_0359_)
  );
  al_nor2 _1802_ (
    .a(\DFF_406.Q ),
    .b(\DFF_114.Q ),
    .y(_0360_)
  );
  al_nand3fft _1803_ (
    .a(\DFF_124.Q ),
    .b(\DFF_177.Q ),
    .c(_0360_),
    .y(_0361_)
  );
  al_or3 _1804_ (
    .a(\DFF_378.Q ),
    .b(\DFF_3.Q ),
    .c(_0361_),
    .y(_0362_)
  );
  al_or3 _1805_ (
    .a(\DFF_419.Q ),
    .b(\DFF_368.Q ),
    .c(\DFF_491.Q ),
    .y(_0363_)
  );
  al_nor2 _1806_ (
    .a(\DFF_217.Q ),
    .b(\DFF_171.Q ),
    .y(_0364_)
  );
  al_and3fft _1807_ (
    .a(\DFF_204.Q ),
    .b(\DFF_394.Q ),
    .c(_0364_),
    .y(_0365_)
  );
  al_or3ftt _1808_ (
    .a(_0365_),
    .b(_0363_),
    .c(_0362_),
    .y(_0366_)
  );
  al_nand3fft _1809_ (
    .a(\DFF_512.Q ),
    .b(\DFF_492.Q ),
    .c(_0366_),
    .y(_0367_)
  );
  al_ao21ftf _1810_ (
    .a(_0359_),
    .b(\DFF_512.Q ),
    .c(_0367_),
    .y(_0368_)
  );
  al_nand2ft _1811_ (
    .a(\DFF_124.Q ),
    .b(\DFF_41.Q ),
    .y(_0369_)
  );
  al_nand2ft _1812_ (
    .a(\DFF_41.Q ),
    .b(\DFF_124.Q ),
    .y(_0370_)
  );
  al_nand2ft _1813_ (
    .a(\DFF_478.Q ),
    .b(\DFF_394.Q ),
    .y(_0371_)
  );
  al_nand2ft _1814_ (
    .a(\DFF_394.Q ),
    .b(\DFF_478.Q ),
    .y(_0372_)
  );
  al_nand2ft _1815_ (
    .a(\DFF_406.Q ),
    .b(\DFF_2.Q ),
    .y(_0373_)
  );
  al_aoi21ftf _1816_ (
    .a(\DFF_65.Q ),
    .b(\DFF_177.Q ),
    .c(_0373_),
    .y(_0374_)
  );
  al_and3 _1817_ (
    .a(_0371_),
    .b(_0372_),
    .c(_0374_),
    .y(_0375_)
  );
  al_and3 _1818_ (
    .a(_0369_),
    .b(_0370_),
    .c(_0375_),
    .y(_0376_)
  );
  al_nand2ft _1819_ (
    .a(\DFF_177.Q ),
    .b(\DFF_65.Q ),
    .y(_0377_)
  );
  al_nand2ft _1820_ (
    .a(\DFF_419.Q ),
    .b(\DFF_239.Q ),
    .y(_0378_)
  );
  al_nand2ft _1821_ (
    .a(\DFF_467.Q ),
    .b(\DFF_114.Q ),
    .y(_0379_)
  );
  al_aoi21ftf _1822_ (
    .a(\DFF_217.Q ),
    .b(\DFF_225.Q ),
    .c(_0379_),
    .y(_0380_)
  );
  al_and3 _1823_ (
    .a(_0377_),
    .b(_0378_),
    .c(_0380_),
    .y(_0381_)
  );
  al_nand2ft _1824_ (
    .a(\DFF_2.Q ),
    .b(\DFF_406.Q ),
    .y(_0382_)
  );
  al_aoi21ftf _1825_ (
    .a(\DFF_225.Q ),
    .b(\DFF_217.Q ),
    .c(_0382_),
    .y(_0383_)
  );
  al_nand2ft _1826_ (
    .a(\DFF_183.Q ),
    .b(\DFF_204.Q ),
    .y(_0384_)
  );
  al_aoi21ftf _1827_ (
    .a(\DFF_114.Q ),
    .b(\DFF_467.Q ),
    .c(_0384_),
    .y(_0385_)
  );
  al_nand2ft _1828_ (
    .a(\DFF_175.Q ),
    .b(\DFF_491.Q ),
    .y(_0386_)
  );
  al_aoi21ftf _1829_ (
    .a(\DFF_239.Q ),
    .b(\DFF_419.Q ),
    .c(_0386_),
    .y(_0387_)
  );
  al_nand2ft _1830_ (
    .a(\DFF_491.Q ),
    .b(\DFF_175.Q ),
    .y(_0388_)
  );
  al_nand2ft _1831_ (
    .a(\DFF_204.Q ),
    .b(\DFF_183.Q ),
    .y(_0389_)
  );
  al_and3 _1832_ (
    .a(_0388_),
    .b(_0389_),
    .c(_0387_),
    .y(_0390_)
  );
  al_and3 _1833_ (
    .a(_0383_),
    .b(_0385_),
    .c(_0390_),
    .y(_0391_)
  );
  al_nand3 _1834_ (
    .a(_0381_),
    .b(_0391_),
    .c(_0376_),
    .y(_0392_)
  );
  al_mux2l _1835_ (
    .a(\DFF_265.Q ),
    .b(_0368_),
    .s(_0392_),
    .y(_0393_)
  );
  al_ao21ftf _1836_ (
    .a(_0358_),
    .b(_0368_),
    .c(_0393_),
    .y(_0394_)
  );
  al_and3 _1837_ (
    .a(_0357_),
    .b(_0394_),
    .c(_0355_),
    .y(\DFF_37.D )
  );
  al_nand2ft _1838_ (
    .a(\DFF_275.Q ),
    .b(g1700),
    .y(\DFF_471.D )
  );
  al_mux2h _1839_ (
    .a(\DFF_77.Q ),
    .b(\DFF_276.Q ),
    .s(g1700),
    .y(_0395_)
  );
  al_aoi21ttf _1840_ (
    .a(\DFF_77.Q ),
    .b(\DFF_276.Q ),
    .c(_0395_),
    .y(\DFF_276.D )
  );
  al_nor2 _1841_ (
    .a(\DFF_362.Q ),
    .b(\DFF_310.Q ),
    .y(_0396_)
  );
  al_mux2l _1842_ (
    .a(\DFF_135.Q ),
    .b(_0396_),
    .s(\DFF_358.Q ),
    .y(\DFF_262.D )
  );
  al_or3 _1843_ (
    .a(g46),
    .b(_0011_),
    .c(_0321_),
    .y(\DFF_526.D )
  );
  al_inv _1844_ (
    .a(\DFF_413.Q ),
    .y(_0397_)
  );
  al_or3 _1845_ (
    .a(g46),
    .b(_0018_),
    .c(_0015_),
    .y(_0398_)
  );
  al_or2ft _1846_ (
    .a(_0398_),
    .b(\DFF_22.D ),
    .y(_0399_)
  );
  al_nand3 _1847_ (
    .a(\DFF_234.Q ),
    .b(_0397_),
    .c(_0399_),
    .y(_0400_)
  );
  al_ao21 _1848_ (
    .a(\DFF_234.Q ),
    .b(_0399_),
    .c(_0397_),
    .y(_0401_)
  );
  al_or3 _1849_ (
    .a(\DFF_202.Q ),
    .b(\DFF_510.Q ),
    .c(\DFF_250.Q ),
    .y(_0402_)
  );
  al_nor2 _1850_ (
    .a(\DFF_486.Q ),
    .b(\DFF_401.Q ),
    .y(_0403_)
  );
  al_nand3fft _1851_ (
    .a(\DFF_231.Q ),
    .b(\DFF_355.Q ),
    .c(_0403_),
    .y(_0404_)
  );
  al_nor2 _1852_ (
    .a(\DFF_334.Q ),
    .b(\DFF_498.Q ),
    .y(_0405_)
  );
  al_or2 _1853_ (
    .a(\DFF_480.Q ),
    .b(\DFF_322.Q ),
    .y(_0406_)
  );
  al_or3 _1854_ (
    .a(\DFF_58.Q ),
    .b(\DFF_61.Q ),
    .c(\DFF_442.Q ),
    .y(_0407_)
  );
  al_and3fft _1855_ (
    .a(_0406_),
    .b(_0407_),
    .c(_0405_),
    .y(_0408_)
  );
  al_nand3fft _1856_ (
    .a(_0402_),
    .b(_0404_),
    .c(_0408_),
    .y(_0409_)
  );
  al_and2 _1857_ (
    .a(\DFF_361.Q ),
    .b(\DFF_418.Q ),
    .y(_0410_)
  );
  al_nand3 _1858_ (
    .a(\DFF_28.Q ),
    .b(\DFF_119.Q ),
    .c(_0410_),
    .y(_0411_)
  );
  al_nand2 _1859_ (
    .a(\DFF_486.Q ),
    .b(\DFF_401.Q ),
    .y(_0412_)
  );
  al_ao21ftt _1860_ (
    .a(_0403_),
    .b(_0412_),
    .c(_0411_),
    .y(_0413_)
  );
  al_oai21ttf _1861_ (
    .a(\DFF_32.Q ),
    .b(_0409_),
    .c(_0413_),
    .y(_0414_)
  );
  al_ao21ttf _1862_ (
    .a(_0400_),
    .b(_0401_),
    .c(_0414_),
    .y(_0415_)
  );
  al_nand2ft _1863_ (
    .a(_0411_),
    .b(_0414_),
    .y(_0416_)
  );
  al_nand3 _1864_ (
    .a(_0416_),
    .b(_0400_),
    .c(_0401_),
    .y(_0417_)
  );
  al_and2ft _1865_ (
    .a(\DFF_334.Q ),
    .b(\DFF_428.Q ),
    .y(_0418_)
  );
  al_and2ft _1866_ (
    .a(\DFF_428.Q ),
    .b(\DFF_334.Q ),
    .y(_0419_)
  );
  al_nand2ft _1867_ (
    .a(\DFF_442.Q ),
    .b(\DFF_87.Q ),
    .y(_0420_)
  );
  al_nand2ft _1868_ (
    .a(\DFF_87.Q ),
    .b(\DFF_442.Q ),
    .y(_0421_)
  );
  al_nand2ft _1869_ (
    .a(\DFF_480.Q ),
    .b(\DFF_515.Q ),
    .y(_0422_)
  );
  al_aoi21ftf _1870_ (
    .a(\DFF_202.Q ),
    .b(\DFF_414.Q ),
    .c(_0422_),
    .y(_0423_)
  );
  al_and3 _1871_ (
    .a(_0420_),
    .b(_0421_),
    .c(_0423_),
    .y(_0424_)
  );
  al_nand3fft _1872_ (
    .a(_0418_),
    .b(_0419_),
    .c(_0424_),
    .y(_0425_)
  );
  al_and2ft _1873_ (
    .a(\DFF_355.Q ),
    .b(\DFF_108.Q ),
    .y(_0426_)
  );
  al_and2ft _1874_ (
    .a(\DFF_108.Q ),
    .b(\DFF_355.Q ),
    .y(_0427_)
  );
  al_nand2ft _1875_ (
    .a(\DFF_231.Q ),
    .b(\DFF_167.Q ),
    .y(_0428_)
  );
  al_aoi21ftf _1876_ (
    .a(\DFF_322.Q ),
    .b(\DFF_192.Q ),
    .c(_0428_),
    .y(_0429_)
  );
  al_nand3fft _1877_ (
    .a(_0426_),
    .b(_0427_),
    .c(_0429_),
    .y(_0430_)
  );
  al_nand2ft _1878_ (
    .a(\DFF_414.Q ),
    .b(\DFF_202.Q ),
    .y(_0431_)
  );
  al_aoi21ftf _1879_ (
    .a(\DFF_192.Q ),
    .b(\DFF_322.Q ),
    .c(_0431_),
    .y(_0432_)
  );
  al_nand2ft _1880_ (
    .a(\DFF_167.Q ),
    .b(\DFF_231.Q ),
    .y(_0433_)
  );
  al_aoi21ftf _1881_ (
    .a(\DFF_510.Q ),
    .b(\DFF_497.Q ),
    .c(_0433_),
    .y(_0434_)
  );
  al_nand2ft _1882_ (
    .a(\DFF_115.Q ),
    .b(\DFF_58.Q ),
    .y(_0435_)
  );
  al_nand2ft _1883_ (
    .a(\DFF_58.Q ),
    .b(\DFF_115.Q ),
    .y(_0436_)
  );
  al_nand2ft _1884_ (
    .a(\DFF_515.Q ),
    .b(\DFF_480.Q ),
    .y(_0437_)
  );
  al_aoi21ftf _1885_ (
    .a(\DFF_497.Q ),
    .b(\DFF_510.Q ),
    .c(_0437_),
    .y(_0438_)
  );
  al_and3 _1886_ (
    .a(_0435_),
    .b(_0436_),
    .c(_0438_),
    .y(_0439_)
  );
  al_and3 _1887_ (
    .a(_0432_),
    .b(_0434_),
    .c(_0439_),
    .y(_0440_)
  );
  al_nand3fft _1888_ (
    .a(_0430_),
    .b(_0425_),
    .c(_0440_),
    .y(_0441_)
  );
  al_ao21 _1889_ (
    .a(_0417_),
    .b(_0415_),
    .c(_0441_),
    .y(_0442_)
  );
  al_or3 _1890_ (
    .a(g1696),
    .b(\DFF_174.Q ),
    .c(\DFF_372.Q ),
    .y(_0443_)
  );
  al_nor3fft _1891_ (
    .a(\DFF_0.Q ),
    .b(_0410_),
    .c(_0443_),
    .y(_0444_)
  );
  al_and3 _1892_ (
    .a(\DFF_28.Q ),
    .b(\DFF_119.Q ),
    .c(_0444_),
    .y(_0445_)
  );
  al_and2 _1893_ (
    .a(_0445_),
    .b(_0442_),
    .y(\DFF_335.D )
  );
  al_and3 _1894_ (
    .a(\DFF_344.Q ),
    .b(\DFF_198.Q ),
    .c(\DFF_470.Q ),
    .y(_0446_)
  );
  al_and2 _1895_ (
    .a(\DFF_506.Q ),
    .b(_0446_),
    .y(\DFF_328.D )
  );
  al_or3 _1896_ (
    .a(g41),
    .b(g31),
    .c(g30),
    .y(g9451)
  );
  al_or3 _1897_ (
    .a(g30),
    .b(_0009_),
    .c(\DFF_242.D ),
    .y(g10459)
  );
  al_and3 _1898_ (
    .a(\DFF_112.Q ),
    .b(\DFF_149.Q ),
    .c(\DFF_407.Q ),
    .y(_0447_)
  );
  al_and3 _1899_ (
    .a(\DFF_253.Q ),
    .b(\DFF_30.Q ),
    .c(_0447_),
    .y(_0448_)
  );
  al_and3 _1900_ (
    .a(\DFF_247.Q ),
    .b(\DFF_301.Q ),
    .c(_0448_),
    .y(_0449_)
  );
  al_nand3 _1901_ (
    .a(\DFF_434.Q ),
    .b(\DFF_38.Q ),
    .c(_0449_),
    .y(_0450_)
  );
  al_ao21 _1902_ (
    .a(\DFF_38.Q ),
    .b(_0449_),
    .c(\DFF_434.Q ),
    .y(_0451_)
  );
  al_and2ft _1903_ (
    .a(\DFF_54.Q ),
    .b(g109),
    .y(_0452_)
  );
  al_and3 _1904_ (
    .a(_0452_),
    .b(_0450_),
    .c(_0451_),
    .y(\DFF_434.D )
  );
  al_and2 _1905_ (
    .a(\DFF_331.Q ),
    .b(g109),
    .y(\DFF_487.D )
  );
  al_and2 _1906_ (
    .a(g109),
    .b(\DFF_525.Q ),
    .y(\DFF_525.D )
  );
  al_and3 _1907_ (
    .a(\DFF_227.Q ),
    .b(\DFF_389.Q ),
    .c(\DFF_429.Q ),
    .y(_0453_)
  );
  al_and2 _1908_ (
    .a(\DFF_127.Q ),
    .b(_0453_),
    .y(_0454_)
  );
  al_and3 _1909_ (
    .a(\DFF_304.Q ),
    .b(g109),
    .c(\DFF_89.Q ),
    .y(_0455_)
  );
  al_mux2h _1910_ (
    .a(\DFF_393.Q ),
    .b(_0454_),
    .s(_0455_),
    .y(_0456_)
  );
  al_aoi21ttf _1911_ (
    .a(\DFF_393.Q ),
    .b(_0454_),
    .c(_0456_),
    .y(\DFF_393.D )
  );
  al_and3fft _1912_ (
    .a(\DFF_141.Q ),
    .b(\DFF_18.Q ),
    .c(\DFF_352.Q ),
    .y(_0457_)
  );
  al_and3ftt _1913_ (
    .a(\DFF_223.Q ),
    .b(\DFF_455.Q ),
    .c(\DFF_297.Q ),
    .y(_0458_)
  );
  al_nand3ftt _1914_ (
    .a(\DFF_111.Q ),
    .b(_0458_),
    .c(_0457_),
    .y(_0459_)
  );
  al_nand3ftt _1915_ (
    .a(\DFF_302.Q ),
    .b(\DFF_369.Q ),
    .c(\DFF_297.Q ),
    .y(_0460_)
  );
  al_nand2ft _1916_ (
    .a(\DFF_297.Q ),
    .b(\DFF_302.Q ),
    .y(_0461_)
  );
  al_and3 _1917_ (
    .a(_0460_),
    .b(_0461_),
    .c(_0459_),
    .y(_0462_)
  );
  al_ao21 _1918_ (
    .a(\DFF_178.Q ),
    .b(_0017_),
    .c(_0458_),
    .y(_0463_)
  );
  al_and3ftt _1919_ (
    .a(\DFF_111.Q ),
    .b(_0457_),
    .c(_0463_),
    .y(_0464_)
  );
  al_inv _1920_ (
    .a(\DFF_212.Q ),
    .y(_0465_)
  );
  al_inv _1921_ (
    .a(\DFF_271.Q ),
    .y(_0466_)
  );
  al_inv _1922_ (
    .a(\DFF_300.Q ),
    .y(_0467_)
  );
  al_inv _1923_ (
    .a(\DFF_44.Q ),
    .y(_0468_)
  );
  al_inv _1924_ (
    .a(\DFF_354.Q ),
    .y(_0469_)
  );
  al_nand3fft _1925_ (
    .a(\DFF_369.Q ),
    .b(\DFF_297.Q ),
    .c(\DFF_302.Q ),
    .y(_0470_)
  );
  al_mux2l _1926_ (
    .a(\DFF_369.Q ),
    .b(\DFF_297.Q ),
    .s(\DFF_302.Q ),
    .y(_0471_)
  );
  al_oai21ftt _1927_ (
    .a(_0470_),
    .b(_0471_),
    .c(\DFF_449.Q ),
    .y(_0472_)
  );
  al_and3fft _1928_ (
    .a(_0469_),
    .b(_0472_),
    .c(\DFF_1.Q ),
    .y(_0473_)
  );
  al_and3 _1929_ (
    .a(\DFF_333.Q ),
    .b(\DFF_461.Q ),
    .c(_0473_),
    .y(_0474_)
  );
  al_nand3fft _1930_ (
    .a(_0467_),
    .b(_0468_),
    .c(_0474_),
    .y(_0475_)
  );
  al_mux2l _1931_ (
    .a(_0465_),
    .b(_0475_),
    .s(_0466_),
    .y(_0476_)
  );
  al_inv _1932_ (
    .a(\DFF_1.Q ),
    .y(_0477_)
  );
  al_and3fft _1933_ (
    .a(\DFF_449.Q ),
    .b(_0471_),
    .c(_0470_),
    .y(_0478_)
  );
  al_and3 _1934_ (
    .a(_0477_),
    .b(_0469_),
    .c(_0478_),
    .y(_0479_)
  );
  al_and3fft _1935_ (
    .a(\DFF_333.Q ),
    .b(\DFF_461.Q ),
    .c(_0479_),
    .y(_0480_)
  );
  al_nand3fft _1936_ (
    .a(\DFF_300.Q ),
    .b(\DFF_44.Q ),
    .c(_0480_),
    .y(_0481_)
  );
  al_mux2l _1937_ (
    .a(\DFF_212.Q ),
    .b(_0481_),
    .s(\DFF_271.Q ),
    .y(_0482_)
  );
  al_nor3ftt _1938_ (
    .a(_0464_),
    .b(_0482_),
    .c(_0476_),
    .y(_0483_)
  );
  al_nand3fft _1939_ (
    .a(_0016_),
    .b(_0462_),
    .c(_0483_),
    .y(_0484_)
  );
  al_ao21ftf _1940_ (
    .a(_0462_),
    .b(_0483_),
    .c(_0016_),
    .y(_0485_)
  );
  al_and3 _1941_ (
    .a(g18),
    .b(_0484_),
    .c(_0485_),
    .y(\DFF_297.D )
  );
  al_and2 _1942_ (
    .a(\DFF_33.Q ),
    .b(g109),
    .y(\DFF_88.D )
  );
  al_oa21ftt _1943_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_23.Q ),
    .y(\DFF_23.D )
  );
  al_or2 _1944_ (
    .a(g82),
    .b(\DFF_533.Q ),
    .y(g8340)
  );
  al_and2 _1945_ (
    .a(g109),
    .b(\DFF_97.Q ),
    .y(\DFF_201.D )
  );
  al_aoi21ftf _1946_ (
    .a(\DFF_436.Q ),
    .b(\DFF_71.D ),
    .c(g109),
    .y(_0486_)
  );
  al_and2 _1947_ (
    .a(\DFF_340.Q ),
    .b(_0486_),
    .y(\DFF_340.D )
  );
  al_inv _1948_ (
    .a(\DFF_128.Q ),
    .y(_0487_)
  );
  al_nand2 _1949_ (
    .a(\DFF_105.Q ),
    .b(g18),
    .y(_0488_)
  );
  al_inv _1950_ (
    .a(g18),
    .y(_0489_)
  );
  al_nor2 _1951_ (
    .a(\DFF_417.Q ),
    .b(\DFF_278.Q ),
    .y(_0490_)
  );
  al_and2 _1952_ (
    .a(\DFF_31.Q ),
    .b(\DFF_158.Q ),
    .y(_0491_)
  );
  al_nand3 _1953_ (
    .a(\DFF_457.Q ),
    .b(_0490_),
    .c(_0491_),
    .y(_0492_)
  );
  al_ao21 _1954_ (
    .a(_0490_),
    .b(_0491_),
    .c(\DFF_457.Q ),
    .y(_0493_)
  );
  al_nand3 _1955_ (
    .a(_0489_),
    .b(_0492_),
    .c(_0493_),
    .y(_0494_)
  );
  al_nand3 _1956_ (
    .a(_0487_),
    .b(_0488_),
    .c(_0494_),
    .y(_0495_)
  );
  al_ao21 _1957_ (
    .a(_0488_),
    .b(_0494_),
    .c(_0487_),
    .y(_0496_)
  );
  al_and3 _1958_ (
    .a(g109),
    .b(_0495_),
    .c(_0496_),
    .y(\DFF_109.D )
  );
  al_mux2h _1959_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .s(\DFF_241.Q ),
    .y(\DFF_241.D )
  );
  al_and2 _1960_ (
    .a(g109),
    .b(\DFF_366.Q ),
    .y(\DFF_366.D )
  );
  al_and2 _1961_ (
    .a(\DFF_327.Q ),
    .b(g109),
    .y(\DFF_331.D )
  );
  al_and2 _1962_ (
    .a(\DFF_487.Q ),
    .b(g109),
    .y(\DFF_5.D )
  );
  al_inv _1963_ (
    .a(\DFF_235.Q ),
    .y(_0497_)
  );
  al_nand2 _1964_ (
    .a(\DFF_331.Q ),
    .b(g18),
    .y(_0498_)
  );
  al_and3fft _1965_ (
    .a(\DFF_278.Q ),
    .b(\DFF_31.Q ),
    .c(\DFF_417.Q ),
    .y(_0499_)
  );
  al_ao21ttf _1966_ (
    .a(\DFF_158.Q ),
    .b(_0499_),
    .c(\DFF_366.Q ),
    .y(_0500_)
  );
  al_nand3ftt _1967_ (
    .a(\DFF_366.Q ),
    .b(\DFF_158.Q ),
    .c(_0499_),
    .y(_0501_)
  );
  al_ao21 _1968_ (
    .a(_0501_),
    .b(_0500_),
    .c(g18),
    .y(_0502_)
  );
  al_nand3 _1969_ (
    .a(_0497_),
    .b(_0498_),
    .c(_0502_),
    .y(_0503_)
  );
  al_ao21 _1970_ (
    .a(_0498_),
    .b(_0502_),
    .c(_0497_),
    .y(_0504_)
  );
  al_and3 _1971_ (
    .a(g109),
    .b(_0503_),
    .c(_0504_),
    .y(\DFF_415.D )
  );
  al_or2 _1972_ (
    .a(g82),
    .b(\DFF_49.Q ),
    .y(g8349)
  );
  al_and2 _1973_ (
    .a(g109),
    .b(\DFF_34.Q ),
    .y(\DFF_97.D )
  );
  al_mux2h _1974_ (
    .a(\DFF_289.Q ),
    .b(\DFF_452.Q ),
    .s(g109),
    .y(_0505_)
  );
  al_and2ft _1975_ (
    .a(\DFF_473.Q ),
    .b(_0505_),
    .y(\DFF_289.D )
  );
  al_nor2ft _1976_ (
    .a(\DFF_330.Q ),
    .b(\DFF_122.D ),
    .y(\DFF_252.D )
  );
  al_and2 _1977_ (
    .a(\DFF_184.Q ),
    .b(\DFF_393.Q ),
    .y(_0506_)
  );
  al_nand3 _1978_ (
    .a(\DFF_127.Q ),
    .b(_0453_),
    .c(_0506_),
    .y(_0507_)
  );
  al_or3fft _1979_ (
    .a(\DFF_99.Q ),
    .b(\DFF_387.Q ),
    .c(_0507_),
    .y(_0508_)
  );
  al_nand2ft _1980_ (
    .a(\DFF_347.Q ),
    .b(_0508_),
    .y(_0509_)
  );
  al_nand3 _1981_ (
    .a(\DFF_387.Q ),
    .b(_0506_),
    .c(_0454_),
    .y(_0510_)
  );
  al_or3fft _1982_ (
    .a(\DFF_99.Q ),
    .b(\DFF_347.Q ),
    .c(_0510_),
    .y(_0511_)
  );
  al_and3 _1983_ (
    .a(_0455_),
    .b(_0511_),
    .c(_0509_),
    .y(\DFF_347.D )
  );
  al_or3 _1984_ (
    .a(\DFF_455.Q ),
    .b(\DFF_297.Q ),
    .c(_0017_),
    .y(_0512_)
  );
  al_nor2ft _1985_ (
    .a(_0512_),
    .b(_0483_),
    .y(_0513_)
  );
  al_and3fft _1986_ (
    .a(\DFF_297.Q ),
    .b(\DFF_302.Q ),
    .c(\DFF_369.Q ),
    .y(_0514_)
  );
  al_or3 _1987_ (
    .a(\DFF_455.Q ),
    .b(\DFF_369.Q ),
    .c(\DFF_302.Q ),
    .y(_0515_)
  );
  al_oa21ttf _1988_ (
    .a(\DFF_297.Q ),
    .b(_0515_),
    .c(_0514_),
    .y(_0516_)
  );
  al_and2 _1989_ (
    .a(\DFF_369.Q ),
    .b(\DFF_297.Q ),
    .y(_0517_)
  );
  al_ao21ttf _1990_ (
    .a(\DFF_302.Q ),
    .b(_0517_),
    .c(_0470_),
    .y(_0518_)
  );
  al_aoi21ftt _1991_ (
    .a(_0518_),
    .b(_0516_),
    .c(_0513_),
    .y(_0519_)
  );
  al_mux2l _1992_ (
    .a(\DFF_369.Q ),
    .b(_0519_),
    .s(_0489_),
    .y(_0520_)
  );
  al_aoi21ttf _1993_ (
    .a(\DFF_369.Q ),
    .b(_0519_),
    .c(_0520_),
    .y(\DFF_369.D )
  );
  al_and2 _1994_ (
    .a(\DFF_303.Q ),
    .b(g109),
    .y(\DFF_142.D )
  );
  al_nand2 _1995_ (
    .a(\DFF_185.Q ),
    .b(g18),
    .y(_0521_)
  );
  al_and3fft _1996_ (
    .a(\DFF_417.Q ),
    .b(\DFF_31.Q ),
    .c(\DFF_278.Q ),
    .y(_0522_)
  );
  al_nand3ftt _1997_ (
    .a(\DFF_158.Q ),
    .b(\DFF_468.Q ),
    .c(_0522_),
    .y(_0523_)
  );
  al_ao21ftt _1998_ (
    .a(\DFF_158.Q ),
    .b(_0522_),
    .c(\DFF_468.Q ),
    .y(_0524_)
  );
  al_nand3 _1999_ (
    .a(_0489_),
    .b(_0523_),
    .c(_0524_),
    .y(_0525_)
  );
  al_aoi21 _2000_ (
    .a(_0521_),
    .b(_0525_),
    .c(\DFF_36.Q ),
    .y(_0526_)
  );
  al_and3 _2001_ (
    .a(\DFF_36.Q ),
    .b(_0521_),
    .c(_0525_),
    .y(_0527_)
  );
  al_mux2l _2002_ (
    .a(_0527_),
    .b(_0526_),
    .s(_0151_),
    .y(\DFF_503.D )
  );
  al_nand3 _2003_ (
    .a(\DFF_344.Q ),
    .b(_0445_),
    .c(_0442_),
    .y(_0528_)
  );
  al_inv _2004_ (
    .a(\DFF_470.Q ),
    .y(_0529_)
  );
  al_and2ft _2005_ (
    .a(\DFF_299.Q ),
    .b(g109),
    .y(_0530_)
  );
  al_or3 _2006_ (
    .a(_0000_),
    .b(_0113_),
    .c(_0530_),
    .y(_0531_)
  );
  al_aoi21ttf _2007_ (
    .a(_0529_),
    .b(_0528_),
    .c(_0531_),
    .y(_0532_)
  );
  al_aoi21ftf _2008_ (
    .a(_0528_),
    .b(\DFF_470.Q ),
    .c(_0532_),
    .y(\DFF_470.D )
  );
  al_and2 _2009_ (
    .a(\DFF_182.Q ),
    .b(g109),
    .y(\DFF_33.D )
  );
  al_nand3 _2010_ (
    .a(\DFF_294.Q ),
    .b(\DFF_14.Q ),
    .c(\DFF_37.D ),
    .y(_0533_)
  );
  al_nand2ft _2011_ (
    .a(\DFF_188.Q ),
    .b(g109),
    .y(_0534_)
  );
  al_nand3ftt _2012_ (
    .a(\DFF_93.Q ),
    .b(g109),
    .c(\DFF_53.Q ),
    .y(_0535_)
  );
  al_aoi21ttf _2013_ (
    .a(\DFF_37.Q ),
    .b(g109),
    .c(_0535_),
    .y(_0536_)
  );
  al_and2 _2014_ (
    .a(_0534_),
    .b(_0536_),
    .y(_0537_)
  );
  al_ao21 _2015_ (
    .a(\DFF_294.Q ),
    .b(\DFF_37.D ),
    .c(\DFF_14.Q ),
    .y(_0538_)
  );
  al_and3ftt _2016_ (
    .a(_0537_),
    .b(_0533_),
    .c(_0538_),
    .y(\DFF_14.D )
  );
  al_and2 _2017_ (
    .a(\DFF_296.Q ),
    .b(g109),
    .y(\DFF_220.D )
  );
  al_mux2l _2018_ (
    .a(_0225_),
    .b(_0284_),
    .s(_0151_),
    .y(_0539_)
  );
  al_and2ft _2019_ (
    .a(_0322_),
    .b(\DFF_242.D ),
    .y(_0540_)
  );
  al_aoi21 _2020_ (
    .a(g877),
    .b(_0539_),
    .c(_0540_),
    .y(_0541_)
  );
  al_nand2ft _2021_ (
    .a(_0535_),
    .b(\DFF_350.D ),
    .y(_0542_)
  );
  al_nand3 _2022_ (
    .a(\DFF_37.Q ),
    .b(g109),
    .c(\DFF_228.D ),
    .y(_0543_)
  );
  al_nand3 _2023_ (
    .a(g881),
    .b(g109),
    .c(\DFF_384.D ),
    .y(_0544_)
  );
  al_and3 _2024_ (
    .a(_0542_),
    .b(_0543_),
    .c(_0544_),
    .y(_0545_)
  );
  al_and2 _2025_ (
    .a(_0541_),
    .b(_0545_),
    .y(g10628)
  );
  al_and3 _2026_ (
    .a(\DFF_12.Q ),
    .b(\DFF_255.Q ),
    .c(\DFF_264.Q ),
    .y(_0546_)
  );
  al_inv _2027_ (
    .a(_0546_),
    .y(_0547_)
  );
  al_ao21ftf _2028_ (
    .a(_0547_),
    .b(\DFF_152.Q ),
    .c(_0355_),
    .y(_0548_)
  );
  al_inv _2029_ (
    .a(\DFF_264.Q ),
    .y(_0549_)
  );
  al_nand2ft _2030_ (
    .a(\DFF_441.Q ),
    .b(g109),
    .y(_0550_)
  );
  al_aoi21 _2031_ (
    .a(_0549_),
    .b(_0548_),
    .c(_0550_),
    .y(_0551_)
  );
  al_aoi21ftf _2032_ (
    .a(_0548_),
    .b(\DFF_264.Q ),
    .c(_0551_),
    .y(\DFF_264.D )
  );
  al_or2 _2033_ (
    .a(g82),
    .b(\DFF_513.Q ),
    .y(g8328)
  );
  al_and2 _2034_ (
    .a(g109),
    .b(\DFF_240.Q ),
    .y(\DFF_240.D )
  );
  al_aoi21 _2035_ (
    .a(\DFF_227.Q ),
    .b(\DFF_429.Q ),
    .c(\DFF_389.Q ),
    .y(_0552_)
  );
  al_and3fft _2036_ (
    .a(_0552_),
    .b(_0453_),
    .c(_0455_),
    .y(\DFF_389.D )
  );
  al_and2 _2037_ (
    .a(g109),
    .b(\DFF_24.Q ),
    .y(\DFF_169.D )
  );
  al_and2 _2038_ (
    .a(g109),
    .b(\DFF_416.Q ),
    .y(\DFF_416.D )
  );
  al_or3fft _2039_ (
    .a(\DFF_12.Q ),
    .b(\DFF_264.Q ),
    .c(_0548_),
    .y(_0553_)
  );
  al_mux2l _2040_ (
    .a(_0549_),
    .b(_0548_),
    .s(\DFF_12.Q ),
    .y(_0554_)
  );
  al_and3fft _2041_ (
    .a(_0550_),
    .b(_0554_),
    .c(_0553_),
    .y(\DFF_12.D )
  );
  al_and2 _2042_ (
    .a(\DFF_163.Q ),
    .b(g109),
    .y(\DFF_132.D )
  );
  al_nor2 _2043_ (
    .a(g30),
    .b(_0009_),
    .y(_0555_)
  );
  al_nand3 _2044_ (
    .a(_0555_),
    .b(_0314_),
    .c(_0313_),
    .y(g10801)
  );
  al_oa21 _2045_ (
    .a(_0331_),
    .b(_0539_),
    .c(_0334_),
    .y(_0556_)
  );
  al_and3 _2046_ (
    .a(_0326_),
    .b(_0327_),
    .c(_0556_),
    .y(_0557_)
  );
  al_nand2ft _2047_ (
    .a(_0347_),
    .b(_0346_),
    .y(_0558_)
  );
  al_and3 _2048_ (
    .a(_0323_),
    .b(_0324_),
    .c(_0558_),
    .y(_0559_)
  );
  al_inv _2049_ (
    .a(\DFF_405.Q ),
    .y(_0560_)
  );
  al_ao21 _2050_ (
    .a(g109),
    .b(\DFF_22.D ),
    .c(_0560_),
    .y(_0561_)
  );
  al_and3 _2051_ (
    .a(g109),
    .b(_0560_),
    .c(\DFF_22.D ),
    .y(_0562_)
  );
  al_and3ftt _2052_ (
    .a(_0562_),
    .b(_0561_),
    .c(_0348_),
    .y(_0563_)
  );
  al_and3ftt _2053_ (
    .a(_0342_),
    .b(_0329_),
    .c(_0343_),
    .y(_0564_)
  );
  al_and2 _2054_ (
    .a(g109),
    .b(\DFF_116.D ),
    .y(_0565_)
  );
  al_ao21ttf _2055_ (
    .a(_0328_),
    .b(_0565_),
    .c(_0335_),
    .y(_0566_)
  );
  al_nand3ftt _2056_ (
    .a(_0566_),
    .b(_0564_),
    .c(_0563_),
    .y(_0567_)
  );
  al_nand3ftt _2057_ (
    .a(_0567_),
    .b(_0557_),
    .c(_0559_),
    .y(_0568_)
  );
  al_ao21 _2058_ (
    .a(_0354_),
    .b(_0568_),
    .c(_0357_),
    .y(_0569_)
  );
  al_inv _2059_ (
    .a(\DFF_19.Q ),
    .y(_0570_)
  );
  al_aoi21 _2060_ (
    .a(_0570_),
    .b(_0569_),
    .c(_0534_),
    .y(_0571_)
  );
  al_aoi21ftf _2061_ (
    .a(_0569_),
    .b(\DFF_19.Q ),
    .c(_0571_),
    .y(\DFF_19.D )
  );
  al_and2 _2062_ (
    .a(g109),
    .b(\DFF_90.Q ),
    .y(\DFF_494.D )
  );
  al_or3fft _2063_ (
    .a(\DFF_361.Q ),
    .b(\DFF_0.Q ),
    .c(_0443_),
    .y(_0572_)
  );
  al_aoi21ftf _2064_ (
    .a(\DFF_418.Q ),
    .b(_0572_),
    .c(_0530_),
    .y(_0573_)
  );
  al_aoi21ttf _2065_ (
    .a(_0411_),
    .b(_0444_),
    .c(_0573_),
    .y(\DFF_418.D )
  );
  al_and2 _2066_ (
    .a(\DFF_142.Q ),
    .b(g109),
    .y(\DFF_185.D )
  );
  al_and2ft _2067_ (
    .a(\DFF_237.Q ),
    .b(\DFF_34.Q ),
    .y(_0574_)
  );
  al_nand2ft _2068_ (
    .a(\DFF_34.Q ),
    .b(\DFF_237.Q ),
    .y(_0575_)
  );
  al_nor2 _2069_ (
    .a(\DFF_201.Q ),
    .b(\DFF_519.Q ),
    .y(_0576_)
  );
  al_nand2 _2070_ (
    .a(\DFF_201.Q ),
    .b(\DFF_519.Q ),
    .y(_0577_)
  );
  al_nand2ft _2071_ (
    .a(_0576_),
    .b(_0577_),
    .y(_0578_)
  );
  al_nand3ftt _2072_ (
    .a(_0574_),
    .b(_0575_),
    .c(_0578_),
    .y(_0579_)
  );
  al_ao21ftt _2073_ (
    .a(_0574_),
    .b(_0575_),
    .c(_0578_),
    .y(_0580_)
  );
  al_and3 _2074_ (
    .a(g109),
    .b(_0579_),
    .c(_0580_),
    .y(\DFF_237.D )
  );
  al_or3fft _2075_ (
    .a(\DFF_198.Q ),
    .b(\DFF_470.Q ),
    .c(_0528_),
    .y(_0581_)
  );
  al_aoi21ttf _2076_ (
    .a(\DFF_328.D ),
    .b(\DFF_335.D ),
    .c(_0531_),
    .y(_0582_)
  );
  al_aoi21ftf _2077_ (
    .a(\DFF_506.Q ),
    .b(_0581_),
    .c(_0582_),
    .y(\DFF_506.D )
  );
  al_inv _2078_ (
    .a(_0356_),
    .y(_0583_)
  );
  al_aoi21 _2079_ (
    .a(_0354_),
    .b(_0568_),
    .c(_0583_),
    .y(_0584_)
  );
  al_mux2l _2080_ (
    .a(\DFF_483.Q ),
    .b(_0584_),
    .s(_0534_),
    .y(\DFF_483.D )
  );
  al_inv _2081_ (
    .a(\DFF_190.Q ),
    .y(_0585_)
  );
  al_nor2 _2082_ (
    .a(\DFF_147.Q ),
    .b(\DFF_296.Q ),
    .y(_0586_)
  );
  al_nand3fft _2083_ (
    .a(\DFF_474.Q ),
    .b(\DFF_490.Q ),
    .c(_0586_),
    .y(_0587_)
  );
  al_and3fft _2084_ (
    .a(\DFF_444.Q ),
    .b(_0587_),
    .c(_0585_),
    .y(_0588_)
  );
  al_nand3ftt _2085_ (
    .a(\DFF_380.Q ),
    .b(\DFF_473.Q ),
    .c(g18),
    .y(_0589_)
  );
  al_or2 _2086_ (
    .a(\DFF_382.Q ),
    .b(\DFF_337.Q ),
    .y(_0590_)
  );
  al_nor3ftt _2087_ (
    .a(\DFF_307.Q ),
    .b(_0589_),
    .c(_0590_),
    .y(_0591_)
  );
  al_and2 _2088_ (
    .a(\DFF_314.Q ),
    .b(\DFF_220.Q ),
    .y(_0592_)
  );
  al_nand2 _2089_ (
    .a(\DFF_102.Q ),
    .b(\DFF_364.Q ),
    .y(_0593_)
  );
  al_and3fft _2090_ (
    .a(\DFF_508.Q ),
    .b(_0593_),
    .c(_0592_),
    .y(_0594_)
  );
  al_and3 _2091_ (
    .a(_0591_),
    .b(_0594_),
    .c(_0588_),
    .y(_0595_)
  );
  al_mux2l _2092_ (
    .a(\DFF_4.Q ),
    .b(_0595_),
    .s(_0151_),
    .y(\DFF_4.D )
  );
  al_and3ftt _2093_ (
    .a(\DFF_372.Q ),
    .b(g1696),
    .c(\DFF_103.Q ),
    .y(_0596_)
  );
  al_nand2 _2094_ (
    .a(\DFF_332.Q ),
    .b(\DFF_523.Q ),
    .y(_0597_)
  );
  al_or3fft _2095_ (
    .a(\DFF_268.Q ),
    .b(_0596_),
    .c(_0597_),
    .y(_0598_)
  );
  al_inv _2096_ (
    .a(\DFF_59.Q ),
    .y(_0599_)
  );
  al_aoi21 _2097_ (
    .a(_0599_),
    .b(_0598_),
    .c(\DFF_174.Q ),
    .y(_0600_)
  );
  al_aoi21ftf _2098_ (
    .a(_0598_),
    .b(\DFF_59.Q ),
    .c(_0600_),
    .y(\DFF_59.D )
  );
  al_nand2 _2099_ (
    .a(\DFF_125.Q ),
    .b(g18),
    .y(_0601_)
  );
  al_aoi21ftf _2100_ (
    .a(g18),
    .b(\DFF_516.Q ),
    .c(_0601_),
    .y(_0602_)
  );
  al_oa21ftf _2101_ (
    .a(\DFF_277.Q ),
    .b(_0602_),
    .c(_0151_),
    .y(_0603_)
  );
  al_aoi21ftf _2102_ (
    .a(\DFF_277.Q ),
    .b(_0602_),
    .c(_0603_),
    .y(\DFF_95.D )
  );
  al_and3fft _2103_ (
    .a(\DFF_54.Q ),
    .b(\DFF_112.Q ),
    .c(g109),
    .y(\DFF_112.D )
  );
  al_ao21ftf _2104_ (
    .a(g18),
    .b(\DFF_288.Q ),
    .c(_0521_),
    .y(\DFF_443.D )
  );
  al_aoi21 _2105_ (
    .a(\DFF_508.Q ),
    .b(\DFF_443.D ),
    .c(_0151_),
    .y(_0604_)
  );
  al_oa21 _2106_ (
    .a(\DFF_508.Q ),
    .b(\DFF_443.D ),
    .c(_0604_),
    .y(\DFF_314.D )
  );
  al_and3ftt _2107_ (
    .a(\DFF_111.Q ),
    .b(\DFF_223.Q ),
    .c(_0457_),
    .y(_0605_)
  );
  al_mux2l _2108_ (
    .a(_0459_),
    .b(_0483_),
    .s(_0605_),
    .y(_0606_)
  );
  al_inv _2109_ (
    .a(\DFF_455.Q ),
    .y(_0607_)
  );
  al_mux2l _2110_ (
    .a(_0607_),
    .b(_0606_),
    .s(_0489_),
    .y(_0608_)
  );
  al_aoi21ftf _2111_ (
    .a(\DFF_455.Q ),
    .b(_0606_),
    .c(_0608_),
    .y(\DFF_455.D )
  );
  al_and2 _2112_ (
    .a(\DFF_237.Q ),
    .b(g109),
    .y(\DFF_165.D )
  );
  al_and2 _2113_ (
    .a(\DFF_189.Q ),
    .b(g109),
    .y(\DFF_105.D )
  );
  al_mux2h _2114_ (
    .a(\DFF_253.Q ),
    .b(_0447_),
    .s(_0452_),
    .y(_0609_)
  );
  al_aoi21ttf _2115_ (
    .a(\DFF_253.Q ),
    .b(_0447_),
    .c(_0609_),
    .y(\DFF_253.D )
  );
  al_nor2 _2116_ (
    .a(\DFF_303.Q ),
    .b(\DFF_125.Q ),
    .y(_0610_)
  );
  al_or3 _2117_ (
    .a(\DFF_67.Q ),
    .b(\DFF_396.Q ),
    .c(\DFF_5.Q ),
    .y(_0611_)
  );
  al_and3fft _2118_ (
    .a(\DFF_185.Q ),
    .b(_0611_),
    .c(_0610_),
    .y(_0612_)
  );
  al_nor2 _2119_ (
    .a(\DFF_189.Q ),
    .b(\DFF_327.Q ),
    .y(_0613_)
  );
  al_nand3fft _2120_ (
    .a(\DFF_88.Q ),
    .b(\DFF_487.Q ),
    .c(_0613_),
    .y(_0614_)
  );
  al_or3 _2121_ (
    .a(\DFF_331.Q ),
    .b(\DFF_163.Q ),
    .c(_0614_),
    .y(_0615_)
  );
  al_nor2 _2122_ (
    .a(\DFF_142.Q ),
    .b(\DFF_132.Q ),
    .y(_0616_)
  );
  al_and3fft _2123_ (
    .a(\DFF_105.Q ),
    .b(\DFF_33.Q ),
    .c(_0616_),
    .y(_0617_)
  );
  al_or3fft _2124_ (
    .a(_0612_),
    .b(_0617_),
    .c(_0615_),
    .y(_0618_)
  );
  al_or3 _2125_ (
    .a(\DFF_484.Q ),
    .b(\DFF_76.Q ),
    .c(\DFF_284.Q ),
    .y(_0619_)
  );
  al_nor2 _2126_ (
    .a(\DFF_424.Q ),
    .b(\DFF_66.Q ),
    .y(_0620_)
  );
  al_or2 _2127_ (
    .a(\DFF_182.Q ),
    .b(\DFF_153.Q ),
    .y(_0621_)
  );
  al_and3fft _2128_ (
    .a(_0621_),
    .b(_0619_),
    .c(_0620_),
    .y(_0622_)
  );
  al_and3fft _2129_ (
    .a(\DFF_400.Q ),
    .b(_0618_),
    .c(_0622_),
    .y(_0623_)
  );
  al_nand2 _2130_ (
    .a(\DFF_424.Q ),
    .b(\DFF_66.Q ),
    .y(_0624_)
  );
  al_nor2 _2131_ (
    .a(\DFF_400.Q ),
    .b(\DFF_396.Q ),
    .y(_0625_)
  );
  al_nand2 _2132_ (
    .a(\DFF_400.Q ),
    .b(\DFF_396.Q ),
    .y(_0626_)
  );
  al_nand2ft _2133_ (
    .a(_0625_),
    .b(_0626_),
    .y(_0627_)
  );
  al_and3ftt _2134_ (
    .a(_0620_),
    .b(_0624_),
    .c(_0627_),
    .y(_0628_)
  );
  al_ao21ftt _2135_ (
    .a(_0620_),
    .b(_0624_),
    .c(_0627_),
    .y(_0629_)
  );
  al_nand2ft _2136_ (
    .a(_0628_),
    .b(_0629_),
    .y(_0630_)
  );
  al_mux2h _2137_ (
    .a(_0630_),
    .b(_0623_),
    .s(g109),
    .y(\DFF_400.D )
  );
  al_nand2 _2138_ (
    .a(\DFF_473.Q ),
    .b(g18),
    .y(_0631_)
  );
  al_aoi21ftf _2139_ (
    .a(\DFF_531.Q ),
    .b(_0631_),
    .c(g109),
    .y(\DFF_531.D )
  );
  al_and3ftt _2140_ (
    .a(\DFF_126.Q ),
    .b(\DFF_278.Q ),
    .c(g109),
    .y(\DFF_278.D )
  );
  al_and2 _2141_ (
    .a(\DFF_153.Q ),
    .b(g109),
    .y(\DFF_76.D )
  );
  al_and2 _2142_ (
    .a(\DFF_13.Q ),
    .b(_0486_),
    .y(\DFF_13.D )
  );
  al_oa21ftt _2143_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_472.Q ),
    .y(\DFF_472.D )
  );
  al_or2 _2144_ (
    .a(g82),
    .b(\DFF_213.Q ),
    .y(g8316)
  );
  al_and2 _2145_ (
    .a(\DFF_66.Q ),
    .b(g109),
    .y(\DFF_284.D )
  );
  al_oa21ftt _2146_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_63.Q ),
    .y(\DFF_63.D )
  );
  al_inv _2147_ (
    .a(\DFF_387.Q ),
    .y(_0632_)
  );
  al_nand2 _2148_ (
    .a(_0632_),
    .b(_0507_),
    .y(_0633_)
  );
  al_and3 _2149_ (
    .a(_0455_),
    .b(_0510_),
    .c(_0633_),
    .y(\DFF_387.D )
  );
  al_mux2l _2150_ (
    .a(_0529_),
    .b(_0528_),
    .s(\DFF_198.Q ),
    .y(_0634_)
  );
  al_nor3fft _2151_ (
    .a(_0531_),
    .b(_0581_),
    .c(_0634_),
    .y(\DFF_198.D )
  );
  al_nor2ft _2152_ (
    .a(\DFF_336.Q ),
    .b(\DFF_262.D ),
    .y(\DFF_136.D )
  );
  al_and2 _2153_ (
    .a(g109),
    .b(\DFF_145.Q ),
    .y(\DFF_145.D )
  );
  al_and2 _2154_ (
    .a(\DFF_400.Q ),
    .b(g109),
    .y(\DFF_484.D )
  );
  al_nor3fft _2155_ (
    .a(_0622_),
    .b(\DFF_484.D ),
    .c(_0618_),
    .y(\DFF_452.D )
  );
  al_and2 _2156_ (
    .a(\DFF_289.Q ),
    .b(\DFF_452.D ),
    .y(\DFF_473.D )
  );
  al_nor2 _2157_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .y(_0635_)
  );
  al_and3ftt _2158_ (
    .a(\DFF_174.Q ),
    .b(\DFF_0.Q ),
    .c(_0635_),
    .y(_0636_)
  );
  al_and3 _2159_ (
    .a(\DFF_119.Q ),
    .b(_0410_),
    .c(_0636_),
    .y(_0637_)
  );
  al_mux2h _2160_ (
    .a(\DFF_28.Q ),
    .b(_0637_),
    .s(_0530_),
    .y(\DFF_28.D )
  );
  al_and3 _2161_ (
    .a(g109),
    .b(g742),
    .c(g741),
    .y(g5658)
  );
  al_aoi21 _2162_ (
    .a(_0354_),
    .b(_0568_),
    .c(_0547_),
    .y(_0638_)
  );
  al_mux2l _2163_ (
    .a(\DFF_152.Q ),
    .b(_0638_),
    .s(_0550_),
    .y(\DFF_152.D )
  );
  al_inv _2164_ (
    .a(\DFF_174.Q ),
    .y(_0639_)
  );
  al_and3fft _2165_ (
    .a(_0599_),
    .b(_0598_),
    .c(\DFF_75.Q ),
    .y(_0640_)
  );
  al_aoi21 _2166_ (
    .a(\DFF_324.Q ),
    .b(_0640_),
    .c(\DFF_104.Q ),
    .y(_0641_)
  );
  al_and3 _2167_ (
    .a(\DFF_324.Q ),
    .b(\DFF_104.Q ),
    .c(_0640_),
    .y(_0642_)
  );
  al_nor3ftt _2168_ (
    .a(_0639_),
    .b(_0642_),
    .c(_0641_),
    .y(\DFF_104.D )
  );
  al_oa21ftt _2169_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_421.Q ),
    .y(\DFF_421.D )
  );
  al_and2 _2170_ (
    .a(\DFF_484.Q ),
    .b(g109),
    .y(\DFF_424.D )
  );
  al_or2ft _2171_ (
    .a(_0555_),
    .b(\DFF_228.D ),
    .y(g10461)
  );
  al_aoi21 _2172_ (
    .a(\DFF_247.Q ),
    .b(_0448_),
    .c(\DFF_301.Q ),
    .y(_0643_)
  );
  al_nor3ftt _2173_ (
    .a(_0452_),
    .b(_0449_),
    .c(_0643_),
    .y(\DFF_301.D )
  );
  al_aoi21ftf _2174_ (
    .a(\DFF_369.Q ),
    .b(_0483_),
    .c(g18),
    .y(_0644_)
  );
  al_oa21 _2175_ (
    .a(\DFF_302.Q ),
    .b(_0483_),
    .c(_0644_),
    .y(\DFF_302.D )
  );
  al_aoi21ftf _2176_ (
    .a(\DFF_179.Q ),
    .b(_0631_),
    .c(g109),
    .y(\DFF_179.D )
  );
  al_aoi21ftf _2177_ (
    .a(g18),
    .b(\DFF_249.Q ),
    .c(_0521_),
    .y(_0645_)
  );
  al_oa21ftf _2178_ (
    .a(\DFF_172.Q ),
    .b(_0645_),
    .c(_0151_),
    .y(_0646_)
  );
  al_aoi21ftf _2179_ (
    .a(\DFF_172.Q ),
    .b(_0645_),
    .c(_0646_),
    .y(\DFF_273.D )
  );
  al_and2 _2180_ (
    .a(\DFF_284.Q ),
    .b(g109),
    .y(\DFF_153.D )
  );
  al_aoi21ftf _2181_ (
    .a(\DFF_111.Q ),
    .b(_0457_),
    .c(_0512_),
    .y(_0647_)
  );
  al_oai21ftt _2182_ (
    .a(\DFF_352.Q ),
    .b(\DFF_141.Q ),
    .c(\DFF_18.Q ),
    .y(_0648_)
  );
  al_aoi21ftf _2183_ (
    .a(_0457_),
    .b(_0648_),
    .c(_0647_),
    .y(\DFF_18.D )
  );
  al_or2ft _2184_ (
    .a(_0555_),
    .b(\DFF_22.D ),
    .y(g10377)
  );
  al_and3 _2185_ (
    .a(g109),
    .b(g744),
    .c(g743),
    .y(g5659)
  );
  al_and2 _2186_ (
    .a(g109),
    .b(\DFF_494.Q ),
    .y(\DFF_315.D )
  );
  al_and2 _2187_ (
    .a(\DFF_340.Q ),
    .b(\DFF_83.Q ),
    .y(_0649_)
  );
  al_and3 _2188_ (
    .a(\DFF_243.Q ),
    .b(\DFF_13.Q ),
    .c(_0649_),
    .y(\DFF_291.D )
  );
  al_mux2l _2189_ (
    .a(_0599_),
    .b(_0598_),
    .s(\DFF_75.Q ),
    .y(_0650_)
  );
  al_nor3ftt _2190_ (
    .a(_0639_),
    .b(_0640_),
    .c(_0650_),
    .y(\DFF_75.D )
  );
  al_and3ftt _2191_ (
    .a(\DFF_126.Q ),
    .b(\DFF_31.Q ),
    .c(g109),
    .y(\DFF_31.D )
  );
  al_nand2 _2192_ (
    .a(\DFF_132.Q ),
    .b(g18),
    .y(_0651_)
  );
  al_ao21ftf _2193_ (
    .a(g18),
    .b(\DFF_208.Q ),
    .c(_0651_),
    .y(\DFF_193.D )
  );
  al_aoi21 _2194_ (
    .a(\DFF_314.Q ),
    .b(\DFF_193.D ),
    .c(_0151_),
    .y(_0652_)
  );
  al_oa21 _2195_ (
    .a(\DFF_314.Q ),
    .b(\DFF_193.D ),
    .c(_0652_),
    .y(\DFF_102.D )
  );
  al_and2ft _2196_ (
    .a(\DFF_118.Q ),
    .b(\DFF_90.Q ),
    .y(_0653_)
  );
  al_and3 _2197_ (
    .a(\DFF_36.Q ),
    .b(\DFF_24.Q ),
    .c(_0653_),
    .y(_0654_)
  );
  al_nand3fft _2198_ (
    .a(_0487_),
    .b(_0497_),
    .c(_0654_),
    .y(_0655_)
  );
  al_nand3ftt _2199_ (
    .a(\DFF_531.Q ),
    .b(\DFF_473.Q ),
    .c(g18),
    .y(_0656_)
  );
  al_nor3fft _2200_ (
    .a(\DFF_494.Q ),
    .b(\DFF_503.Q ),
    .c(_0656_),
    .y(_0657_)
  );
  al_inv _2201_ (
    .a(\DFF_47.Q ),
    .y(_0658_)
  );
  al_and2ft _2202_ (
    .a(\DFF_169.Q ),
    .b(\DFF_143.Q ),
    .y(_0659_)
  );
  al_and3ftt _2203_ (
    .a(\DFF_415.Q ),
    .b(\DFF_315.Q ),
    .c(_0659_),
    .y(_0660_)
  );
  al_nand3fft _2204_ (
    .a(\DFF_109.Q ),
    .b(_0658_),
    .c(_0660_),
    .y(_0661_)
  );
  al_nor3ftt _2205_ (
    .a(_0657_),
    .b(_0655_),
    .c(_0661_),
    .y(_0662_)
  );
  al_mux2l _2206_ (
    .a(\DFF_528.Q ),
    .b(_0662_),
    .s(_0151_),
    .y(\DFF_528.D )
  );
  al_and2 _2207_ (
    .a(\DFF_5.Q ),
    .b(g109),
    .y(\DFF_189.D )
  );
  al_or2 _2208_ (
    .a(g82),
    .b(\DFF_287.Q ),
    .y(g8323)
  );
  al_oa21ftt _2209_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_224.Q ),
    .y(\DFF_224.D )
  );
  al_ao21 _2210_ (
    .a(_0320_),
    .b(\DFF_37.D ),
    .c(\DFF_293.Q ),
    .y(_0663_)
  );
  al_nand2 _2211_ (
    .a(\DFF_53.D ),
    .b(\DFF_37.D ),
    .y(_0664_)
  );
  al_and3ftt _2212_ (
    .a(_0537_),
    .b(_0664_),
    .c(_0663_),
    .y(\DFF_293.D )
  );
  al_and2 _2213_ (
    .a(g109),
    .b(\DFF_307.Q ),
    .y(\DFF_364.D )
  );
  al_or3 _2214_ (
    .a(g30),
    .b(_0009_),
    .c(\DFF_384.D ),
    .y(g10457)
  );
  al_and2 _2215_ (
    .a(g109),
    .b(\DFF_353.Q ),
    .y(\DFF_353.D )
  );
  al_or2 _2216_ (
    .a(g82),
    .b(\DFF_91.Q ),
    .y(g8318)
  );
  al_and3fft _2217_ (
    .a(\DFF_518.Q ),
    .b(\DFF_64.Q ),
    .c(\DFF_191.Q ),
    .y(_0665_)
  );
  al_or2ft _2218_ (
    .a(\DFF_403.Q ),
    .b(_0665_),
    .y(_0666_)
  );
  al_and2ft _2219_ (
    .a(\DFF_403.Q ),
    .b(_0665_),
    .y(_0667_)
  );
  al_or3 _2220_ (
    .a(\DFF_362.Q ),
    .b(\DFF_310.Q ),
    .c(\DFF_135.Q ),
    .y(_0668_)
  );
  al_nand3fft _2221_ (
    .a(\DFF_403.Q ),
    .b(\DFF_196.Q ),
    .c(_0665_),
    .y(_0669_)
  );
  al_oa21 _2222_ (
    .a(\DFF_358.Q ),
    .b(_0668_),
    .c(_0669_),
    .y(_0670_)
  );
  al_aoi21ftf _2223_ (
    .a(_0667_),
    .b(_0666_),
    .c(_0670_),
    .y(\DFF_403.D )
  );
  al_and3ftt _2224_ (
    .a(\DFF_126.Q ),
    .b(\DFF_158.Q ),
    .c(g109),
    .y(\DFF_158.D )
  );
  al_inv _2225_ (
    .a(\DFF_155.Q ),
    .y(_0671_)
  );
  al_nand3fft _2226_ (
    .a(\DFF_455.Q ),
    .b(_0671_),
    .c(_0605_),
    .y(_0672_)
  );
  al_and2ft _2227_ (
    .a(\DFF_111.Q ),
    .b(_0457_),
    .y(_0673_)
  );
  al_or3ftt _2228_ (
    .a(\DFF_297.Q ),
    .b(\DFF_223.Q ),
    .c(_0515_),
    .y(_0674_)
  );
  al_ao21ftt _2229_ (
    .a(_0674_),
    .b(_0673_),
    .c(\DFF_223.Q ),
    .y(_0675_)
  );
  al_and3 _2230_ (
    .a(g18),
    .b(_0672_),
    .c(_0675_),
    .y(\DFF_223.D )
  );
  al_and2 _2231_ (
    .a(\DFF_337.Q ),
    .b(g109),
    .y(\DFF_307.D )
  );
  al_mux2l _2232_ (
    .a(_0632_),
    .b(_0507_),
    .s(\DFF_99.Q ),
    .y(_0676_)
  );
  al_nor3fft _2233_ (
    .a(_0455_),
    .b(_0508_),
    .c(_0676_),
    .y(\DFF_99.D )
  );
  al_or3fft _2234_ (
    .a(_0120_),
    .b(_0555_),
    .c(_0284_),
    .y(g10455)
  );
  al_and2 _2235_ (
    .a(\DFF_105.Q ),
    .b(g109),
    .y(\DFF_396.D )
  );
  al_nor2ft _2236_ (
    .a(\DFF_117.Q ),
    .b(\DFF_262.D ),
    .y(\DFF_157.D )
  );
  al_and3ftt _2237_ (
    .a(\DFF_261.Q ),
    .b(\DFF_358.Q ),
    .c(\DFF_135.Q ),
    .y(_0677_)
  );
  al_inv _2238_ (
    .a(\DFF_359.Q ),
    .y(_0678_)
  );
  al_inv _2239_ (
    .a(\DFF_6.Q ),
    .y(_0679_)
  );
  al_inv _2240_ (
    .a(\DFF_286.Q ),
    .y(_0680_)
  );
  al_and3fft _2241_ (
    .a(\DFF_358.Q ),
    .b(\DFF_310.Q ),
    .c(\DFF_362.Q ),
    .y(_0681_)
  );
  al_and2ft _2242_ (
    .a(\DFF_362.Q ),
    .b(\DFF_310.Q ),
    .y(_0682_)
  );
  al_aoi21ftt _2243_ (
    .a(\DFF_358.Q ),
    .b(_0682_),
    .c(_0681_),
    .y(_0683_)
  );
  al_ao21ftf _2244_ (
    .a(\DFF_310.Q ),
    .b(\DFF_358.Q ),
    .c(_0683_),
    .y(_0684_)
  );
  al_and3 _2245_ (
    .a(\DFF_381.Q ),
    .b(\DFF_395.Q ),
    .c(_0684_),
    .y(_0685_)
  );
  al_and3 _2246_ (
    .a(\DFF_316.Q ),
    .b(\DFF_450.Q ),
    .c(_0685_),
    .y(_0686_)
  );
  al_and3 _2247_ (
    .a(\DFF_57.Q ),
    .b(\DFF_11.Q ),
    .c(_0686_),
    .y(_0687_)
  );
  al_nand3fft _2248_ (
    .a(_0679_),
    .b(_0680_),
    .c(_0687_),
    .y(_0688_)
  );
  al_inv _2249_ (
    .a(\DFF_72.Q ),
    .y(_0689_)
  );
  al_or3 _2250_ (
    .a(_0689_),
    .b(_0396_),
    .c(_0669_),
    .y(_0690_)
  );
  al_aoi21ftf _2251_ (
    .a(_0669_),
    .b(_0677_),
    .c(_0690_),
    .y(_0691_)
  );
  al_inv _2252_ (
    .a(\DFF_57.Q ),
    .y(_0692_)
  );
  al_inv _2253_ (
    .a(\DFF_11.Q ),
    .y(_0693_)
  );
  al_inv _2254_ (
    .a(\DFF_450.Q ),
    .y(_0694_)
  );
  al_inv _2255_ (
    .a(\DFF_381.Q ),
    .y(_0695_)
  );
  al_and3fft _2256_ (
    .a(\DFF_395.Q ),
    .b(_0684_),
    .c(_0695_),
    .y(_0696_)
  );
  al_and3ftt _2257_ (
    .a(\DFF_316.Q ),
    .b(_0694_),
    .c(_0696_),
    .y(_0697_)
  );
  al_and3 _2258_ (
    .a(_0692_),
    .b(_0693_),
    .c(_0697_),
    .y(_0698_)
  );
  al_and3 _2259_ (
    .a(_0679_),
    .b(_0680_),
    .c(_0698_),
    .y(_0699_)
  );
  al_mux2l _2260_ (
    .a(\DFF_359.Q ),
    .b(_0699_),
    .s(_0691_),
    .y(_0700_)
  );
  al_aoi21ftf _2261_ (
    .a(_0678_),
    .b(_0688_),
    .c(_0700_),
    .y(_0701_)
  );
  al_or3ftt _2262_ (
    .a(_0677_),
    .b(_0669_),
    .c(_0701_),
    .y(_0702_)
  );
  al_or3ftt _2263_ (
    .a(_0677_),
    .b(\DFF_43.Q ),
    .c(_0669_),
    .y(_0703_)
  );
  al_and3ftt _2264_ (
    .a(\DFF_196.Q ),
    .b(\DFF_261.Q ),
    .c(_0667_),
    .y(_0704_)
  );
  al_and3ftt _2265_ (
    .a(_0704_),
    .b(_0703_),
    .c(_0702_),
    .y(_0705_)
  );
  al_inv _2266_ (
    .a(\DFF_135.Q ),
    .y(_0706_)
  );
  al_mux2l _2267_ (
    .a(_0706_),
    .b(_0705_),
    .s(_0489_),
    .y(_0707_)
  );
  al_aoi21ftf _2268_ (
    .a(\DFF_135.Q ),
    .b(_0705_),
    .c(_0707_),
    .y(\DFF_135.D )
  );
  al_and2 _2269_ (
    .a(g109),
    .b(\DFF_7.Q ),
    .y(\DFF_7.D )
  );
  al_nand2 _2270_ (
    .a(\DFF_303.Q ),
    .b(g18),
    .y(_0708_)
  );
  al_ao21ftf _2271_ (
    .a(g18),
    .b(\DFF_524.Q ),
    .c(_0708_),
    .y(\DFF_244.D )
  );
  al_aoi21 _2272_ (
    .a(\DFF_444.Q ),
    .b(\DFF_244.D ),
    .c(_0151_),
    .y(_0709_)
  );
  al_oa21 _2273_ (
    .a(\DFF_444.Q ),
    .b(\DFF_244.D ),
    .c(_0709_),
    .y(\DFF_508.D )
  );
  al_aoi21 _2274_ (
    .a(\DFF_253.Q ),
    .b(_0447_),
    .c(\DFF_30.Q ),
    .y(_0710_)
  );
  al_nor3ftt _2275_ (
    .a(_0452_),
    .b(_0448_),
    .c(_0710_),
    .y(\DFF_30.D )
  );
  al_aoi21 _2276_ (
    .a(_0320_),
    .b(\DFF_37.D ),
    .c(_0537_),
    .y(_0711_)
  );
  al_aoi21ftf _2277_ (
    .a(\DFF_52.Q ),
    .b(_0533_),
    .c(_0711_),
    .y(\DFF_52.D )
  );
  al_and2 _2278_ (
    .a(g109),
    .b(\DFF_457.Q ),
    .y(\DFF_457.D )
  );
  al_nand2 _2279_ (
    .a(\DFF_284.Q ),
    .b(g18),
    .y(_0712_)
  );
  al_aoi21ftf _2280_ (
    .a(g18),
    .b(\DFF_435.Q ),
    .c(_0712_),
    .y(_0713_)
  );
  al_oa21ftf _2281_ (
    .a(\DFF_165.Q ),
    .b(_0713_),
    .c(_0151_),
    .y(_0714_)
  );
  al_aoi21ftf _2282_ (
    .a(\DFF_165.Q ),
    .b(_0713_),
    .c(_0714_),
    .y(\DFF_306.D )
  );
  al_ao21ftf _2283_ (
    .a(g18),
    .b(\DFF_260.Q ),
    .c(_0601_),
    .y(\DFF_446.D )
  );
  al_aoi21 _2284_ (
    .a(\DFF_102.Q ),
    .b(\DFF_446.D ),
    .c(_0151_),
    .y(_0715_)
  );
  al_oa21 _2285_ (
    .a(\DFF_102.Q ),
    .b(\DFF_446.D ),
    .c(_0715_),
    .y(\DFF_490.D )
  );
  al_mux2l _2286_ (
    .a(\DFF_268.Q ),
    .b(_0596_),
    .s(\DFF_174.Q ),
    .y(_0716_)
  );
  al_aoi21ttf _2287_ (
    .a(\DFF_268.Q ),
    .b(_0596_),
    .c(_0716_),
    .y(\DFF_268.D )
  );
  al_and2 _2288_ (
    .a(g109),
    .b(\DFF_109.Q ),
    .y(\DFF_24.D )
  );
  al_and2 _2289_ (
    .a(\DFF_132.Q ),
    .b(g109),
    .y(\DFF_67.D )
  );
  al_mux2h _2290_ (
    .a(\DFF_247.Q ),
    .b(_0448_),
    .s(_0452_),
    .y(_0717_)
  );
  al_aoi21ttf _2291_ (
    .a(\DFF_247.Q ),
    .b(_0448_),
    .c(_0717_),
    .y(\DFF_247.D )
  );
  al_oa21ftt _2292_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_513.Q ),
    .y(\DFF_513.D )
  );
  al_and2 _2293_ (
    .a(\DFF_125.Q ),
    .b(g109),
    .y(\DFF_327.D )
  );
  al_and2 _2294_ (
    .a(\DFF_424.Q ),
    .b(g109),
    .y(\DFF_66.D )
  );
  al_ao21ftf _2295_ (
    .a(g18),
    .b(\DFF_159.Q ),
    .c(_0712_),
    .y(\DFF_270.D )
  );
  al_aoi21 _2296_ (
    .a(\DFF_220.Q ),
    .b(\DFF_270.D ),
    .c(_0151_),
    .y(_0718_)
  );
  al_oa21 _2297_ (
    .a(\DFF_220.Q ),
    .b(\DFF_270.D ),
    .c(_0718_),
    .y(\DFF_382.D )
  );
  al_mux2h _2298_ (
    .a(\DFF_38.Q ),
    .b(_0449_),
    .s(_0452_),
    .y(_0719_)
  );
  al_aoi21ttf _2299_ (
    .a(\DFF_38.Q ),
    .b(_0449_),
    .c(_0719_),
    .y(\DFF_38.D )
  );
  al_aoi21ftf _2300_ (
    .a(g18),
    .b(\DFF_482.Q ),
    .c(_0498_),
    .y(_0720_)
  );
  al_oa21ftf _2301_ (
    .a(\DFF_95.Q ),
    .b(_0720_),
    .c(_0151_),
    .y(_0721_)
  );
  al_aoi21ftf _2302_ (
    .a(\DFF_95.Q ),
    .b(_0720_),
    .c(_0721_),
    .y(\DFF_437.D )
  );
  al_or2 _2303_ (
    .a(g82),
    .b(\DFF_479.Q ),
    .y(g8331)
  );
  al_or2 _2304_ (
    .a(g82),
    .b(\DFF_224.Q ),
    .y(g8335)
  );
  al_oa21ftt _2305_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_323.Q ),
    .y(\DFF_323.D )
  );
  al_and2 _2306_ (
    .a(g109),
    .b(\DFF_399.Q ),
    .y(\DFF_399.D )
  );
  al_inv _2307_ (
    .a(\DFF_416.Q ),
    .y(_0722_)
  );
  al_ao21 _2308_ (
    .a(\DFF_158.Q ),
    .b(_0522_),
    .c(_0722_),
    .y(_0723_)
  );
  al_nand3ftt _2309_ (
    .a(\DFF_416.Q ),
    .b(\DFF_158.Q ),
    .c(_0522_),
    .y(_0724_)
  );
  al_ao21 _2310_ (
    .a(_0724_),
    .b(_0723_),
    .c(g18),
    .y(_0725_)
  );
  al_aoi21 _2311_ (
    .a(_0708_),
    .b(_0725_),
    .c(\DFF_143.Q ),
    .y(_0726_)
  );
  al_and3 _2312_ (
    .a(\DFF_143.Q ),
    .b(_0708_),
    .c(_0725_),
    .y(_0727_)
  );
  al_mux2l _2313_ (
    .a(_0727_),
    .b(_0726_),
    .s(_0151_),
    .y(\DFF_36.D )
  );
  al_aoi21ftf _2314_ (
    .a(\DFF_380.Q ),
    .b(_0631_),
    .c(g109),
    .y(\DFF_380.D )
  );
  al_nand2 _2315_ (
    .a(\DFF_76.Q ),
    .b(g18),
    .y(_0728_)
  );
  al_aoi21ftf _2316_ (
    .a(g18),
    .b(\DFF_404.Q ),
    .c(_0728_),
    .y(_0729_)
  );
  al_oa21ftf _2317_ (
    .a(\DFF_306.Q ),
    .b(_0729_),
    .c(_0151_),
    .y(_0730_)
  );
  al_aoi21ftf _2318_ (
    .a(\DFF_306.Q ),
    .b(_0729_),
    .c(_0730_),
    .y(\DFF_139.D )
  );
  al_inv _2319_ (
    .a(\DFF_346.Q ),
    .y(_0731_)
  );
  al_aoi21 _2320_ (
    .a(\DFF_346.Q ),
    .b(_0642_),
    .c(\DFF_174.Q ),
    .y(_0732_)
  );
  al_aoi21ftf _2321_ (
    .a(_0642_),
    .b(_0731_),
    .c(_0732_),
    .y(\DFF_346.D )
  );
  al_aoi21 _2322_ (
    .a(\DFF_294.Q ),
    .b(\DFF_37.D ),
    .c(_0537_),
    .y(_0733_)
  );
  al_oa21 _2323_ (
    .a(\DFF_294.Q ),
    .b(\DFF_37.D ),
    .c(_0733_),
    .y(\DFF_294.D )
  );
  al_nand2 _2324_ (
    .a(\DFF_5.Q ),
    .b(g18),
    .y(_0734_)
  );
  al_ao21ftf _2325_ (
    .a(g18),
    .b(\DFF_50.Q ),
    .c(_0734_),
    .y(\DFF_500.D )
  );
  al_aoi21 _2326_ (
    .a(\DFF_190.Q ),
    .b(\DFF_500.D ),
    .c(_0151_),
    .y(_0735_)
  );
  al_aoi21ftf _2327_ (
    .a(\DFF_500.D ),
    .b(_0585_),
    .c(_0735_),
    .y(\DFF_147.D )
  );
  al_oa21ftt _2328_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_363.Q ),
    .y(\DFF_363.D )
  );
  al_nand2 _2329_ (
    .a(\DFF_33.Q ),
    .b(g18),
    .y(_0736_)
  );
  al_ao21ftf _2330_ (
    .a(g18),
    .b(\DFF_166.Q ),
    .c(_0736_),
    .y(\DFF_222.D )
  );
  al_aoi21 _2331_ (
    .a(\DFF_474.Q ),
    .b(\DFF_222.D ),
    .c(_0151_),
    .y(_0737_)
  );
  al_oa21 _2332_ (
    .a(\DFF_474.Q ),
    .b(\DFF_222.D ),
    .c(_0737_),
    .y(\DFF_444.D )
  );
  al_or2 _2333_ (
    .a(g82),
    .b(\DFF_63.Q ),
    .y(g8313)
  );
  al_nand3ftt _2334_ (
    .a(\DFF_158.Q ),
    .b(\DFF_399.Q ),
    .c(_0499_),
    .y(_0738_)
  );
  al_ao21ftt _2335_ (
    .a(\DFF_158.Q ),
    .b(_0499_),
    .c(\DFF_399.Q ),
    .y(_0739_)
  );
  al_nand3 _2336_ (
    .a(_0489_),
    .b(_0738_),
    .c(_0739_),
    .y(_0740_)
  );
  al_aoi21 _2337_ (
    .a(_0734_),
    .b(_0740_),
    .c(\DFF_415.Q ),
    .y(_0741_)
  );
  al_and3 _2338_ (
    .a(\DFF_415.Q ),
    .b(_0734_),
    .c(_0740_),
    .y(_0742_)
  );
  al_mux2l _2339_ (
    .a(_0742_),
    .b(_0741_),
    .s(_0151_),
    .y(\DFF_128.D )
  );
  al_ao21 _2340_ (
    .a(_0445_),
    .b(_0442_),
    .c(\DFF_344.Q ),
    .y(_0743_)
  );
  al_and3 _2341_ (
    .a(_0531_),
    .b(_0528_),
    .c(_0743_),
    .y(\DFF_344.D )
  );
  al_mux2h _2342_ (
    .a(\DFF_119.Q ),
    .b(_0444_),
    .s(_0530_),
    .y(_0744_)
  );
  al_aoi21ftf _2343_ (
    .a(\DFF_28.Q ),
    .b(_0637_),
    .c(_0744_),
    .y(\DFF_119.D )
  );
  al_or2ft _2344_ (
    .a(_0555_),
    .b(\DFF_116.D ),
    .y(g10465)
  );
  al_and2 _2345_ (
    .a(g109),
    .b(\DFF_214.Q ),
    .y(\DFF_214.D )
  );
  al_or2 _2346_ (
    .a(\DFF_127.Q ),
    .b(_0453_),
    .y(_0745_)
  );
  al_nor3fft _2347_ (
    .a(_0455_),
    .b(_0745_),
    .c(_0454_),
    .y(\DFF_127.D )
  );
  al_nor2ft _2348_ (
    .a(\DFF_136.Q ),
    .b(\DFF_262.D ),
    .y(\DFF_117.D )
  );
  al_oa21ftt _2349_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_507.Q ),
    .y(\DFF_507.D )
  );
  al_and2 _2350_ (
    .a(g109),
    .b(\DFF_383.Q ),
    .y(\DFF_383.D )
  );
  al_ao21ftf _2351_ (
    .a(g18),
    .b(\DFF_460.Q ),
    .c(_0488_),
    .y(\DFF_397.D )
  );
  al_aoi21 _2352_ (
    .a(\DFF_147.Q ),
    .b(\DFF_397.D ),
    .c(_0151_),
    .y(_0746_)
  );
  al_oa21 _2353_ (
    .a(\DFF_147.Q ),
    .b(\DFF_397.D ),
    .c(_0746_),
    .y(\DFF_337.D )
  );
  al_ao21ftf _2354_ (
    .a(g18),
    .b(\DFF_74.Q ),
    .c(_0734_),
    .y(_0747_)
  );
  al_aoi21 _2355_ (
    .a(\DFF_437.Q ),
    .b(_0747_),
    .c(_0151_),
    .y(_0748_)
  );
  al_oa21 _2356_ (
    .a(\DFF_437.Q ),
    .b(_0747_),
    .c(_0748_),
    .y(\DFF_519.D )
  );
  al_and2 _2357_ (
    .a(\DFF_268.Q ),
    .b(_0596_),
    .y(_0749_)
  );
  al_mux2l _2358_ (
    .a(\DFF_523.Q ),
    .b(_0749_),
    .s(\DFF_174.Q ),
    .y(_0750_)
  );
  al_aoi21ttf _2359_ (
    .a(\DFF_523.Q ),
    .b(_0749_),
    .c(_0750_),
    .y(\DFF_523.D )
  );
  al_and3fft _2360_ (
    .a(g1696),
    .b(\DFF_275.Q ),
    .c(g1700),
    .y(g6842)
  );
  al_and3 _2361_ (
    .a(_0541_),
    .b(_0545_),
    .c(_0192_),
    .y(g11206)
  );
  al_and2 _2362_ (
    .a(\DFF_88.Q ),
    .b(g109),
    .y(\DFF_303.D )
  );
  al_aoi21ftf _2363_ (
    .a(g18),
    .b(\DFF_509.Q ),
    .c(_0488_),
    .y(_0751_)
  );
  al_oa21ftf _2364_ (
    .a(\DFF_519.Q ),
    .b(_0751_),
    .c(_0151_),
    .y(_0752_)
  );
  al_aoi21ftf _2365_ (
    .a(\DFF_519.Q ),
    .b(_0751_),
    .c(_0752_),
    .y(\DFF_34.D )
  );
  al_and2 _2366_ (
    .a(\DFF_76.Q ),
    .b(g109),
    .y(\DFF_182.D )
  );
  al_oai21ftt _2367_ (
    .a(\DFF_191.Q ),
    .b(\DFF_518.Q ),
    .c(\DFF_64.Q ),
    .y(_0753_)
  );
  al_aoi21ftf _2368_ (
    .a(_0665_),
    .b(_0753_),
    .c(_0670_),
    .y(\DFF_64.D )
  );
  al_or2ft _2369_ (
    .a(_0555_),
    .b(\DFF_350.D ),
    .y(g10463)
  );
  al_and2ft _2370_ (
    .a(\DFF_278.Q ),
    .b(\DFF_417.Q ),
    .y(_0754_)
  );
  al_nand3 _2371_ (
    .a(\DFF_353.Q ),
    .b(_0754_),
    .c(_0491_),
    .y(_0755_)
  );
  al_ao21 _2372_ (
    .a(_0754_),
    .b(_0491_),
    .c(\DFF_353.Q ),
    .y(_0756_)
  );
  al_nand3 _2373_ (
    .a(_0489_),
    .b(_0755_),
    .c(_0756_),
    .y(_0757_)
  );
  al_aoi21 _2374_ (
    .a(_0651_),
    .b(_0757_),
    .c(\DFF_503.Q ),
    .y(_0758_)
  );
  al_and3 _2375_ (
    .a(\DFF_503.Q ),
    .b(_0651_),
    .c(_0757_),
    .y(_0759_)
  );
  al_mux2l _2376_ (
    .a(_0759_),
    .b(_0758_),
    .s(_0151_),
    .y(\DFF_47.D )
  );
  al_nor2ft _2377_ (
    .a(\DFF_157.Q ),
    .b(\DFF_262.D ),
    .y(\DFF_191.D )
  );
  al_inv _2378_ (
    .a(\DFF_86.Q ),
    .y(_0760_)
  );
  al_nand3fft _2379_ (
    .a(\DFF_135.Q ),
    .b(_0760_),
    .c(_0704_),
    .y(_0761_)
  );
  al_and3fft _2380_ (
    .a(\DFF_261.Q ),
    .b(_0668_),
    .c(\DFF_358.Q ),
    .y(_0762_)
  );
  al_ao21ftt _2381_ (
    .a(_0669_),
    .b(_0762_),
    .c(\DFF_261.Q ),
    .y(_0763_)
  );
  al_and3 _2382_ (
    .a(g18),
    .b(_0763_),
    .c(_0761_),
    .y(\DFF_261.D )
  );
  al_or2 _2383_ (
    .a(g82),
    .b(\DFF_363.Q ),
    .y(g8352)
  );
  al_ao21 _2384_ (
    .a(\DFF_393.Q ),
    .b(_0454_),
    .c(\DFF_184.Q ),
    .y(_0764_)
  );
  al_and3 _2385_ (
    .a(_0455_),
    .b(_0507_),
    .c(_0764_),
    .y(\DFF_184.D )
  );
  al_and2 _2386_ (
    .a(g109),
    .b(\DFF_438.Q ),
    .y(\DFF_438.D )
  );
  al_and2 _2387_ (
    .a(\DFF_400.Q ),
    .b(g18),
    .y(_0765_)
  );
  al_nor2 _2388_ (
    .a(\DFF_472.Q ),
    .b(\DFF_421.Q ),
    .y(_0766_)
  );
  al_nand3fft _2389_ (
    .a(\DFF_507.Q ),
    .b(\DFF_23.Q ),
    .c(_0766_),
    .y(_0767_)
  );
  al_nor3fft _2390_ (
    .a(_0398_),
    .b(_0767_),
    .c(\DFF_116.D ),
    .y(_0768_)
  );
  al_oai21ftf _2391_ (
    .a(\DFF_420.Q ),
    .b(_0767_),
    .c(g18),
    .y(_0769_)
  );
  al_mux2l _2392_ (
    .a(_0769_),
    .b(_0768_),
    .s(_0765_),
    .y(_0770_)
  );
  al_nor2 _2393_ (
    .a(\DFF_494.Q ),
    .b(\DFF_143.Q ),
    .y(_0771_)
  );
  al_nand2 _2394_ (
    .a(\DFF_494.Q ),
    .b(\DFF_143.Q ),
    .y(_0772_)
  );
  al_nand2ft _2395_ (
    .a(_0771_),
    .b(_0772_),
    .y(_0773_)
  );
  al_nand2ft _2396_ (
    .a(\DFF_90.Q ),
    .b(\DFF_118.Q ),
    .y(_0774_)
  );
  al_and3ftt _2397_ (
    .a(_0653_),
    .b(_0774_),
    .c(_0773_),
    .y(_0775_)
  );
  al_ao21ftt _2398_ (
    .a(_0653_),
    .b(_0774_),
    .c(_0773_),
    .y(_0776_)
  );
  al_nand2ft _2399_ (
    .a(_0775_),
    .b(_0776_),
    .y(_0777_)
  );
  al_mux2l _2400_ (
    .a(_0777_),
    .b(_0770_),
    .s(_0151_),
    .y(_0778_)
  );
  al_aoi21ttf _2401_ (
    .a(_0770_),
    .b(_0777_),
    .c(_0778_),
    .y(\DFF_143.D )
  );
  al_nor2ft _2402_ (
    .a(\DFF_252.Q ),
    .b(\DFF_122.D ),
    .y(\DFF_489.D )
  );
  al_aoi21ftf _2403_ (
    .a(_0357_),
    .b(_0355_),
    .c(\DFF_409.Q ),
    .y(_0779_)
  );
  al_ao21 _2404_ (
    .a(\DFF_19.Q ),
    .b(\DFF_207.Q ),
    .c(\DFF_409.Q ),
    .y(_0780_)
  );
  al_and3 _2405_ (
    .a(_0583_),
    .b(_0780_),
    .c(_0355_),
    .y(_0781_)
  );
  al_mux2l _2406_ (
    .a(_0781_),
    .b(_0779_),
    .s(_0534_),
    .y(\DFF_409.D )
  );
  al_or3 _2407_ (
    .a(g30),
    .b(_0009_),
    .c(\DFF_319.D ),
    .y(g10379)
  );
  al_oa21ftt _2408_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_91.Q ),
    .y(\DFF_91.D )
  );
  al_mux2l _2409_ (
    .a(\DFF_324.Q ),
    .b(_0640_),
    .s(\DFF_174.Q ),
    .y(_0782_)
  );
  al_aoi21ttf _2410_ (
    .a(\DFF_324.Q ),
    .b(_0640_),
    .c(_0782_),
    .y(\DFF_324.D )
  );
  al_oa21ftt _2411_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_49.Q ),
    .y(\DFF_49.D )
  );
  al_aoi21ftf _2412_ (
    .a(g18),
    .b(\DFF_199.Q ),
    .c(_0736_),
    .y(_0783_)
  );
  al_oa21ftf _2413_ (
    .a(\DFF_139.Q ),
    .b(_0783_),
    .c(_0151_),
    .y(_0784_)
  );
  al_aoi21ftf _2414_ (
    .a(\DFF_139.Q ),
    .b(_0783_),
    .c(_0784_),
    .y(\DFF_98.D )
  );
  al_and2 _2415_ (
    .a(\DFF_147.Q ),
    .b(\DFF_296.Q ),
    .y(_0785_)
  );
  al_and2ft _2416_ (
    .a(\DFF_364.Q ),
    .b(\DFF_337.Q ),
    .y(_0786_)
  );
  al_nand2ft _2417_ (
    .a(\DFF_337.Q ),
    .b(\DFF_364.Q ),
    .y(_0787_)
  );
  al_nand2ft _2418_ (
    .a(_0786_),
    .b(_0787_),
    .y(_0788_)
  );
  al_oai21ttf _2419_ (
    .a(_0586_),
    .b(_0785_),
    .c(_0788_),
    .y(_0789_)
  );
  al_nand3fft _2420_ (
    .a(_0586_),
    .b(_0785_),
    .c(_0788_),
    .y(_0790_)
  );
  al_and3 _2421_ (
    .a(g109),
    .b(_0790_),
    .c(_0789_),
    .y(\DFF_296.D )
  );
  al_nand3ftt _2422_ (
    .a(\DFF_310.Q ),
    .b(\DFF_362.Q ),
    .c(\DFF_358.Q ),
    .y(_0791_)
  );
  al_ao21ftf _2423_ (
    .a(\DFF_358.Q ),
    .b(\DFF_310.Q ),
    .c(_0791_),
    .y(_0792_)
  );
  al_oai21ftf _2424_ (
    .a(_0677_),
    .b(_0669_),
    .c(_0792_),
    .y(_0793_)
  );
  al_ao21 _2425_ (
    .a(_0793_),
    .b(_0701_),
    .c(\DFF_358.Q ),
    .y(_0794_)
  );
  al_nand3 _2426_ (
    .a(\DFF_358.Q ),
    .b(_0793_),
    .c(_0701_),
    .y(_0795_)
  );
  al_and3 _2427_ (
    .a(g18),
    .b(_0795_),
    .c(_0794_),
    .y(\DFF_358.D )
  );
  al_or2 _2428_ (
    .a(g82),
    .b(\DFF_496.Q ),
    .y(g8347)
  );
  al_aoi21ftf _2429_ (
    .a(g18),
    .b(\DFF_374.Q ),
    .c(_0651_),
    .y(_0796_)
  );
  al_inv _2430_ (
    .a(\DFF_273.Q ),
    .y(_0797_)
  );
  al_mux2l _2431_ (
    .a(_0797_),
    .b(_0796_),
    .s(_0151_),
    .y(_0798_)
  );
  al_aoi21ftf _2432_ (
    .a(\DFF_273.Q ),
    .b(_0796_),
    .c(_0798_),
    .y(\DFF_277.D )
  );
  al_and2 _2433_ (
    .a(g109),
    .b(\DFF_232.Q ),
    .y(\DFF_232.D )
  );
  al_and2 _2434_ (
    .a(\DFF_243.Q ),
    .b(_0486_),
    .y(\DFF_243.D )
  );
  al_and2 _2435_ (
    .a(g109),
    .b(\DFF_315.Q ),
    .y(\DFF_118.D )
  );
  al_nor2ft _2436_ (
    .a(\DFF_385.Q ),
    .b(\DFF_122.D ),
    .y(\DFF_330.D )
  );
  al_and2 _2437_ (
    .a(g109),
    .b(\DFF_468.Q ),
    .y(\DFF_468.D )
  );
  al_ao21 _2438_ (
    .a(\DFF_523.Q ),
    .b(_0749_),
    .c(\DFF_332.Q ),
    .y(_0799_)
  );
  al_and3 _2439_ (
    .a(_0639_),
    .b(_0598_),
    .c(_0799_),
    .y(\DFF_332.D )
  );
  al_nand3fft _2440_ (
    .a(\DFF_358.Q ),
    .b(\DFF_135.Q ),
    .c(_0396_),
    .y(_0800_)
  );
  al_ao21 _2441_ (
    .a(_0677_),
    .b(_0701_),
    .c(\DFF_43.Q ),
    .y(_0801_)
  );
  al_nand3 _2442_ (
    .a(\DFF_43.Q ),
    .b(_0677_),
    .c(_0701_),
    .y(_0802_)
  );
  al_and3 _2443_ (
    .a(_0800_),
    .b(_0802_),
    .c(_0801_),
    .y(\DFF_43.D )
  );
  al_and2ft _2444_ (
    .a(\DFF_158.Q ),
    .b(\DFF_31.Q ),
    .y(_0803_)
  );
  al_ao21ttf _2445_ (
    .a(_0754_),
    .b(_0803_),
    .c(\DFF_145.Q ),
    .y(_0804_)
  );
  al_nand3ftt _2446_ (
    .a(\DFF_145.Q ),
    .b(_0754_),
    .c(_0803_),
    .y(_0805_)
  );
  al_ao21 _2447_ (
    .a(_0805_),
    .b(_0804_),
    .c(g18),
    .y(_0806_)
  );
  al_nand3 _2448_ (
    .a(_0658_),
    .b(_0601_),
    .c(_0806_),
    .y(_0807_)
  );
  al_ao21 _2449_ (
    .a(_0601_),
    .b(_0806_),
    .c(_0658_),
    .y(_0808_)
  );
  al_and3 _2450_ (
    .a(g109),
    .b(_0807_),
    .c(_0808_),
    .y(\DFF_235.D )
  );
  al_nand2 _2451_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .y(_0809_)
  );
  al_and3fft _2452_ (
    .a(\DFF_471.D ),
    .b(_0635_),
    .c(_0809_),
    .y(\DFF_372.D )
  );
  al_ao21ftf _2453_ (
    .a(g18),
    .b(\DFF_186.Q ),
    .c(_0498_),
    .y(\DFF_356.D )
  );
  al_aoi21 _2454_ (
    .a(\DFF_490.Q ),
    .b(\DFF_356.D ),
    .c(_0151_),
    .y(_0810_)
  );
  al_oa21 _2455_ (
    .a(\DFF_490.Q ),
    .b(\DFF_356.D ),
    .c(_0810_),
    .y(\DFF_190.D )
  );
  al_and2 _2456_ (
    .a(g109),
    .b(\DFF_169.Q ),
    .y(\DFF_90.D )
  );
  al_inv _2457_ (
    .a(\DFF_362.Q ),
    .y(_0811_)
  );
  al_nand3 _2458_ (
    .a(\DFF_362.Q ),
    .b(\DFF_358.Q ),
    .c(\DFF_310.Q ),
    .y(_0812_)
  );
  al_nand3 _2459_ (
    .a(_0683_),
    .b(_0812_),
    .c(_0703_),
    .y(_0813_)
  );
  al_ao21ttf _2460_ (
    .a(_0813_),
    .b(_0701_),
    .c(_0800_),
    .y(_0814_)
  );
  al_mux2l _2461_ (
    .a(\DFF_362.Q ),
    .b(_0814_),
    .s(_0489_),
    .y(_0815_)
  );
  al_aoi21ftf _2462_ (
    .a(_0811_),
    .b(_0814_),
    .c(_0815_),
    .y(\DFF_362.D )
  );
  al_nor3fft _2463_ (
    .a(\DFF_97.Q ),
    .b(\DFF_306.Q ),
    .c(_0575_),
    .y(_0816_)
  );
  al_nand3fft _2464_ (
    .a(\DFF_165.Q ),
    .b(\DFF_277.Q ),
    .c(_0816_),
    .y(_0817_)
  );
  al_nor3fft _2465_ (
    .a(\DFF_172.Q ),
    .b(\DFF_201.Q ),
    .c(_0656_),
    .y(_0818_)
  );
  al_inv _2466_ (
    .a(\DFF_98.Q ),
    .y(_0819_)
  );
  al_and2ft _2467_ (
    .a(\DFF_95.Q ),
    .b(\DFF_519.Q ),
    .y(_0820_)
  );
  al_and3ftt _2468_ (
    .a(\DFF_139.Q ),
    .b(\DFF_437.Q ),
    .c(_0820_),
    .y(_0821_)
  );
  al_nand3fft _2469_ (
    .a(_0819_),
    .b(_0797_),
    .c(_0821_),
    .y(_0822_)
  );
  al_nor3ftt _2470_ (
    .a(_0818_),
    .b(_0822_),
    .c(_0817_),
    .y(_0823_)
  );
  al_mux2l _2471_ (
    .a(\DFF_29.Q ),
    .b(_0823_),
    .s(_0151_),
    .y(\DFF_29.D )
  );
  al_aoi21 _2472_ (
    .a(\DFF_112.Q ),
    .b(\DFF_407.Q ),
    .c(\DFF_149.Q ),
    .y(_0824_)
  );
  al_and3fft _2473_ (
    .a(_0824_),
    .b(_0447_),
    .c(_0452_),
    .y(\DFF_149.D )
  );
  al_and2 _2474_ (
    .a(\DFF_67.Q ),
    .b(g109),
    .y(\DFF_125.D )
  );
  al_and2 _2475_ (
    .a(\DFF_83.Q ),
    .b(_0486_),
    .y(\DFF_83.D )
  );
  al_ao21ftf _2476_ (
    .a(g18),
    .b(\DFF_211.Q ),
    .c(_0728_),
    .y(\DFF_246.D )
  );
  al_aoi21 _2477_ (
    .a(\DFF_382.Q ),
    .b(\DFF_246.D ),
    .c(_0151_),
    .y(_0825_)
  );
  al_oa21 _2478_ (
    .a(\DFF_382.Q ),
    .b(\DFF_246.D ),
    .c(_0825_),
    .y(\DFF_474.D )
  );
  al_and2 _2479_ (
    .a(g109),
    .b(\DFF_517.Q ),
    .y(\DFF_517.D )
  );
  al_and2ft _2480_ (
    .a(\DFF_141.Q ),
    .b(\DFF_352.Q ),
    .y(_0826_)
  );
  al_nand2ft _2481_ (
    .a(\DFF_352.Q ),
    .b(\DFF_141.Q ),
    .y(_0827_)
  );
  al_aoi21ftf _2482_ (
    .a(_0826_),
    .b(_0827_),
    .c(_0647_),
    .y(\DFF_141.D )
  );
  al_mux2h _2483_ (
    .a(\DFF_361.Q ),
    .b(_0636_),
    .s(_0530_),
    .y(_0828_)
  );
  al_aoi21ftf _2484_ (
    .a(_0572_),
    .b(_0411_),
    .c(_0828_),
    .y(\DFF_361.D )
  );
  al_mux2l _2485_ (
    .a(_0570_),
    .b(_0569_),
    .s(\DFF_207.Q ),
    .y(_0829_)
  );
  al_or3fft _2486_ (
    .a(\DFF_19.Q ),
    .b(\DFF_207.Q ),
    .c(_0569_),
    .y(_0830_)
  );
  al_and3fft _2487_ (
    .a(_0534_),
    .b(_0829_),
    .c(_0830_),
    .y(\DFF_207.D )
  );
  al_aoi21ftf _2488_ (
    .a(g18),
    .b(\DFF_495.Q ),
    .c(_0708_),
    .y(_0831_)
  );
  al_mux2l _2489_ (
    .a(_0819_),
    .b(_0831_),
    .s(_0151_),
    .y(_0832_)
  );
  al_aoi21ftf _2490_ (
    .a(\DFF_98.Q ),
    .b(_0831_),
    .c(_0832_),
    .y(\DFF_172.D )
  );
  al_oa21 _2491_ (
    .a(\DFF_112.Q ),
    .b(\DFF_407.Q ),
    .c(_0452_),
    .y(_0833_)
  );
  al_aoi21ttf _2492_ (
    .a(\DFF_112.Q ),
    .b(\DFF_407.Q ),
    .c(_0833_),
    .y(\DFF_407.D )
  );
  al_and3ftt _2493_ (
    .a(\DFF_126.Q ),
    .b(\DFF_417.Q ),
    .c(g109),
    .y(\DFF_417.D )
  );
  al_aoi21 _2494_ (
    .a(_0811_),
    .b(_0701_),
    .c(_0489_),
    .y(_0834_)
  );
  al_oa21 _2495_ (
    .a(\DFF_310.Q ),
    .b(_0701_),
    .c(_0834_),
    .y(\DFF_310.D )
  );
  al_and2 _2496_ (
    .a(\DFF_185.Q ),
    .b(g109),
    .y(\DFF_163.D )
  );
  al_nor2ft _2497_ (
    .a(\DFF_489.Q ),
    .b(\DFF_122.D ),
    .y(\DFF_352.D )
  );
  al_and2 _2498_ (
    .a(\DFF_255.Q ),
    .b(_0548_),
    .y(_0835_)
  );
  al_ao21 _2499_ (
    .a(\DFF_12.Q ),
    .b(\DFF_264.Q ),
    .c(\DFF_255.Q ),
    .y(_0836_)
  );
  al_and3 _2500_ (
    .a(_0547_),
    .b(_0836_),
    .c(_0355_),
    .y(_0837_)
  );
  al_mux2l _2501_ (
    .a(_0837_),
    .b(_0835_),
    .s(_0550_),
    .y(\DFF_255.D )
  );
  al_or3 _2502_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_173.Q ),
    .y(_0838_)
  );
  al_mux2h _2503_ (
    .a(\DFF_515.Q ),
    .b(_0635_),
    .s(_0838_),
    .y(\DFF_515.D )
  );
  al_oai21ftf _2504_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_287.Q ),
    .y(\DFF_287.D )
  );
  al_oa21ftf _2505_ (
    .a(\DFF_0.Q ),
    .b(_0443_),
    .c(_0151_),
    .y(_0839_)
  );
  al_nor3fft _2506_ (
    .a(\DFF_510.Q ),
    .b(\DFF_0.Q ),
    .c(_0443_),
    .y(_0840_)
  );
  al_ao21 _2507_ (
    .a(\DFF_202.Q ),
    .b(_0839_),
    .c(_0840_),
    .y(\DFF_202.D )
  );
  al_inv _2508_ (
    .a(_0635_),
    .y(_0841_)
  );
  al_nand3 _2509_ (
    .a(_0635_),
    .b(_0734_),
    .c(_0740_),
    .y(_0842_)
  );
  al_aoi21ftf _2510_ (
    .a(\DFF_516.Q ),
    .b(_0841_),
    .c(_0842_),
    .y(\DFF_516.D )
  );
  al_oa21ftf _2511_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_266.Q ),
    .y(_0843_)
  );
  al_nand2ft _2512_ (
    .a(\DFF_255.Q ),
    .b(\DFF_152.Q ),
    .y(_0844_)
  );
  al_and3fft _2513_ (
    .a(\DFF_12.Q ),
    .b(_0844_),
    .c(\DFF_264.Q ),
    .y(_0845_)
  );
  al_and2 _2514_ (
    .a(\DFF_245.Q ),
    .b(_0845_),
    .y(_0846_)
  );
  al_or2 _2515_ (
    .a(\DFF_245.Q ),
    .b(_0845_),
    .y(_0847_)
  );
  al_nand2ft _2516_ (
    .a(_0846_),
    .b(_0847_),
    .y(_0848_)
  );
  al_nand3 _2517_ (
    .a(\DFF_183.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_0849_)
  );
  al_ao21ftf _2518_ (
    .a(_0848_),
    .b(_0355_),
    .c(_0849_),
    .y(_0850_)
  );
  al_or3 _2519_ (
    .a(\DFF_12.Q ),
    .b(\DFF_264.Q ),
    .c(_0844_),
    .y(_0851_)
  );
  al_or2 _2520_ (
    .a(\DFF_529.Q ),
    .b(_0851_),
    .y(_0852_)
  );
  al_and2 _2521_ (
    .a(\DFF_529.Q ),
    .b(_0851_),
    .y(_0853_)
  );
  al_nand2ft _2522_ (
    .a(_0853_),
    .b(_0852_),
    .y(_0854_)
  );
  al_nand3ftt _2523_ (
    .a(\DFF_175.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_0855_)
  );
  al_ao21ftf _2524_ (
    .a(_0854_),
    .b(_0355_),
    .c(_0855_),
    .y(_0856_)
  );
  al_and2 _2525_ (
    .a(_0850_),
    .b(_0856_),
    .y(_0857_)
  );
  al_nor2 _2526_ (
    .a(_0850_),
    .b(_0856_),
    .y(_0858_)
  );
  al_nand3 _2527_ (
    .a(\DFF_239.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_0859_)
  );
  al_nand3ftt _2528_ (
    .a(\DFF_152.Q ),
    .b(\DFF_459.Q ),
    .c(_0546_),
    .y(_0860_)
  );
  al_ao21ftt _2529_ (
    .a(\DFF_152.Q ),
    .b(_0546_),
    .c(\DFF_459.Q ),
    .y(_0861_)
  );
  al_nand3 _2530_ (
    .a(_0860_),
    .b(_0861_),
    .c(_0355_),
    .y(_0862_)
  );
  al_nand2ft _2531_ (
    .a(\DFF_264.Q ),
    .b(\DFF_12.Q ),
    .y(_0863_)
  );
  al_and3fft _2532_ (
    .a(\DFF_152.Q ),
    .b(_0863_),
    .c(\DFF_255.Q ),
    .y(_0864_)
  );
  al_and2 _2533_ (
    .a(\DFF_221.Q ),
    .b(_0864_),
    .y(_0865_)
  );
  al_or2 _2534_ (
    .a(\DFF_221.Q ),
    .b(_0864_),
    .y(_0866_)
  );
  al_nand2ft _2535_ (
    .a(_0865_),
    .b(_0866_),
    .y(_0867_)
  );
  al_nand3 _2536_ (
    .a(\DFF_65.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_0868_)
  );
  al_ao21ftf _2537_ (
    .a(_0867_),
    .b(_0355_),
    .c(_0868_),
    .y(_0869_)
  );
  al_or3fft _2538_ (
    .a(_0859_),
    .b(_0862_),
    .c(_0869_),
    .y(_0870_)
  );
  al_ao21ttf _2539_ (
    .a(_0859_),
    .b(_0862_),
    .c(_0869_),
    .y(_0871_)
  );
  al_and2 _2540_ (
    .a(_0871_),
    .b(_0870_),
    .y(_0872_)
  );
  al_oa21 _2541_ (
    .a(_0857_),
    .b(_0858_),
    .c(_0872_),
    .y(_0873_)
  );
  al_nand2 _2542_ (
    .a(_0871_),
    .b(_0870_),
    .y(_0874_)
  );
  al_and3fft _2543_ (
    .a(_0857_),
    .b(_0858_),
    .c(_0874_),
    .y(_0875_)
  );
  al_nand3 _2544_ (
    .a(\DFF_225.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_0876_)
  );
  al_or2 _2545_ (
    .a(\DFF_152.Q ),
    .b(\DFF_255.Q ),
    .y(_0877_)
  );
  al_nor3fft _2546_ (
    .a(\DFF_12.Q ),
    .b(\DFF_264.Q ),
    .c(_0877_),
    .y(_0878_)
  );
  al_and2 _2547_ (
    .a(\DFF_151.Q ),
    .b(_0878_),
    .y(_0879_)
  );
  al_or2 _2548_ (
    .a(\DFF_151.Q ),
    .b(_0878_),
    .y(_0880_)
  );
  al_nand3ftt _2549_ (
    .a(_0879_),
    .b(_0880_),
    .c(_0355_),
    .y(_0881_)
  );
  al_or3 _2550_ (
    .a(\DFF_430.Q ),
    .b(_0863_),
    .c(_0877_),
    .y(_0882_)
  );
  al_mux2h _2551_ (
    .a(_0863_),
    .b(_0877_),
    .s(\DFF_430.Q ),
    .y(_0883_)
  );
  al_or2ft _2552_ (
    .a(_0882_),
    .b(_0883_),
    .y(_0884_)
  );
  al_inv _2553_ (
    .a(\DFF_41.Q ),
    .y(_0885_)
  );
  al_nand3 _2554_ (
    .a(_0885_),
    .b(_0354_),
    .c(_0568_),
    .y(_0886_)
  );
  al_ao21ftf _2555_ (
    .a(_0884_),
    .b(_0355_),
    .c(_0886_),
    .y(_0887_)
  );
  al_and3 _2556_ (
    .a(_0876_),
    .b(_0881_),
    .c(_0887_),
    .y(_0888_)
  );
  al_ao21 _2557_ (
    .a(_0876_),
    .b(_0881_),
    .c(_0887_),
    .y(_0889_)
  );
  al_nand2ft _2558_ (
    .a(_0888_),
    .b(_0889_),
    .y(_0890_)
  );
  al_and3fft _2559_ (
    .a(\DFF_12.Q ),
    .b(\DFF_152.Q ),
    .c(\DFF_255.Q ),
    .y(_0891_)
  );
  al_and3 _2560_ (
    .a(\DFF_264.Q ),
    .b(\DFF_51.Q ),
    .c(_0891_),
    .y(_0892_)
  );
  al_ao21 _2561_ (
    .a(\DFF_264.Q ),
    .b(_0891_),
    .c(\DFF_51.Q ),
    .y(_0893_)
  );
  al_nand2ft _2562_ (
    .a(_0892_),
    .b(_0893_),
    .y(_0894_)
  );
  al_nand3ftt _2563_ (
    .a(\DFF_467.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_0895_)
  );
  al_ao21ttf _2564_ (
    .a(_0894_),
    .b(_0355_),
    .c(_0895_),
    .y(_0896_)
  );
  al_and3ftt _2565_ (
    .a(\DFF_264.Q ),
    .b(\DFF_329.Q ),
    .c(_0891_),
    .y(_0897_)
  );
  al_ao21ftt _2566_ (
    .a(\DFF_264.Q ),
    .b(_0891_),
    .c(\DFF_329.Q ),
    .y(_0898_)
  );
  al_nand2ft _2567_ (
    .a(_0897_),
    .b(_0898_),
    .y(_0899_)
  );
  al_nand3 _2568_ (
    .a(\DFF_478.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_0900_)
  );
  al_ao21ftf _2569_ (
    .a(_0899_),
    .b(_0355_),
    .c(_0900_),
    .y(_0901_)
  );
  al_nand2ft _2570_ (
    .a(_0901_),
    .b(_0896_),
    .y(_0902_)
  );
  al_nand2ft _2571_ (
    .a(_0896_),
    .b(_0901_),
    .y(_0903_)
  );
  al_and3 _2572_ (
    .a(_0902_),
    .b(_0903_),
    .c(_0890_),
    .y(_0904_)
  );
  al_ao21 _2573_ (
    .a(_0902_),
    .b(_0903_),
    .c(_0890_),
    .y(_0905_)
  );
  al_nand2ft _2574_ (
    .a(_0904_),
    .b(_0905_),
    .y(_0906_)
  );
  al_nand3fft _2575_ (
    .a(_0873_),
    .b(_0875_),
    .c(_0906_),
    .y(_0907_)
  );
  al_and3fft _2576_ (
    .a(_0857_),
    .b(_0858_),
    .c(_0872_),
    .y(_0908_)
  );
  al_oa21 _2577_ (
    .a(_0857_),
    .b(_0858_),
    .c(_0874_),
    .y(_0909_)
  );
  al_and2ft _2578_ (
    .a(_0904_),
    .b(_0905_),
    .y(_0910_)
  );
  al_nand3fft _2579_ (
    .a(_0908_),
    .b(_0909_),
    .c(_0910_),
    .y(_0911_)
  );
  al_or3 _2580_ (
    .a(\DFF_379.Q ),
    .b(_0844_),
    .c(_0863_),
    .y(_0912_)
  );
  al_mux2h _2581_ (
    .a(_0844_),
    .b(_0863_),
    .s(\DFF_379.Q ),
    .y(_0913_)
  );
  al_or2ft _2582_ (
    .a(_0912_),
    .b(_0913_),
    .y(_0914_)
  );
  al_nand3 _2583_ (
    .a(\DFF_2.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_0915_)
  );
  al_ao21ttf _2584_ (
    .a(_0914_),
    .b(_0355_),
    .c(_0915_),
    .y(_0916_)
  );
  al_inv _2585_ (
    .a(_0916_),
    .y(_0917_)
  );
  al_nand3 _2586_ (
    .a(_0917_),
    .b(_0907_),
    .c(_0911_),
    .y(_0918_)
  );
  al_nand3fft _2587_ (
    .a(_0873_),
    .b(_0875_),
    .c(_0910_),
    .y(_0919_)
  );
  al_nand3fft _2588_ (
    .a(_0908_),
    .b(_0909_),
    .c(_0906_),
    .y(_0920_)
  );
  al_nand3 _2589_ (
    .a(_0916_),
    .b(_0920_),
    .c(_0919_),
    .y(_0921_)
  );
  al_and3fft _2590_ (
    .a(\DFF_12.Q ),
    .b(_0877_),
    .c(\DFF_264.Q ),
    .y(_0922_)
  );
  al_nor2 _2591_ (
    .a(\DFF_379.Q ),
    .b(\DFF_210.Q ),
    .y(_0923_)
  );
  al_nand3fft _2592_ (
    .a(\DFF_522.Q ),
    .b(\DFF_51.Q ),
    .c(_0923_),
    .y(_0924_)
  );
  al_or3 _2593_ (
    .a(\DFF_430.Q ),
    .b(\DFF_459.Q ),
    .c(\DFF_205.Q ),
    .y(_0925_)
  );
  al_nor2 _2594_ (
    .a(\DFF_529.Q ),
    .b(\DFF_329.Q ),
    .y(_0926_)
  );
  al_nand3fft _2595_ (
    .a(\DFF_151.Q ),
    .b(\DFF_203.Q ),
    .c(_0926_),
    .y(_0927_)
  );
  al_or3 _2596_ (
    .a(\DFF_245.Q ),
    .b(\DFF_221.Q ),
    .c(_0927_),
    .y(_0928_)
  );
  al_or3 _2597_ (
    .a(_0924_),
    .b(_0925_),
    .c(_0928_),
    .y(_0929_)
  );
  al_nand3fft _2598_ (
    .a(\DFF_475.Q ),
    .b(\DFF_447.Q ),
    .c(_0929_),
    .y(_0930_)
  );
  al_ao21ttf _2599_ (
    .a(\DFF_475.Q ),
    .b(\DFF_447.Q ),
    .c(_0930_),
    .y(_0931_)
  );
  al_and2 _2600_ (
    .a(_0922_),
    .b(_0931_),
    .y(_0932_)
  );
  al_or2 _2601_ (
    .a(_0922_),
    .b(_0931_),
    .y(_0933_)
  );
  al_nand2ft _2602_ (
    .a(_0932_),
    .b(_0933_),
    .y(_0934_)
  );
  al_nand3 _2603_ (
    .a(_0358_),
    .b(_0354_),
    .c(_0568_),
    .y(_0935_)
  );
  al_ao21ftf _2604_ (
    .a(_0934_),
    .b(_0355_),
    .c(_0935_),
    .y(_0936_)
  );
  al_aoi21 _2605_ (
    .a(_0918_),
    .b(_0921_),
    .c(_0936_),
    .y(_0937_)
  );
  al_nand3 _2606_ (
    .a(_0936_),
    .b(_0918_),
    .c(_0921_),
    .y(_0938_)
  );
  al_nand2 _2607_ (
    .a(_0006_),
    .b(_0938_),
    .y(_0939_)
  );
  al_mux2l _2608_ (
    .a(_0937_),
    .b(_0939_),
    .s(_0843_),
    .y(\DFF_266.D )
  );
  al_nand2 _2609_ (
    .a(_0467_),
    .b(_0480_),
    .y(_0940_)
  );
  al_or3fft _2610_ (
    .a(_0465_),
    .b(_0468_),
    .c(_0940_),
    .y(_0941_)
  );
  al_aoi21ftf _2611_ (
    .a(_0475_),
    .b(\DFF_212.Q ),
    .c(_0941_),
    .y(_0942_)
  );
  al_inv _2612_ (
    .a(\DFF_223.Q ),
    .y(_0943_)
  );
  al_ao21ttf _2613_ (
    .a(_0943_),
    .b(_0674_),
    .c(_0673_),
    .y(_0944_)
  );
  al_nand3 _2614_ (
    .a(_0673_),
    .b(_0463_),
    .c(_0944_),
    .y(_0945_)
  );
  al_nor2 _2615_ (
    .a(_0671_),
    .b(_0944_),
    .y(_0946_)
  );
  al_mux2l _2616_ (
    .a(_0945_),
    .b(_0942_),
    .s(_0946_),
    .y(_0947_)
  );
  al_or2 _2617_ (
    .a(_0466_),
    .b(_0947_),
    .y(_0948_)
  );
  al_aoi21ftf _2618_ (
    .a(\DFF_271.Q ),
    .b(_0947_),
    .c(_0513_),
    .y(_0949_)
  );
  al_aoi21ftt _2619_ (
    .a(\DFF_369.Q ),
    .b(\DFF_302.Q ),
    .c(_0458_),
    .y(_0950_)
  );
  al_and3 _2620_ (
    .a(_0516_),
    .b(_0950_),
    .c(_0483_),
    .y(_0951_)
  );
  al_ao21 _2621_ (
    .a(_0948_),
    .b(_0949_),
    .c(_0951_),
    .y(\DFF_271.D )
  );
  al_nand3 _2622_ (
    .a(\DFF_379.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_0952_)
  );
  al_ao21ttf _2623_ (
    .a(\DFF_245.Q ),
    .b(_0355_),
    .c(_0952_),
    .y(\DFF_379.D )
  );
  al_inv _2624_ (
    .a(\DFF_261.Q ),
    .y(_0953_)
  );
  al_and3fft _2625_ (
    .a(_0953_),
    .b(_0669_),
    .c(_0706_),
    .y(_0954_)
  );
  al_or3fft _2626_ (
    .a(\DFF_86.Q ),
    .b(_0800_),
    .c(_0954_),
    .y(_0955_)
  );
  al_ao21ttf _2627_ (
    .a(\DFF_427.Q ),
    .b(_0954_),
    .c(_0955_),
    .y(\DFF_86.D )
  );
  al_and2 _2628_ (
    .a(g109),
    .b(_0589_),
    .y(_0956_)
  );
  al_nand3ftt _2629_ (
    .a(\DFF_197.Q ),
    .b(g109),
    .c(_0589_),
    .y(_0957_)
  );
  al_mux2h _2630_ (
    .a(\DFF_474.Q ),
    .b(_0956_),
    .s(_0957_),
    .y(\DFF_197.D )
  );
  al_and2ft _2631_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .y(_0958_)
  );
  al_nand3ftt _2632_ (
    .a(\DFF_113.Q ),
    .b(\DFF_241.Q ),
    .c(_0958_),
    .y(_0959_)
  );
  al_mux2l _2633_ (
    .a(_0151_),
    .b(\DFF_228.D ),
    .s(_0959_),
    .y(_0960_)
  );
  al_ao21ftt _2634_ (
    .a(_0958_),
    .b(\DFF_162.Q ),
    .c(_0960_),
    .y(\DFF_162.D )
  );
  al_and2 _2635_ (
    .a(g109),
    .b(_0656_),
    .y(_0961_)
  );
  al_nand3ftt _2636_ (
    .a(\DFF_140.Q ),
    .b(g109),
    .c(_0656_),
    .y(_0962_)
  );
  al_mux2h _2637_ (
    .a(\DFF_315.Q ),
    .b(_0961_),
    .s(_0962_),
    .y(\DFF_140.D )
  );
  al_nand3 _2638_ (
    .a(\DFF_3.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_0963_)
  );
  al_ao21ttf _2639_ (
    .a(\DFF_406.Q ),
    .b(_0355_),
    .c(_0963_),
    .y(\DFF_3.D )
  );
  al_or3 _2640_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_402.Q ),
    .y(_0964_)
  );
  al_mux2h _2641_ (
    .a(\DFF_497.Q ),
    .b(_0635_),
    .s(_0964_),
    .y(\DFF_497.D )
  );
  al_nand3ftt _2642_ (
    .a(\DFF_485.Q ),
    .b(g109),
    .c(_0589_),
    .y(_0965_)
  );
  al_mux2h _2643_ (
    .a(\DFF_307.Q ),
    .b(_0956_),
    .s(_0965_),
    .y(\DFF_485.D )
  );
  al_nand2 _2644_ (
    .a(\DFF_323.Q ),
    .b(\DFF_320.Q ),
    .y(_0966_)
  );
  al_ao21 _2645_ (
    .a(\DFF_323.Q ),
    .b(\DFF_320.Q ),
    .c(\DFF_501.Q ),
    .y(_0967_)
  );
  al_mux2h _2646_ (
    .a(\DFF_59.Q ),
    .b(_0966_),
    .s(_0967_),
    .y(\DFF_501.D )
  );
  al_oa21ftt _2647_ (
    .a(\DFF_372.Q ),
    .b(g1696),
    .c(\DFF_16.Q ),
    .y(_0968_)
  );
  al_ao21 _2648_ (
    .a(\DFF_283.Q ),
    .b(_0958_),
    .c(_0968_),
    .y(\DFF_16.D )
  );
  al_nand3ftt _2649_ (
    .a(\DFF_511.Q ),
    .b(g109),
    .c(_0589_),
    .y(_0969_)
  );
  al_mux2h _2650_ (
    .a(\DFF_220.Q ),
    .b(_0956_),
    .s(_0969_),
    .y(\DFF_511.D )
  );
  al_and2ft _2651_ (
    .a(\DFF_417.Q ),
    .b(\DFF_278.Q ),
    .y(_0970_)
  );
  al_nand3 _2652_ (
    .a(\DFF_517.Q ),
    .b(_0970_),
    .c(_0803_),
    .y(_0971_)
  );
  al_ao21 _2653_ (
    .a(_0970_),
    .b(_0803_),
    .c(\DFF_517.Q ),
    .y(_0972_)
  );
  al_ao21 _2654_ (
    .a(_0971_),
    .b(_0972_),
    .c(_0841_),
    .y(_0973_)
  );
  al_aoi21ftf _2655_ (
    .a(\DFF_435.Q ),
    .b(_0841_),
    .c(_0973_),
    .y(\DFF_435.D )
  );
  al_nand3ftt _2656_ (
    .a(_0368_),
    .b(_0357_),
    .c(_0355_),
    .y(_0974_)
  );
  al_nand3ftt _2657_ (
    .a(_0357_),
    .b(\DFF_265.Q ),
    .c(_0355_),
    .y(_0975_)
  );
  al_nand3 _2658_ (
    .a(\DFF_124.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_0976_)
  );
  al_nand3 _2659_ (
    .a(_0976_),
    .b(_0974_),
    .c(_0975_),
    .y(\DFF_124.D )
  );
  al_nand2 _2660_ (
    .a(_0536_),
    .b(\DFF_37.D ),
    .y(_0977_)
  );
  al_and3 _2661_ (
    .a(\DFF_338.Q ),
    .b(_0536_),
    .c(\DFF_37.D ),
    .y(_0978_)
  );
  al_ao21 _2662_ (
    .a(\DFF_454.Q ),
    .b(_0977_),
    .c(_0978_),
    .y(\DFF_454.D )
  );
  al_ao21 _2663_ (
    .a(\DFF_323.Q ),
    .b(\DFF_320.Q ),
    .c(\DFF_131.Q ),
    .y(_0979_)
  );
  al_mux2h _2664_ (
    .a(\DFF_268.Q ),
    .b(_0966_),
    .s(_0979_),
    .y(\DFF_131.D )
  );
  al_nand3 _2665_ (
    .a(_0635_),
    .b(_0498_),
    .c(_0502_),
    .y(_0980_)
  );
  al_aoi21ftf _2666_ (
    .a(\DFF_374.Q ),
    .b(_0841_),
    .c(_0980_),
    .y(\DFF_374.D )
  );
  al_inv _2667_ (
    .a(\DFF_241.Q ),
    .y(_0981_)
  );
  al_and3fft _2668_ (
    .a(\DFF_113.Q ),
    .b(_0602_),
    .c(_0981_),
    .y(_0982_)
  );
  al_and3ftt _2669_ (
    .a(\DFF_113.Q ),
    .b(\DFF_241.Q ),
    .c(g109),
    .y(_0983_)
  );
  al_ao21 _2670_ (
    .a(_0983_),
    .b(\DFF_228.D ),
    .c(_0982_),
    .y(_0984_)
  );
  al_nand2 _2671_ (
    .a(_0635_),
    .b(_0984_),
    .y(_0985_)
  );
  al_ao21ftf _2672_ (
    .a(_0635_),
    .b(\DFF_206.Q ),
    .c(_0985_),
    .y(\DFF_206.D )
  );
  al_nand3ftt _2673_ (
    .a(\DFF_123.Q ),
    .b(g109),
    .c(_0589_),
    .y(_0986_)
  );
  al_mux2h _2674_ (
    .a(\DFF_314.Q ),
    .b(_0956_),
    .s(_0986_),
    .y(\DFF_123.D )
  );
  al_nand2ft _2675_ (
    .a(g85),
    .b(g86),
    .y(_0987_)
  );
  al_ao21ttf _2676_ (
    .a(g85),
    .b(\DFF_274.Q ),
    .c(_0987_),
    .y(\DFF_274.D )
  );
  al_oa21ftt _2677_ (
    .a(\DFF_372.Q ),
    .b(g1696),
    .c(\DFF_82.Q ),
    .y(_0988_)
  );
  al_ao21 _2678_ (
    .a(\DFF_308.Q ),
    .b(_0958_),
    .c(_0988_),
    .y(\DFF_82.D )
  );
  al_and3 _2679_ (
    .a(\DFF_248.Q ),
    .b(_0536_),
    .c(\DFF_37.D ),
    .y(_0989_)
  );
  al_ao21 _2680_ (
    .a(\DFF_351.Q ),
    .b(_0977_),
    .c(_0989_),
    .y(\DFF_351.D )
  );
  al_aoi21ftf _2681_ (
    .a(_0944_),
    .b(\DFF_532.Q ),
    .c(_0945_),
    .y(_0990_)
  );
  al_and2 _2682_ (
    .a(\DFF_449.Q ),
    .b(_0990_),
    .y(_0991_)
  );
  al_or2 _2683_ (
    .a(\DFF_449.Q ),
    .b(_0990_),
    .y(_0992_)
  );
  al_nand2ft _2684_ (
    .a(_0991_),
    .b(_0992_),
    .y(_0993_)
  );
  al_ao21 _2685_ (
    .a(_0993_),
    .b(_0513_),
    .c(_0951_),
    .y(\DFF_449.D )
  );
  al_nand3 _2686_ (
    .a(\DFF_204.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_0994_)
  );
  al_ao21ttf _2687_ (
    .a(\DFF_491.Q ),
    .b(_0355_),
    .c(_0994_),
    .y(\DFF_204.D )
  );
  al_nand3 _2688_ (
    .a(\DFF_491.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_0995_)
  );
  al_ao21ttf _2689_ (
    .a(\DFF_419.Q ),
    .b(_0355_),
    .c(_0995_),
    .y(\DFF_491.D )
  );
  al_nand3ftt _2690_ (
    .a(\DFF_456.Q ),
    .b(g109),
    .c(_0656_),
    .y(_0996_)
  );
  al_mux2h _2691_ (
    .a(\DFF_47.Q ),
    .b(_0961_),
    .s(_0996_),
    .y(\DFF_456.D )
  );
  al_nand3 _2692_ (
    .a(\DFF_459.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_0997_)
  );
  al_ao21ttf _2693_ (
    .a(\DFF_221.Q ),
    .b(_0355_),
    .c(_0997_),
    .y(\DFF_459.D )
  );
  al_oa21ftf _2694_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_308.Q ),
    .y(_0998_)
  );
  al_aoi21 _2695_ (
    .a(_0006_),
    .b(_0856_),
    .c(_0998_),
    .y(\DFF_308.D )
  );
  al_aoi21ftf _2696_ (
    .a(_0467_),
    .b(_0474_),
    .c(_0940_),
    .y(_0999_)
  );
  al_nor2ft _2697_ (
    .a(\DFF_373.Q ),
    .b(_0944_),
    .y(_1000_)
  );
  al_mux2l _2698_ (
    .a(_0945_),
    .b(_0999_),
    .s(_1000_),
    .y(_1001_)
  );
  al_nand2 _2699_ (
    .a(\DFF_44.Q ),
    .b(_1001_),
    .y(_1002_)
  );
  al_or2 _2700_ (
    .a(\DFF_44.Q ),
    .b(_1001_),
    .y(_1003_)
  );
  al_ao21ttf _2701_ (
    .a(_1002_),
    .b(_1003_),
    .c(_0513_),
    .y(_1004_)
  );
  al_nand2ft _2702_ (
    .a(_0951_),
    .b(_1004_),
    .y(\DFF_44.D )
  );
  al_ao21ttf _2703_ (
    .a(_0416_),
    .b(_0415_),
    .c(_0636_),
    .y(_1005_)
  );
  al_ao21ttf _2704_ (
    .a(\DFF_480.Q ),
    .b(_0839_),
    .c(_1005_),
    .y(\DFF_480.D )
  );
  al_ao21 _2705_ (
    .a(\DFF_323.Q ),
    .b(\DFF_320.Q ),
    .c(\DFF_272.Q ),
    .y(_1006_)
  );
  al_mux2h _2706_ (
    .a(\DFF_103.Q ),
    .b(_0966_),
    .s(_1006_),
    .y(\DFF_272.D )
  );
  al_or2ft _2707_ (
    .a(_0317_),
    .b(_0316_),
    .y(\DFF_92.D )
  );
  al_inv _2708_ (
    .a(\DFF_521.Q ),
    .y(_1007_)
  );
  al_or3fft _2709_ (
    .a(\DFF_281.Q ),
    .b(_0800_),
    .c(_0954_),
    .y(_1008_)
  );
  al_ao21ftf _2710_ (
    .a(_1007_),
    .b(_0954_),
    .c(_1008_),
    .y(\DFF_281.D )
  );
  al_oai21ftf _2711_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_103.Q ),
    .y(_1009_)
  );
  al_oai21ftf _2712_ (
    .a(_1009_),
    .b(_0596_),
    .c(\DFF_174.Q ),
    .y(\DFF_103.D )
  );
  al_and3 _2713_ (
    .a(\DFF_433.Q ),
    .b(_0536_),
    .c(\DFF_37.D ),
    .y(_1010_)
  );
  al_ao21 _2714_ (
    .a(\DFF_408.Q ),
    .b(_0977_),
    .c(_1010_),
    .y(\DFF_408.D )
  );
  al_inv _2715_ (
    .a(\DFF_339.Q ),
    .y(_1011_)
  );
  al_and3 _2716_ (
    .a(\DFF_223.Q ),
    .b(_0607_),
    .c(_0673_),
    .y(_1012_)
  );
  al_or3fft _2717_ (
    .a(\DFF_373.Q ),
    .b(_0512_),
    .c(_1012_),
    .y(_1013_)
  );
  al_ao21ftf _2718_ (
    .a(_1011_),
    .b(_1012_),
    .c(_1013_),
    .y(\DFF_373.D )
  );
  al_nor3fft _2719_ (
    .a(\DFF_322.Q ),
    .b(\DFF_0.Q ),
    .c(_0443_),
    .y(_1014_)
  );
  al_ao21 _2720_ (
    .a(\DFF_32.Q ),
    .b(_0839_),
    .c(_1014_),
    .y(\DFF_32.D )
  );
  al_oa21ftt _2721_ (
    .a(\DFF_372.Q ),
    .b(g1696),
    .c(\DFF_402.Q ),
    .y(_1015_)
  );
  al_ao21 _2722_ (
    .a(\DFF_79.Q ),
    .b(_0958_),
    .c(_1015_),
    .y(\DFF_402.D )
  );
  al_nand3ftt _2723_ (
    .a(\DFF_520.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1016_)
  );
  al_mux2h _2724_ (
    .a(\DFF_118.Q ),
    .b(_0961_),
    .s(_1016_),
    .y(\DFF_520.D )
  );
  al_inv _2725_ (
    .a(_0006_),
    .y(_1017_)
  );
  al_oa21ftf _2726_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_499.Q ),
    .y(_1018_)
  );
  al_mux2l _2727_ (
    .a(_1017_),
    .b(_0916_),
    .s(_1018_),
    .y(\DFF_499.D )
  );
  al_nand3 _2728_ (
    .a(_0006_),
    .b(_0859_),
    .c(_0862_),
    .y(_1019_)
  );
  al_aoi21ftf _2729_ (
    .a(\DFF_238.Q ),
    .b(_1017_),
    .c(_1019_),
    .y(\DFF_238.D )
  );
  al_or3fft _2730_ (
    .a(\DFF_313.Q ),
    .b(_0512_),
    .c(_1012_),
    .y(_1020_)
  );
  al_ao21ttf _2731_ (
    .a(\DFF_373.Q ),
    .b(_1012_),
    .c(_1020_),
    .y(\DFF_313.D )
  );
  al_nand3ftt _2732_ (
    .a(\DFF_138.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1021_)
  );
  al_mux2h _2733_ (
    .a(\DFF_128.Q ),
    .b(_0961_),
    .s(_1021_),
    .y(\DFF_138.D )
  );
  al_or3 _2734_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_27.Q ),
    .y(_1022_)
  );
  al_mux2h _2735_ (
    .a(\DFF_234.Q ),
    .b(_0635_),
    .s(_1022_),
    .y(\DFF_234.D )
  );
  al_nor3fft _2736_ (
    .a(\DFF_355.Q ),
    .b(\DFF_0.Q ),
    .c(_0443_),
    .y(_1023_)
  );
  al_ao21 _2737_ (
    .a(\DFF_442.Q ),
    .b(_0839_),
    .c(_1023_),
    .y(\DFF_442.D )
  );
  al_nand3 _2738_ (
    .a(\DFF_221.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1024_)
  );
  al_ao21ttf _2739_ (
    .a(\DFF_51.Q ),
    .b(_0355_),
    .c(_1024_),
    .y(\DFF_221.D )
  );
  al_nor2ft _2740_ (
    .a(_0800_),
    .b(_0701_),
    .y(_1025_)
  );
  al_and2 _2741_ (
    .a(\DFF_11.Q ),
    .b(_0686_),
    .y(_1026_)
  );
  al_nand3fft _2742_ (
    .a(_0679_),
    .b(_0692_),
    .c(_1026_),
    .y(_1027_)
  );
  al_oai21ftf _2743_ (
    .a(_0953_),
    .b(_0762_),
    .c(_0669_),
    .y(_1028_)
  );
  al_inv _2744_ (
    .a(_1028_),
    .y(_1029_)
  );
  al_aoi21 _2745_ (
    .a(_0679_),
    .b(_0698_),
    .c(_1029_),
    .y(_1030_)
  );
  al_or2 _2746_ (
    .a(\DFF_427.Q ),
    .b(_1028_),
    .y(_1031_)
  );
  al_ao21ttf _2747_ (
    .a(_1028_),
    .b(_0691_),
    .c(_1031_),
    .y(_1032_)
  );
  al_aoi21 _2748_ (
    .a(_1027_),
    .b(_1030_),
    .c(_1032_),
    .y(_1033_)
  );
  al_nand2 _2749_ (
    .a(\DFF_286.Q ),
    .b(_1033_),
    .y(_1034_)
  );
  al_or2 _2750_ (
    .a(\DFF_286.Q ),
    .b(_1033_),
    .y(_1035_)
  );
  al_nand3 _2751_ (
    .a(_1034_),
    .b(_1035_),
    .c(_1025_),
    .y(_1036_)
  );
  al_ao21ftt _2752_ (
    .a(\DFF_362.Q ),
    .b(\DFF_310.Q ),
    .c(_0677_),
    .y(_1037_)
  );
  al_and3fft _2753_ (
    .a(_0681_),
    .b(_1037_),
    .c(_0800_),
    .y(_1038_)
  );
  al_and2 _2754_ (
    .a(_1038_),
    .b(_0701_),
    .y(_1039_)
  );
  al_nand2ft _2755_ (
    .a(_1039_),
    .b(_1036_),
    .y(\DFF_286.D )
  );
  al_nand2ft _2756_ (
    .a(\DFF_518.Q ),
    .b(\DFF_191.Q ),
    .y(_1040_)
  );
  al_nand2ft _2757_ (
    .a(\DFF_191.Q ),
    .b(\DFF_518.Q ),
    .y(_1041_)
  );
  al_nand3 _2758_ (
    .a(_1040_),
    .b(_1041_),
    .c(_0670_),
    .y(\DFF_518.D )
  );
  al_and2ft _2759_ (
    .a(\DFF_113.Q ),
    .b(\DFF_241.Q ),
    .y(_1042_)
  );
  al_mux2h _2760_ (
    .a(_0151_),
    .b(\DFF_116.D ),
    .s(_1042_),
    .y(_1043_)
  );
  al_inv _2761_ (
    .a(\DFF_113.Q ),
    .y(_1044_)
  );
  al_or3fft _2762_ (
    .a(_0981_),
    .b(_1044_),
    .c(_0645_),
    .y(_1045_)
  );
  al_oai21ftf _2763_ (
    .a(_1045_),
    .b(_1043_),
    .c(_0841_),
    .y(_1046_)
  );
  al_ao21ftf _2764_ (
    .a(_0635_),
    .b(\DFF_288.Q ),
    .c(_1046_),
    .y(\DFF_288.D )
  );
  al_mux2h _2765_ (
    .a(_0151_),
    .b(\DFF_350.D ),
    .s(_1042_),
    .y(_1047_)
  );
  al_or3fft _2766_ (
    .a(_0981_),
    .b(_1044_),
    .c(_0796_),
    .y(_1048_)
  );
  al_oai21ftf _2767_ (
    .a(_1048_),
    .b(_1047_),
    .c(_0841_),
    .y(_1049_)
  );
  al_ao21ftf _2768_ (
    .a(_0635_),
    .b(\DFF_208.Q ),
    .c(_1049_),
    .y(\DFF_208.D )
  );
  al_ao21ftt _2769_ (
    .a(_0478_),
    .b(_0472_),
    .c(_0945_),
    .y(_1050_)
  );
  al_aoi21ftf _2770_ (
    .a(_0944_),
    .b(\DFF_349.Q ),
    .c(_1050_),
    .y(_1051_)
  );
  al_and2 _2771_ (
    .a(\DFF_1.Q ),
    .b(_1051_),
    .y(_1052_)
  );
  al_or2 _2772_ (
    .a(\DFF_1.Q ),
    .b(_1051_),
    .y(_1053_)
  );
  al_nand2ft _2773_ (
    .a(_1052_),
    .b(_1053_),
    .y(_1054_)
  );
  al_ao21 _2774_ (
    .a(_1054_),
    .b(_0513_),
    .c(_0951_),
    .y(\DFF_1.D )
  );
  al_inv _2775_ (
    .a(\DFF_276.Q ),
    .y(_1055_)
  );
  al_ao21ftt _2776_ (
    .a(_0731_),
    .b(_1055_),
    .c(_0512_),
    .y(_1056_)
  );
  al_aoi21 _2777_ (
    .a(\DFF_276.Q ),
    .b(\DFF_168.D ),
    .c(_1056_),
    .y(_1057_)
  );
  al_inv _2778_ (
    .a(\DFF_178.Q ),
    .y(_1058_)
  );
  al_aoi21 _2779_ (
    .a(\DFF_223.Q ),
    .b(\DFF_455.Q ),
    .c(_0517_),
    .y(_1059_)
  );
  al_nand3fft _2780_ (
    .a(\DFF_178.Q ),
    .b(_0458_),
    .c(_1059_),
    .y(_1060_)
  );
  al_ao21ftf _2781_ (
    .a(_1058_),
    .b(_0461_),
    .c(_1060_),
    .y(_1061_)
  );
  al_or3fft _2782_ (
    .a(g109),
    .b(_1061_),
    .c(\DFF_350.D ),
    .y(_1062_)
  );
  al_mux2l _2783_ (
    .a(_0151_),
    .b(\DFF_350.D ),
    .s(_1061_),
    .y(_1063_)
  );
  al_and3 _2784_ (
    .a(_0461_),
    .b(_0674_),
    .c(_1059_),
    .y(_1064_)
  );
  al_aoi21ttf _2785_ (
    .a(_0950_),
    .b(_1064_),
    .c(\DFF_489.D ),
    .y(_1065_)
  );
  al_or3fft _2786_ (
    .a(_1065_),
    .b(_1062_),
    .c(_1063_),
    .y(_1066_)
  );
  al_ao21 _2787_ (
    .a(\DFF_311.Q ),
    .b(_1066_),
    .c(_0514_),
    .y(_1067_)
  );
  al_ao21 _2788_ (
    .a(_0512_),
    .b(_1067_),
    .c(_1057_),
    .y(\DFF_311.D )
  );
  al_nand3 _2789_ (
    .a(\DFF_114.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1068_)
  );
  al_ao21ttf _2790_ (
    .a(\DFF_394.Q ),
    .b(_0355_),
    .c(_1068_),
    .y(\DFF_114.D )
  );
  al_nand2 _2791_ (
    .a(_1028_),
    .b(_0691_),
    .y(_1069_)
  );
  al_or3ftt _2792_ (
    .a(_1028_),
    .b(_0686_),
    .c(_0697_),
    .y(_1070_)
  );
  al_or2 _2793_ (
    .a(\DFF_281.Q ),
    .b(_1028_),
    .y(_1071_)
  );
  al_and3 _2794_ (
    .a(_1069_),
    .b(_1071_),
    .c(_1070_),
    .y(_1072_)
  );
  al_and2 _2795_ (
    .a(_0693_),
    .b(_1072_),
    .y(_1073_)
  );
  al_or2 _2796_ (
    .a(_0693_),
    .b(_1072_),
    .y(_1074_)
  );
  al_nand2ft _2797_ (
    .a(_1073_),
    .b(_1074_),
    .y(_1075_)
  );
  al_ao21 _2798_ (
    .a(_1075_),
    .b(_1025_),
    .c(_1039_),
    .y(\DFF_11.D )
  );
  al_nand3ftt _2799_ (
    .a(\DFF_466.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1076_)
  );
  al_mux2h _2800_ (
    .a(\DFF_109.Q ),
    .b(_0961_),
    .s(_1076_),
    .y(\DFF_466.D )
  );
  al_or3fft _2801_ (
    .a(\DFF_48.Q ),
    .b(_0800_),
    .c(_0954_),
    .y(_1077_)
  );
  al_ao21ttf _2802_ (
    .a(\DFF_15.Q ),
    .b(_0954_),
    .c(_1077_),
    .y(\DFF_48.D )
  );
  al_and3ftt _2803_ (
    .a(\DFF_31.Q ),
    .b(\DFF_158.Q ),
    .c(_0490_),
    .y(_1078_)
  );
  al_or2ft _2804_ (
    .a(\DFF_323.Q ),
    .b(_1078_),
    .y(_1079_)
  );
  al_and2ft _2805_ (
    .a(\DFF_323.Q ),
    .b(_1078_),
    .y(_1080_)
  );
  al_nand2ft _2806_ (
    .a(_1080_),
    .b(_1079_),
    .y(_1081_)
  );
  al_nor2 _2807_ (
    .a(\DFF_525.Q ),
    .b(\DFF_366.Q ),
    .y(_1082_)
  );
  al_nand3fft _2808_ (
    .a(\DFF_240.Q ),
    .b(\DFF_353.Q ),
    .c(_1082_),
    .y(_1083_)
  );
  al_or3 _2809_ (
    .a(\DFF_399.Q ),
    .b(\DFF_214.Q ),
    .c(\DFF_468.Q ),
    .y(_1084_)
  );
  al_nor2 _2810_ (
    .a(\DFF_232.Q ),
    .b(\DFF_517.Q ),
    .y(_1085_)
  );
  al_nand3fft _2811_ (
    .a(\DFF_457.Q ),
    .b(\DFF_438.Q ),
    .c(_1085_),
    .y(_1086_)
  );
  al_and3fft _2812_ (
    .a(\DFF_145.Q ),
    .b(_1086_),
    .c(_0722_),
    .y(_1087_)
  );
  al_nand3fft _2813_ (
    .a(_1083_),
    .b(_1084_),
    .c(_1087_),
    .y(_1088_)
  );
  al_nand3fft _2814_ (
    .a(\DFF_7.Q ),
    .b(\DFF_383.Q ),
    .c(_1088_),
    .y(_1089_)
  );
  al_aoi21ttf _2815_ (
    .a(\DFF_7.Q ),
    .b(\DFF_383.Q ),
    .c(_1089_),
    .y(_1090_)
  );
  al_and2ft _2816_ (
    .a(_1081_),
    .b(_1090_),
    .y(_1091_)
  );
  al_or2ft _2817_ (
    .a(_1081_),
    .b(_1090_),
    .y(_1092_)
  );
  al_nand2ft _2818_ (
    .a(_1091_),
    .b(_1092_),
    .y(_1093_)
  );
  al_aoi21 _2819_ (
    .a(_1093_),
    .b(_0770_),
    .c(_0841_),
    .y(_1094_)
  );
  al_oai21 _2820_ (
    .a(_0770_),
    .b(_1093_),
    .c(_1094_),
    .y(_1095_)
  );
  al_aoi21ftf _2821_ (
    .a(\DFF_509.Q ),
    .b(_0841_),
    .c(_1095_),
    .y(\DFF_509.D )
  );
  al_nand3ftt _2822_ (
    .a(_0809_),
    .b(g109),
    .c(\DFF_384.D ),
    .y(_1096_)
  );
  al_ao21ttf _2823_ (
    .a(\DFF_530.Q ),
    .b(_0809_),
    .c(_1096_),
    .y(\DFF_530.D )
  );
  al_nand3ftt _2824_ (
    .a(\DFF_505.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1097_)
  );
  al_mux2h _2825_ (
    .a(\DFF_97.Q ),
    .b(_0961_),
    .s(_1097_),
    .y(\DFF_505.D )
  );
  al_oai21ftf _2826_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_213.Q ),
    .y(\DFF_213.D )
  );
  al_nand3ftt _2827_ (
    .a(\DFF_426.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1098_)
  );
  al_mux2h _2828_ (
    .a(\DFF_437.Q ),
    .b(_0961_),
    .s(_1098_),
    .y(\DFF_426.D )
  );
  al_ao21 _2829_ (
    .a(\DFF_323.Q ),
    .b(\DFF_320.Q ),
    .c(\DFF_282.Q ),
    .y(_1099_)
  );
  al_mux2h _2830_ (
    .a(\DFF_346.Q ),
    .b(_0966_),
    .s(_1099_),
    .y(\DFF_282.D )
  );
  al_and2 _2831_ (
    .a(\DFF_227.Q ),
    .b(\DFF_429.Q ),
    .y(_1100_)
  );
  al_or2 _2832_ (
    .a(\DFF_227.Q ),
    .b(\DFF_429.Q ),
    .y(_1101_)
  );
  al_oai21ftt _2833_ (
    .a(_1101_),
    .b(_1100_),
    .c(_0455_),
    .y(\DFF_429.D )
  );
  al_nand3ftt _2834_ (
    .a(\DFF_256.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1102_)
  );
  al_mux2h _2835_ (
    .a(\DFF_165.Q ),
    .b(_0961_),
    .s(_1102_),
    .y(\DFF_256.D )
  );
  al_nor3fft _2836_ (
    .a(\DFF_58.Q ),
    .b(\DFF_0.Q ),
    .c(_0443_),
    .y(_1103_)
  );
  al_ao21 _2837_ (
    .a(\DFF_322.Q ),
    .b(_0839_),
    .c(_1103_),
    .y(\DFF_322.D )
  );
  al_nand2ft _2838_ (
    .a(g85),
    .b(g92),
    .y(_1104_)
  );
  al_ao21ttf _2839_ (
    .a(g85),
    .b(\DFF_305.Q ),
    .c(_1104_),
    .y(\DFF_305.D )
  );
  al_or3 _2840_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_94.Q ),
    .y(_1105_)
  );
  al_mux2h _2841_ (
    .a(\DFF_414.Q ),
    .b(_0635_),
    .s(_1105_),
    .y(\DFF_414.D )
  );
  al_nand3ftt _2842_ (
    .a(\DFF_463.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1106_)
  );
  al_mux2h _2843_ (
    .a(\DFF_98.Q ),
    .b(_0961_),
    .s(_1106_),
    .y(\DFF_463.D )
  );
  al_nand3 _2844_ (
    .a(\DFF_394.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1107_)
  );
  al_ao21ttf _2845_ (
    .a(\DFF_217.Q ),
    .b(_0355_),
    .c(_1107_),
    .y(\DFF_394.D )
  );
  al_and3fft _2846_ (
    .a(\DFF_113.Q ),
    .b(_0720_),
    .c(_0981_),
    .y(_1108_)
  );
  al_ao21 _2847_ (
    .a(_0983_),
    .b(\DFF_242.D ),
    .c(_1108_),
    .y(_1109_)
  );
  al_nand2 _2848_ (
    .a(_0635_),
    .b(_1109_),
    .y(_1110_)
  );
  al_ao21ftf _2849_ (
    .a(_0635_),
    .b(\DFF_186.Q ),
    .c(_1110_),
    .y(\DFF_186.D )
  );
  al_nand3 _2850_ (
    .a(\DFF_215.Q ),
    .b(_0445_),
    .c(_0442_),
    .y(_1111_)
  );
  al_nand2 _2851_ (
    .a(\DFF_325.Q ),
    .b(_1111_),
    .y(_1112_)
  );
  al_ao21ftf _2852_ (
    .a(_1111_),
    .b(\DFF_75.Q ),
    .c(_1112_),
    .y(\DFF_325.D )
  );
  al_nand2ft _2853_ (
    .a(\DFF_276.Q ),
    .b(\DFF_285.Q ),
    .y(_1113_)
  );
  al_ao21ttf _2854_ (
    .a(\DFF_276.Q ),
    .b(\DFF_69.Q ),
    .c(_1113_),
    .y(g6926)
  );
  al_nor3fft _2855_ (
    .a(\DFF_0.Q ),
    .b(\DFF_250.Q ),
    .c(_0443_),
    .y(_1114_)
  );
  al_ao21 _2856_ (
    .a(\DFF_486.Q ),
    .b(_0839_),
    .c(_1114_),
    .y(\DFF_486.D )
  );
  al_ao21ftf _2857_ (
    .a(_0457_),
    .b(\DFF_111.Q ),
    .c(_0647_),
    .y(\DFF_111.D )
  );
  al_ao21 _2858_ (
    .a(\DFF_323.Q ),
    .b(\DFF_320.Q ),
    .c(\DFF_410.Q ),
    .y(_1115_)
  );
  al_mux2h _2859_ (
    .a(\DFF_324.Q ),
    .b(_0966_),
    .s(_1115_),
    .y(\DFF_410.D )
  );
  al_and2 _2860_ (
    .a(_0477_),
    .b(_0478_),
    .y(_1116_)
  );
  al_nand3fft _2861_ (
    .a(\DFF_333.Q ),
    .b(\DFF_354.Q ),
    .c(_1116_),
    .y(_1117_)
  );
  al_aoi21ttf _2862_ (
    .a(\DFF_333.Q ),
    .b(_0473_),
    .c(_1117_),
    .y(_1118_)
  );
  al_nor2ft _2863_ (
    .a(\DFF_209.Q ),
    .b(_0944_),
    .y(_1119_)
  );
  al_mux2l _2864_ (
    .a(_0945_),
    .b(_1118_),
    .s(_1119_),
    .y(_1120_)
  );
  al_and2 _2865_ (
    .a(\DFF_461.Q ),
    .b(_1120_),
    .y(_1121_)
  );
  al_or2 _2866_ (
    .a(\DFF_461.Q ),
    .b(_1120_),
    .y(_1122_)
  );
  al_nand2ft _2867_ (
    .a(_1121_),
    .b(_1122_),
    .y(_1123_)
  );
  al_ao21 _2868_ (
    .a(_1123_),
    .b(_0513_),
    .c(_0951_),
    .y(\DFF_461.D )
  );
  al_nand3 _2869_ (
    .a(\DFF_522.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1124_)
  );
  al_ao21ttf _2870_ (
    .a(\DFF_203.Q ),
    .b(_0355_),
    .c(_1124_),
    .y(\DFF_522.D )
  );
  al_nand2 _2871_ (
    .a(\DFF_458.Q ),
    .b(_1111_),
    .y(_1125_)
  );
  al_ao21ftf _2872_ (
    .a(_1111_),
    .b(\DFF_59.Q ),
    .c(_1125_),
    .y(\DFF_458.D )
  );
  al_and3 _2873_ (
    .a(\DFF_309.Q ),
    .b(_0536_),
    .c(\DFF_37.D ),
    .y(_1126_)
  );
  al_ao21 _2874_ (
    .a(\DFF_365.Q ),
    .b(_0977_),
    .c(_1126_),
    .y(\DFF_365.D )
  );
  al_nand3ftt _2875_ (
    .a(\DFF_254.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1127_)
  );
  al_mux2h _2876_ (
    .a(\DFF_24.Q ),
    .b(_0961_),
    .s(_1127_),
    .y(\DFF_254.D )
  );
  al_or3 _2877_ (
    .a(\DFF_72.Q ),
    .b(_0396_),
    .c(_0669_),
    .y(_1128_)
  );
  al_nand2 _2878_ (
    .a(\DFF_72.Q ),
    .b(_0669_),
    .y(_1129_)
  );
  al_nand3 _2879_ (
    .a(_0800_),
    .b(_1129_),
    .c(_1128_),
    .y(\DFF_72.D )
  );
  al_aoi21 _2880_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_120.Q ),
    .y(_1130_)
  );
  al_mux2l _2881_ (
    .a(_0809_),
    .b(_0539_),
    .s(_1130_),
    .y(\DFF_120.D )
  );
  al_oa21ftf _2882_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_70.Q ),
    .y(_1131_)
  );
  al_mux2l _2883_ (
    .a(_1017_),
    .b(_0901_),
    .s(_1131_),
    .y(\DFF_70.D )
  );
  al_nand3ftt _2884_ (
    .a(\DFF_39.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1132_)
  );
  al_mux2h _2885_ (
    .a(\DFF_277.Q ),
    .b(_0961_),
    .s(_1132_),
    .y(\DFF_39.D )
  );
  al_inv _2886_ (
    .a(_0958_),
    .y(_1133_)
  );
  al_nor2 _2887_ (
    .a(\DFF_241.Q ),
    .b(\DFF_113.Q ),
    .y(_1134_)
  );
  al_ao21ttf _2888_ (
    .a(g109),
    .b(\DFF_319.D ),
    .c(_1042_),
    .y(_1135_)
  );
  al_aoi21ttf _2889_ (
    .a(_0783_),
    .b(_1134_),
    .c(_1135_),
    .y(_1136_)
  );
  al_oa21ftf _2890_ (
    .a(\DFF_372.Q ),
    .b(g1696),
    .c(\DFF_285.Q ),
    .y(_1137_)
  );
  al_mux2l _2891_ (
    .a(_1133_),
    .b(_1136_),
    .s(_1137_),
    .y(\DFF_285.D )
  );
  al_nand3 _2892_ (
    .a(\DFF_203.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1138_)
  );
  al_ao21ttf _2893_ (
    .a(\DFF_205.Q ),
    .b(_0355_),
    .c(_1138_),
    .y(\DFF_203.D )
  );
  al_mux2l _2894_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .s(\DFF_161.Q ),
    .y(_1139_)
  );
  al_and2ft _2895_ (
    .a(\DFF_428.Q ),
    .b(\DFF_414.Q ),
    .y(_1140_)
  );
  al_nand2ft _2896_ (
    .a(\DFF_414.Q ),
    .b(\DFF_428.Q ),
    .y(_1141_)
  );
  al_nand2ft _2897_ (
    .a(_1140_),
    .b(_1141_),
    .y(_1142_)
  );
  al_nand2 _2898_ (
    .a(\DFF_515.Q ),
    .b(\DFF_497.Q ),
    .y(_1143_)
  );
  al_nor2 _2899_ (
    .a(\DFF_515.Q ),
    .b(\DFF_497.Q ),
    .y(_1144_)
  );
  al_and3ftt _2900_ (
    .a(_1144_),
    .b(_1143_),
    .c(_1142_),
    .y(_1145_)
  );
  al_ao21ftt _2901_ (
    .a(_1144_),
    .b(_1143_),
    .c(_1142_),
    .y(_1146_)
  );
  al_nand2ft _2902_ (
    .a(_1145_),
    .b(_1146_),
    .y(_1147_)
  );
  al_and2ft _2903_ (
    .a(\DFF_115.Q ),
    .b(\DFF_167.Q ),
    .y(_1148_)
  );
  al_nand2ft _2904_ (
    .a(\DFF_167.Q ),
    .b(\DFF_115.Q ),
    .y(_1149_)
  );
  al_nand2ft _2905_ (
    .a(_1148_),
    .b(_1149_),
    .y(_1150_)
  );
  al_and2ft _2906_ (
    .a(\DFF_108.Q ),
    .b(\DFF_192.Q ),
    .y(_1151_)
  );
  al_nand2ft _2907_ (
    .a(\DFF_192.Q ),
    .b(\DFF_108.Q ),
    .y(_1152_)
  );
  al_and2ft _2908_ (
    .a(\DFF_87.Q ),
    .b(\DFF_413.Q ),
    .y(_1153_)
  );
  al_nand2ft _2909_ (
    .a(\DFF_413.Q ),
    .b(\DFF_87.Q ),
    .y(_1154_)
  );
  al_nand2ft _2910_ (
    .a(_1153_),
    .b(_1154_),
    .y(_1155_)
  );
  al_nand3ftt _2911_ (
    .a(_1151_),
    .b(_1152_),
    .c(_1155_),
    .y(_1156_)
  );
  al_aoi21ftt _2912_ (
    .a(_1151_),
    .b(_1152_),
    .c(_1155_),
    .y(_1157_)
  );
  al_nor3fft _2913_ (
    .a(_1150_),
    .b(_1156_),
    .c(_1157_),
    .y(_1158_)
  );
  al_oai21ftf _2914_ (
    .a(_1156_),
    .b(_1157_),
    .c(_1150_),
    .y(_1159_)
  );
  al_aoi21ftt _2915_ (
    .a(_1158_),
    .b(_1159_),
    .c(_1147_),
    .y(_1160_)
  );
  al_and3ftt _2916_ (
    .a(_1158_),
    .b(_1147_),
    .c(_1159_),
    .y(_1161_)
  );
  al_mux2h _2917_ (
    .a(_1161_),
    .b(_1160_),
    .s(_0635_),
    .y(_1162_)
  );
  al_aoi21 _2918_ (
    .a(_1162_),
    .b(_0399_),
    .c(_1139_),
    .y(\DFF_161.D )
  );
  al_nand3ftt _2919_ (
    .a(\DFF_81.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1163_)
  );
  al_mux2h _2920_ (
    .a(\DFF_36.Q ),
    .b(_0961_),
    .s(_1163_),
    .y(\DFF_81.D )
  );
  al_mux2l _2921_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .s(\DFF_166.Q ),
    .y(_1164_)
  );
  al_mux2l _2922_ (
    .a(_0841_),
    .b(_1136_),
    .s(_1164_),
    .y(\DFF_166.D )
  );
  al_nor3fft _2923_ (
    .a(\DFF_498.Q ),
    .b(\DFF_0.Q ),
    .c(_0443_),
    .y(_1165_)
  );
  al_ao21 _2924_ (
    .a(\DFF_61.Q ),
    .b(_0839_),
    .c(_1165_),
    .y(\DFF_61.D )
  );
  al_ao21ttf _2925_ (
    .a(g109),
    .b(\DFF_384.D ),
    .c(_1042_),
    .y(_1166_)
  );
  al_aoi21ttf _2926_ (
    .a(_0713_),
    .b(_1134_),
    .c(_1166_),
    .y(_1167_)
  );
  al_oa21ftf _2927_ (
    .a(\DFF_372.Q ),
    .b(g1696),
    .c(\DFF_280.Q ),
    .y(_1168_)
  );
  al_mux2l _2928_ (
    .a(_1133_),
    .b(_1167_),
    .s(_1168_),
    .y(\DFF_280.D )
  );
  al_nand3ftt _2929_ (
    .a(\DFF_477.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1169_)
  );
  al_mux2h _2930_ (
    .a(\DFF_143.Q ),
    .b(_0961_),
    .s(_1169_),
    .y(\DFF_477.D )
  );
  al_nand3ftt _2931_ (
    .a(\DFF_164.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1170_)
  );
  al_mux2h _2932_ (
    .a(\DFF_34.Q ),
    .b(_0961_),
    .s(_1170_),
    .y(\DFF_164.D )
  );
  al_inv _2933_ (
    .a(\DFF_180.Q ),
    .y(_1171_)
  );
  al_mux2h _2934_ (
    .a(_1171_),
    .b(_0954_),
    .s(_0800_),
    .y(_1172_)
  );
  al_ao21ftf _2935_ (
    .a(_0760_),
    .b(_0954_),
    .c(_1172_),
    .y(\DFF_180.D )
  );
  al_ao21ftf _2936_ (
    .a(_0635_),
    .b(\DFF_465.Q ),
    .c(_1046_),
    .y(\DFF_465.D )
  );
  al_and2 _2937_ (
    .a(_1134_),
    .b(_0729_),
    .y(_1173_)
  );
  al_oa21ftf _2938_ (
    .a(_0983_),
    .b(\DFF_168.D ),
    .c(_1173_),
    .y(_1174_)
  );
  al_oa21ftf _2939_ (
    .a(\DFF_372.Q ),
    .b(g1696),
    .c(\DFF_45.Q ),
    .y(_1175_)
  );
  al_mux2l _2940_ (
    .a(_1133_),
    .b(_1174_),
    .s(_1175_),
    .y(\DFF_45.D )
  );
  al_nor3fft _2941_ (
    .a(\DFF_334.Q ),
    .b(\DFF_0.Q ),
    .c(_0443_),
    .y(_1176_)
  );
  al_ao21 _2942_ (
    .a(\DFF_231.Q ),
    .b(_0839_),
    .c(_1176_),
    .y(\DFF_231.D )
  );
  al_or3fft _2943_ (
    .a(_0981_),
    .b(_1044_),
    .c(_0751_),
    .y(_1177_)
  );
  al_mux2h _2944_ (
    .a(_0225_),
    .b(_0284_),
    .s(_0983_),
    .y(_1178_)
  );
  al_oai21ftf _2945_ (
    .a(_1177_),
    .b(_1178_),
    .c(_0841_),
    .y(_1179_)
  );
  al_ao21ftf _2946_ (
    .a(_0635_),
    .b(\DFF_26.Q ),
    .c(_1179_),
    .y(\DFF_26.D )
  );
  al_nand3 _2947_ (
    .a(\DFF_214.Q ),
    .b(_0803_),
    .c(_0490_),
    .y(_1180_)
  );
  al_ao21 _2948_ (
    .a(_0803_),
    .b(_0490_),
    .c(\DFF_214.Q ),
    .y(_1181_)
  );
  al_ao21 _2949_ (
    .a(_1180_),
    .b(_1181_),
    .c(_0841_),
    .y(_1182_)
  );
  al_aoi21ftf _2950_ (
    .a(\DFF_74.Q ),
    .b(_0841_),
    .c(_1182_),
    .y(\DFF_74.D )
  );
  al_or3 _2951_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_292.Q ),
    .y(_1183_)
  );
  al_mux2h _2952_ (
    .a(\DFF_192.Q ),
    .b(_0635_),
    .s(_1183_),
    .y(\DFF_192.D )
  );
  al_nand2ft _2953_ (
    .a(\DFF_276.Q ),
    .b(\DFF_45.Q ),
    .y(_1184_)
  );
  al_ao21ttf _2954_ (
    .a(\DFF_276.Q ),
    .b(\DFF_101.Q ),
    .c(_1184_),
    .y(g6932)
  );
  al_or3 _2955_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_290.Q ),
    .y(_1185_)
  );
  al_mux2h _2956_ (
    .a(\DFF_428.Q ),
    .b(_0635_),
    .s(_1185_),
    .y(\DFF_428.D )
  );
  al_oai21ttf _2957_ (
    .a(_0479_),
    .b(_0473_),
    .c(_0945_),
    .y(_1186_)
  );
  al_aoi21ftf _2958_ (
    .a(_0944_),
    .b(\DFF_493.Q ),
    .c(_1186_),
    .y(_1187_)
  );
  al_and2 _2959_ (
    .a(\DFF_333.Q ),
    .b(_1187_),
    .y(_1188_)
  );
  al_or2 _2960_ (
    .a(\DFF_333.Q ),
    .b(_1187_),
    .y(_1189_)
  );
  al_nand2ft _2961_ (
    .a(_1188_),
    .b(_1189_),
    .y(_1190_)
  );
  al_ao21 _2962_ (
    .a(_1190_),
    .b(_0513_),
    .c(_0951_),
    .y(\DFF_333.D )
  );
  al_oa21ftt _2963_ (
    .a(\DFF_372.Q ),
    .b(g1696),
    .c(\DFF_292.Q ),
    .y(_1191_)
  );
  al_ao21 _2964_ (
    .a(\DFF_499.Q ),
    .b(_0958_),
    .c(_1191_),
    .y(\DFF_292.D )
  );
  al_nand3 _2965_ (
    .a(_0006_),
    .b(_0876_),
    .c(_0881_),
    .y(_1192_)
  );
  al_aoi21ftf _2966_ (
    .a(\DFF_79.Q ),
    .b(_1017_),
    .c(_1192_),
    .y(\DFF_79.D )
  );
  al_nand2ft _2967_ (
    .a(g85),
    .b(g91),
    .y(_1193_)
  );
  al_ao21ttf _2968_ (
    .a(g85),
    .b(\DFF_110.Q ),
    .c(_1193_),
    .y(\DFF_110.D )
  );
  al_oa21ftt _2969_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_263.Q ),
    .y(_1194_)
  );
  al_nand3 _2970_ (
    .a(_0399_),
    .b(_0918_),
    .c(_0921_),
    .y(_1195_)
  );
  al_mux2l _2971_ (
    .a(_0399_),
    .b(_0936_),
    .s(_1017_),
    .y(_1196_)
  );
  al_ao21 _2972_ (
    .a(_1196_),
    .b(_1195_),
    .c(_1194_),
    .y(\DFF_263.D )
  );
  al_or3 _2973_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_471.Q ),
    .y(_1197_)
  );
  al_mux2h _2974_ (
    .a(\DFF_174.Q ),
    .b(_0635_),
    .s(_1197_),
    .y(\DFF_174.D )
  );
  al_nand3 _2975_ (
    .a(\DFF_151.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1198_)
  );
  al_ao21ttf _2976_ (
    .a(\DFF_430.Q ),
    .b(_0355_),
    .c(_1198_),
    .y(\DFF_151.D )
  );
  al_nor3fft _2977_ (
    .a(\DFF_486.Q ),
    .b(\DFF_0.Q ),
    .c(_0443_),
    .y(_1199_)
  );
  al_ao21 _2978_ (
    .a(\DFF_401.Q ),
    .b(_0839_),
    .c(_1199_),
    .y(\DFF_401.D )
  );
  al_nand3ftt _2979_ (
    .a(\DFF_326.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1200_)
  );
  al_mux2h _2980_ (
    .a(\DFF_95.Q ),
    .b(_0961_),
    .s(_1200_),
    .y(\DFF_326.D )
  );
  al_or3fft _2981_ (
    .a(\DFF_209.Q ),
    .b(_0512_),
    .c(_1012_),
    .y(_1201_)
  );
  al_ao21ttf _2982_ (
    .a(\DFF_493.Q ),
    .b(_1012_),
    .c(_1201_),
    .y(\DFF_209.D )
  );
  al_nand2ft _2983_ (
    .a(g85),
    .b(g93),
    .y(_1202_)
  );
  al_ao21ttf _2984_ (
    .a(g85),
    .b(\DFF_348.Q ),
    .c(_1202_),
    .y(\DFF_348.D )
  );
  al_nand3ftt _2985_ (
    .a(\DFF_259.Q ),
    .b(g109),
    .c(_0589_),
    .y(_1203_)
  );
  al_mux2h _2986_ (
    .a(\DFF_508.Q ),
    .b(_0956_),
    .s(_1203_),
    .y(\DFF_259.D )
  );
  al_ao21ttf _2987_ (
    .a(_0607_),
    .b(_0605_),
    .c(\DFF_532.Q ),
    .y(_1204_)
  );
  al_nand3 _2988_ (
    .a(_0512_),
    .b(_0672_),
    .c(_1204_),
    .y(\DFF_532.D )
  );
  al_oai21ftt _2989_ (
    .a(_1134_),
    .b(_0747_),
    .c(_0635_),
    .y(_1205_)
  );
  al_oai21ftf _2990_ (
    .a(_0983_),
    .b(\DFF_384.D ),
    .c(_1205_),
    .y(_1206_)
  );
  al_ao21ftf _2991_ (
    .a(_0635_),
    .b(\DFF_69.Q ),
    .c(_1206_),
    .y(\DFF_69.D )
  );
  al_aoi21ftf _2992_ (
    .a(_1028_),
    .b(_1171_),
    .c(_1069_),
    .y(_1207_)
  );
  al_and2ft _2993_ (
    .a(\DFF_395.Q ),
    .b(_1207_),
    .y(_1208_)
  );
  al_or2ft _2994_ (
    .a(\DFF_395.Q ),
    .b(_1207_),
    .y(_1209_)
  );
  al_nand2ft _2995_ (
    .a(_1208_),
    .b(_1209_),
    .y(_1210_)
  );
  al_ao21 _2996_ (
    .a(_1210_),
    .b(_1025_),
    .c(_1039_),
    .y(\DFF_395.D )
  );
  al_and3 _2997_ (
    .a(\DFF_405.Q ),
    .b(_0536_),
    .c(\DFF_37.D ),
    .y(_1211_)
  );
  al_ao21 _2998_ (
    .a(\DFF_148.Q ),
    .b(_0977_),
    .c(_1211_),
    .y(\DFF_148.D )
  );
  al_nand3ftt _2999_ (
    .a(\DFF_20.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1212_)
  );
  al_mux2h _3000_ (
    .a(\DFF_169.Q ),
    .b(_0961_),
    .s(_1212_),
    .y(\DFF_20.D )
  );
  al_mux2l _3001_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .s(\DFF_159.Q ),
    .y(_1213_)
  );
  al_mux2l _3002_ (
    .a(_0841_),
    .b(_1167_),
    .s(_1213_),
    .y(\DFF_159.D )
  );
  al_nand2 _3003_ (
    .a(\DFF_481.Q ),
    .b(_1111_),
    .y(_1214_)
  );
  al_ao21ftf _3004_ (
    .a(_1111_),
    .b(\DFF_268.Q ),
    .c(_1214_),
    .y(\DFF_481.D )
  );
  al_or2 _3005_ (
    .a(\DFF_191.Q ),
    .b(\DFF_262.D ),
    .y(\DFF_336.D )
  );
  al_nand3ftt _3006_ (
    .a(\DFF_453.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1215_)
  );
  al_mux2h _3007_ (
    .a(\DFF_172.Q ),
    .b(_0961_),
    .s(_1215_),
    .y(\DFF_453.D )
  );
  al_nand3ftt _3008_ (
    .a(_0809_),
    .b(g109),
    .c(\DFF_228.D ),
    .y(_1216_)
  );
  al_ao21ttf _3009_ (
    .a(\DFF_96.Q ),
    .b(_0809_),
    .c(_1216_),
    .y(\DFF_96.D )
  );
  al_nor3fft _3010_ (
    .a(\DFF_202.Q ),
    .b(\DFF_0.Q ),
    .c(_0443_),
    .y(_1217_)
  );
  al_ao21 _3011_ (
    .a(\DFF_334.Q ),
    .b(_0839_),
    .c(_1217_),
    .y(\DFF_334.D )
  );
  al_nand3ftt _3012_ (
    .a(\DFF_258.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1218_)
  );
  al_mux2h _3013_ (
    .a(\DFF_273.Q ),
    .b(_0961_),
    .s(_1218_),
    .y(\DFF_258.D )
  );
  al_oa21ftt _3014_ (
    .a(\DFF_372.Q ),
    .b(g1696),
    .c(\DFF_170.Q ),
    .y(_1219_)
  );
  al_ao21 _3015_ (
    .a(\DFF_230.Q ),
    .b(_0958_),
    .c(_1219_),
    .y(\DFF_170.D )
  );
  al_or3fft _3016_ (
    .a(\DFF_85.Q ),
    .b(_0512_),
    .c(_1012_),
    .y(_1220_)
  );
  al_ao21ttf _3017_ (
    .a(\DFF_349.Q ),
    .b(_1012_),
    .c(_1220_),
    .y(\DFF_85.D )
  );
  al_oai21ftf _3018_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_533.Q ),
    .y(\DFF_533.D )
  );
  al_and3 _3019_ (
    .a(\DFF_55.Q ),
    .b(_0536_),
    .c(\DFF_37.D ),
    .y(_1221_)
  );
  al_ao21 _3020_ (
    .a(\DFF_312.Q ),
    .b(_0977_),
    .c(_1221_),
    .y(\DFF_312.D )
  );
  al_ao21ftf _3021_ (
    .a(_0635_),
    .b(\DFF_73.Q ),
    .c(_1049_),
    .y(\DFF_73.D )
  );
  al_nand3ftt _3022_ (
    .a(\DFF_514.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1222_)
  );
  al_mux2h _3023_ (
    .a(\DFF_139.Q ),
    .b(_0961_),
    .s(_1222_),
    .y(\DFF_514.D )
  );
  al_nand3 _3024_ (
    .a(_0635_),
    .b(_0651_),
    .c(_0757_),
    .y(_1223_)
  );
  al_aoi21ftf _3025_ (
    .a(\DFF_495.Q ),
    .b(_0841_),
    .c(_1223_),
    .y(\DFF_495.D )
  );
  al_nand2ft _3026_ (
    .a(g85),
    .b(g89),
    .y(_1224_)
  );
  al_ao21ttf _3027_ (
    .a(g85),
    .b(\DFF_236.Q ),
    .c(_1224_),
    .y(\DFF_236.D )
  );
  al_nand3 _3028_ (
    .a(\DFF_512.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1225_)
  );
  al_ao21ttf _3029_ (
    .a(\DFF_378.Q ),
    .b(_0355_),
    .c(_1225_),
    .y(\DFF_512.D )
  );
  al_nand3ftt _3030_ (
    .a(\DFF_391.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1226_)
  );
  al_mux2h _3031_ (
    .a(\DFF_201.Q ),
    .b(_0961_),
    .s(_1226_),
    .y(\DFF_391.D )
  );
  al_nand3ftt _3032_ (
    .a(\DFF_279.Q ),
    .b(g109),
    .c(_0589_),
    .y(_1227_)
  );
  al_mux2h _3033_ (
    .a(\DFF_382.Q ),
    .b(_0956_),
    .s(_1227_),
    .y(\DFF_279.D )
  );
  al_nand3 _3034_ (
    .a(_0635_),
    .b(_0521_),
    .c(_0525_),
    .y(_1228_)
  );
  al_aoi21ftf _3035_ (
    .a(\DFF_199.Q ),
    .b(_0841_),
    .c(_1228_),
    .y(\DFF_199.D )
  );
  al_nand2ft _3036_ (
    .a(g85),
    .b(g94),
    .y(_1229_)
  );
  al_ao21ttf _3037_ (
    .a(g85),
    .b(\DFF_298.Q ),
    .c(_1229_),
    .y(\DFF_298.D )
  );
  al_nor3fft _3038_ (
    .a(\DFF_32.Q ),
    .b(\DFF_0.Q ),
    .c(_0443_),
    .y(_1230_)
  );
  al_ao21 _3039_ (
    .a(\DFF_498.Q ),
    .b(_0839_),
    .c(_1230_),
    .y(\DFF_498.D )
  );
  al_nand3 _3040_ (
    .a(\DFF_447.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1231_)
  );
  al_ao21ttf _3041_ (
    .a(\DFF_475.Q ),
    .b(_0355_),
    .c(_1231_),
    .y(\DFF_447.D )
  );
  al_nand3ftt _3042_ (
    .a(_0809_),
    .b(g109),
    .c(\DFF_242.D ),
    .y(_1232_)
  );
  al_ao21ttf _3043_ (
    .a(\DFF_370.Q ),
    .b(_0809_),
    .c(_1232_),
    .y(\DFF_370.D )
  );
  al_nand3 _3044_ (
    .a(\DFF_171.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1233_)
  );
  al_ao21ttf _3045_ (
    .a(\DFF_368.Q ),
    .b(_0355_),
    .c(_1233_),
    .y(\DFF_171.D )
  );
  al_oa21ftt _3046_ (
    .a(\DFF_372.Q ),
    .b(g1696),
    .c(\DFF_27.Q ),
    .y(_1234_)
  );
  al_ao21 _3047_ (
    .a(\DFF_266.Q ),
    .b(_0958_),
    .c(_1234_),
    .y(\DFF_27.D )
  );
  al_nand3 _3048_ (
    .a(\DFF_368.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1235_)
  );
  al_ao21ttf _3049_ (
    .a(\DFF_3.Q ),
    .b(_0355_),
    .c(_1235_),
    .y(\DFF_368.D )
  );
  al_oa21ftt _3050_ (
    .a(\DFF_372.Q ),
    .b(g1696),
    .c(\DFF_376.Q ),
    .y(_1236_)
  );
  al_ao21 _3051_ (
    .a(\DFF_263.Q ),
    .b(_0958_),
    .c(_1236_),
    .y(\DFF_376.D )
  );
  al_nand2 _3052_ (
    .a(\DFF_134.Q ),
    .b(_1111_),
    .y(_1237_)
  );
  al_ao21ftf _3053_ (
    .a(_1111_),
    .b(\DFF_103.Q ),
    .c(_1237_),
    .y(\DFF_134.D )
  );
  al_nand3 _3054_ (
    .a(\DFF_245.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1238_)
  );
  al_ao21ttf _3055_ (
    .a(\DFF_529.Q ),
    .b(_0355_),
    .c(_1238_),
    .y(\DFF_245.D )
  );
  al_or2 _3056_ (
    .a(\DFF_15.Q ),
    .b(_1028_),
    .y(_1239_)
  );
  al_and2 _3057_ (
    .a(_0694_),
    .b(_0696_),
    .y(_1240_)
  );
  al_nand3fft _3058_ (
    .a(\DFF_316.Q ),
    .b(\DFF_11.Q ),
    .c(_1240_),
    .y(_1241_)
  );
  al_or3fft _3059_ (
    .a(_1028_),
    .b(_1241_),
    .c(_1026_),
    .y(_1242_)
  );
  al_and3 _3060_ (
    .a(_1069_),
    .b(_1239_),
    .c(_1242_),
    .y(_1243_)
  );
  al_and2 _3061_ (
    .a(_0692_),
    .b(_1243_),
    .y(_1244_)
  );
  al_or2 _3062_ (
    .a(_0692_),
    .b(_1243_),
    .y(_1245_)
  );
  al_nand2ft _3063_ (
    .a(_1244_),
    .b(_1245_),
    .y(_1246_)
  );
  al_ao21 _3064_ (
    .a(_1025_),
    .b(_1246_),
    .c(_1039_),
    .y(\DFF_57.D )
  );
  al_or3fft _3065_ (
    .a(\DFF_339.Q ),
    .b(_0512_),
    .c(_1012_),
    .y(_1247_)
  );
  al_ao21ttf _3066_ (
    .a(\DFF_209.Q ),
    .b(_1012_),
    .c(_1247_),
    .y(\DFF_339.D )
  );
  al_ao21ftf _3067_ (
    .a(_0635_),
    .b(\DFF_460.Q ),
    .c(_1179_),
    .y(\DFF_460.D )
  );
  al_nand3 _3068_ (
    .a(\DFF_529.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1248_)
  );
  al_ao21ttf _3069_ (
    .a(\DFF_459.Q ),
    .b(_0355_),
    .c(_1248_),
    .y(\DFF_529.D )
  );
  al_aoi21ftf _3070_ (
    .a(_1028_),
    .b(_0760_),
    .c(_1069_),
    .y(_1249_)
  );
  al_nand2 _3071_ (
    .a(_1028_),
    .b(_0688_),
    .y(_1250_)
  );
  al_mux2h _3072_ (
    .a(_0699_),
    .b(_1250_),
    .s(_1249_),
    .y(_1251_)
  );
  al_or2 _3073_ (
    .a(\DFF_359.Q ),
    .b(_1251_),
    .y(_1252_)
  );
  al_aoi21ftf _3074_ (
    .a(_0678_),
    .b(_1251_),
    .c(_1025_),
    .y(_1253_)
  );
  al_ao21 _3075_ (
    .a(_1252_),
    .b(_1253_),
    .c(_1039_),
    .y(\DFF_359.D )
  );
  al_nand2ft _3076_ (
    .a(g85),
    .b(g88),
    .y(_1254_)
  );
  al_ao21ttf _3077_ (
    .a(g85),
    .b(\DFF_527.Q ),
    .c(_1254_),
    .y(\DFF_527.D )
  );
  al_nor3fft _3078_ (
    .a(\DFF_61.Q ),
    .b(\DFF_0.Q ),
    .c(_0443_),
    .y(_1255_)
  );
  al_ao21 _3079_ (
    .a(\DFF_250.Q ),
    .b(_0839_),
    .c(_1255_),
    .y(\DFF_250.D )
  );
  al_mux2l _3080_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .s(\DFF_211.Q ),
    .y(_1256_)
  );
  al_mux2l _3081_ (
    .a(_0841_),
    .b(_1174_),
    .s(_1256_),
    .y(\DFF_211.D )
  );
  al_and3 _3082_ (
    .a(\DFF_343.Q ),
    .b(_0536_),
    .c(\DFF_37.D ),
    .y(_1257_)
  );
  al_ao21 _3083_ (
    .a(\DFF_106.Q ),
    .b(_0977_),
    .c(_1257_),
    .y(\DFF_106.D )
  );
  al_oa21ftf _3084_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_420.Q ),
    .y(_1258_)
  );
  al_and3ftt _3085_ (
    .a(\DFF_372.Q ),
    .b(g1696),
    .c(_0398_),
    .y(_1259_)
  );
  al_or3ftt _3086_ (
    .a(_1259_),
    .b(\DFF_242.D ),
    .c(_0302_),
    .y(_1260_)
  );
  al_nand3fft _3087_ (
    .a(_0151_),
    .b(\DFF_350.D ),
    .c(\DFF_228.D ),
    .y(_1261_)
  );
  al_mux2l _3088_ (
    .a(_1261_),
    .b(_1260_),
    .s(_1258_),
    .y(\DFF_420.D )
  );
  al_nand3ftt _3089_ (
    .a(\DFF_371.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1262_)
  );
  al_mux2h _3090_ (
    .a(\DFF_415.Q ),
    .b(_0961_),
    .s(_1262_),
    .y(\DFF_371.D )
  );
  al_nand3ftt _3091_ (
    .a(\DFF_386.Q ),
    .b(g109),
    .c(_0589_),
    .y(_1263_)
  );
  al_mux2h _3092_ (
    .a(\DFF_364.Q ),
    .b(_0956_),
    .s(_1263_),
    .y(\DFF_386.D )
  );
  al_ao21ftf _3093_ (
    .a(_1028_),
    .b(_1007_),
    .c(_1069_),
    .y(_1264_)
  );
  al_aoi21ttf _3094_ (
    .a(\DFF_450.Q ),
    .b(_0685_),
    .c(_1028_),
    .y(_1265_)
  );
  al_aoi21ftt _3095_ (
    .a(_1240_),
    .b(_1265_),
    .c(_1264_),
    .y(_1266_)
  );
  al_and2 _3096_ (
    .a(\DFF_316.Q ),
    .b(_1266_),
    .y(_1267_)
  );
  al_or2 _3097_ (
    .a(\DFF_316.Q ),
    .b(_1266_),
    .y(_1268_)
  );
  al_and2ft _3098_ (
    .a(_1267_),
    .b(_1268_),
    .y(_1269_)
  );
  al_ao21 _3099_ (
    .a(_1269_),
    .b(_1025_),
    .c(_1039_),
    .y(\DFF_316.D )
  );
  al_nand3 _3100_ (
    .a(\DFF_378.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1270_)
  );
  al_ao21ttf _3101_ (
    .a(\DFF_171.Q ),
    .b(_0355_),
    .c(_1270_),
    .y(\DFF_378.D )
  );
  al_oa21ftf _3102_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_230.Q ),
    .y(_1271_)
  );
  al_mux2l _3103_ (
    .a(_1017_),
    .b(_0850_),
    .s(_1271_),
    .y(\DFF_230.D )
  );
  al_or2 _3104_ (
    .a(\DFF_299.Q ),
    .b(\DFF_0.Q ),
    .y(\DFF_0.D )
  );
  al_inv _3105_ (
    .a(\DFF_313.Q ),
    .y(_1272_)
  );
  al_or3fft _3106_ (
    .a(\DFF_155.Q ),
    .b(_0512_),
    .c(_1012_),
    .y(_1273_)
  );
  al_ao21ftf _3107_ (
    .a(_1272_),
    .b(_1012_),
    .c(_1273_),
    .y(\DFF_155.D )
  );
  al_or2 _3108_ (
    .a(\DFF_352.Q ),
    .b(\DFF_122.D ),
    .y(\DFF_385.D )
  );
  al_nand2 _3109_ (
    .a(\DFF_146.Q ),
    .b(_1111_),
    .y(_1274_)
  );
  al_ao21ftf _3110_ (
    .a(_1111_),
    .b(\DFF_346.Q ),
    .c(_1274_),
    .y(\DFF_146.D )
  );
  al_nand3 _3111_ (
    .a(\DFF_406.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1275_)
  );
  al_ao21ttf _3112_ (
    .a(\DFF_204.Q ),
    .b(_0355_),
    .c(_1275_),
    .y(\DFF_406.D )
  );
  al_nand2ft _3113_ (
    .a(g85),
    .b(g95),
    .y(_1276_)
  );
  al_ao21ttf _3114_ (
    .a(g85),
    .b(\DFF_160.Q ),
    .c(_1276_),
    .y(\DFF_160.D )
  );
  al_oa21ftt _3115_ (
    .a(\DFF_372.Q ),
    .b(g1696),
    .c(\DFF_173.Q ),
    .y(_1277_)
  );
  al_ao21 _3116_ (
    .a(\DFF_440.Q ),
    .b(_0958_),
    .c(_1277_),
    .y(\DFF_173.D )
  );
  al_nand3 _3117_ (
    .a(\DFF_419.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1278_)
  );
  al_ao21ttf _3118_ (
    .a(\DFF_177.Q ),
    .b(_0355_),
    .c(_1278_),
    .y(\DFF_419.D )
  );
  al_aoi21 _3119_ (
    .a(\DFF_75.Q ),
    .b(\DFF_59.Q ),
    .c(\DFF_276.Q ),
    .y(_1279_)
  );
  al_oai21ftf _3120_ (
    .a(\DFF_276.Q ),
    .b(_0306_),
    .c(_1279_),
    .y(_1280_)
  );
  al_and3ftt _3121_ (
    .a(\DFF_276.Q ),
    .b(\DFF_324.Q ),
    .c(\DFF_104.Q ),
    .y(_1281_)
  );
  al_ao21 _3122_ (
    .a(\DFF_276.Q ),
    .b(_0310_),
    .c(_1281_),
    .y(_1282_)
  );
  al_aoi21 _3123_ (
    .a(\DFF_242.D ),
    .b(\DFF_228.D ),
    .c(_1055_),
    .y(_1283_)
  );
  al_and3fft _3124_ (
    .a(\DFF_276.Q ),
    .b(_0002_),
    .c(_0597_),
    .y(_1284_)
  );
  al_aoi21 _3125_ (
    .a(_0285_),
    .b(_1283_),
    .c(_1284_),
    .y(_1285_)
  );
  al_ao21ftf _3126_ (
    .a(_1282_),
    .b(_1280_),
    .c(_1285_),
    .y(_1286_)
  );
  al_ao21ftt _3127_ (
    .a(\DFF_178.Q ),
    .b(_0017_),
    .c(_0647_),
    .y(_1287_)
  );
  al_ao21ftf _3128_ (
    .a(_0673_),
    .b(_1058_),
    .c(_1287_),
    .y(_1288_)
  );
  al_ao21ftf _3129_ (
    .a(_0512_),
    .b(_1286_),
    .c(_1288_),
    .y(\DFF_178.D )
  );
  al_nand2ft _3130_ (
    .a(g85),
    .b(g87),
    .y(_1289_)
  );
  al_ao21ttf _3131_ (
    .a(g85),
    .b(\DFF_422.Q ),
    .c(_1289_),
    .y(\DFF_422.D )
  );
  al_mux2h _3132_ (
    .a(\DFF_113.Q ),
    .b(_0635_),
    .s(_0443_),
    .y(\DFF_113.D )
  );
  al_nand2ft _3133_ (
    .a(g85),
    .b(g96),
    .y(_1290_)
  );
  al_ao21ttf _3134_ (
    .a(g85),
    .b(\DFF_35.Q ),
    .c(_1290_),
    .y(\DFF_35.D )
  );
  al_nand3 _3135_ (
    .a(_0635_),
    .b(_0488_),
    .c(_0494_),
    .y(_1291_)
  );
  al_aoi21ftf _3136_ (
    .a(\DFF_482.Q ),
    .b(_0841_),
    .c(_1291_),
    .y(\DFF_482.D )
  );
  al_nand3 _3137_ (
    .a(\DFF_177.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1292_)
  );
  al_ao21ttf _3138_ (
    .a(\DFF_114.Q ),
    .b(_0355_),
    .c(_1292_),
    .y(\DFF_177.D )
  );
  al_ao21 _3139_ (
    .a(g109),
    .b(\DFF_242.D ),
    .c(\DFF_113.Q ),
    .y(_1293_)
  );
  al_nand3fft _3140_ (
    .a(_1133_),
    .b(_1134_),
    .c(_1293_),
    .y(_1294_)
  );
  al_ao21ftf _3141_ (
    .a(_0958_),
    .b(\DFF_504.Q ),
    .c(_1294_),
    .y(\DFF_504.D )
  );
  al_or3fft _3142_ (
    .a(\DFF_60.Q ),
    .b(_0800_),
    .c(_0954_),
    .y(_1295_)
  );
  al_ao21ttf _3143_ (
    .a(\DFF_488.Q ),
    .b(_0954_),
    .c(_1295_),
    .y(\DFF_60.D )
  );
  al_or3fft _3144_ (
    .a(\DFF_349.Q ),
    .b(_0512_),
    .c(_1012_),
    .y(_1296_)
  );
  al_ao21ttf _3145_ (
    .a(\DFF_532.Q ),
    .b(_1012_),
    .c(_1296_),
    .y(\DFF_349.D )
  );
  al_nand3ftt _3146_ (
    .a(\DFF_345.Q ),
    .b(g109),
    .c(_0589_),
    .y(_1297_)
  );
  al_mux2h _3147_ (
    .a(\DFF_147.Q ),
    .b(_0956_),
    .s(_1297_),
    .y(\DFF_345.D )
  );
  al_and3 _3148_ (
    .a(\DFF_412.Q ),
    .b(_0536_),
    .c(\DFF_37.D ),
    .y(_1298_)
  );
  al_ao21 _3149_ (
    .a(\DFF_317.Q ),
    .b(_0977_),
    .c(_1298_),
    .y(\DFF_317.D )
  );
  al_nand3ftt _3150_ (
    .a(\DFF_10.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1299_)
  );
  al_mux2h _3151_ (
    .a(\DFF_306.Q ),
    .b(_0961_),
    .s(_1299_),
    .y(\DFF_10.D )
  );
  al_oa21ftt _3152_ (
    .a(\DFF_372.Q ),
    .b(g1696),
    .c(\DFF_56.Q ),
    .y(_1300_)
  );
  al_ao21 _3153_ (
    .a(\DFF_238.Q ),
    .b(_0958_),
    .c(_1300_),
    .y(\DFF_56.D )
  );
  al_oa21ftf _3154_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_283.Q ),
    .y(_1301_)
  );
  al_mux2l _3155_ (
    .a(_1017_),
    .b(_0869_),
    .s(_1301_),
    .y(\DFF_283.D )
  );
  al_ao21ftf _3156_ (
    .a(_0635_),
    .b(\DFF_260.Q ),
    .c(_0985_),
    .y(\DFF_260.D )
  );
  al_nand2ft _3157_ (
    .a(\DFF_276.Q ),
    .b(\DFF_504.Q ),
    .y(_1302_)
  );
  al_ao21ttf _3158_ (
    .a(\DFF_276.Q ),
    .b(\DFF_73.Q ),
    .c(_1302_),
    .y(g6949)
  );
  al_or3 _3159_ (
    .a(_0151_),
    .b(_0809_),
    .c(\DFF_350.D ),
    .y(_1303_)
  );
  al_aoi21ftf _3160_ (
    .a(\DFF_321.Q ),
    .b(_0809_),
    .c(_1303_),
    .y(\DFF_321.D )
  );
  al_inv _3161_ (
    .a(\DFF_85.Q ),
    .y(_1304_)
  );
  al_or3fft _3162_ (
    .a(\DFF_493.Q ),
    .b(_0512_),
    .c(_1012_),
    .y(_1305_)
  );
  al_ao21ftf _3163_ (
    .a(_1304_),
    .b(_1012_),
    .c(_1305_),
    .y(\DFF_493.D )
  );
  al_or2 _3164_ (
    .a(\DFF_48.Q ),
    .b(_1028_),
    .y(_1306_)
  );
  al_or3ftt _3165_ (
    .a(_1028_),
    .b(_0687_),
    .c(_0698_),
    .y(_1307_)
  );
  al_and3 _3166_ (
    .a(_1069_),
    .b(_1306_),
    .c(_1307_),
    .y(_1308_)
  );
  al_and2 _3167_ (
    .a(_0679_),
    .b(_1308_),
    .y(_1309_)
  );
  al_or2 _3168_ (
    .a(_0679_),
    .b(_1308_),
    .y(_1310_)
  );
  al_nand2ft _3169_ (
    .a(_1309_),
    .b(_1310_),
    .y(_1311_)
  );
  al_ao21 _3170_ (
    .a(_1025_),
    .b(_1311_),
    .c(_1039_),
    .y(\DFF_6.D )
  );
  al_ao21ftf _3171_ (
    .a(_0635_),
    .b(\DFF_101.Q ),
    .c(_1110_),
    .y(\DFF_101.D )
  );
  al_nand3 _3172_ (
    .a(\DFF_51.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1312_)
  );
  al_ao21ttf _3173_ (
    .a(\DFF_329.Q ),
    .b(_0355_),
    .c(_1312_),
    .y(\DFF_51.D )
  );
  al_oa21ftt _3174_ (
    .a(\DFF_372.Q ),
    .b(g1696),
    .c(\DFF_290.Q ),
    .y(_1313_)
  );
  al_ao21 _3175_ (
    .a(\DFF_216.Q ),
    .b(_0958_),
    .c(_1313_),
    .y(\DFF_290.D )
  );
  al_nand3ftt _3176_ (
    .a(\DFF_392.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1314_)
  );
  al_mux2h _3177_ (
    .a(\DFF_90.Q ),
    .b(_0961_),
    .s(_1314_),
    .y(\DFF_392.D )
  );
  al_oa21ftf _3178_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_216.Q ),
    .y(_1315_)
  );
  al_aoi21 _3179_ (
    .a(_0006_),
    .b(_0896_),
    .c(_1315_),
    .y(\DFF_216.D )
  );
  al_nand2 _3180_ (
    .a(\DFF_432.Q ),
    .b(_1111_),
    .y(_1316_)
  );
  al_ao21ftf _3181_ (
    .a(_1111_),
    .b(\DFF_104.Q ),
    .c(_1316_),
    .y(\DFF_432.D )
  );
  al_inv _3182_ (
    .a(_0944_),
    .y(_1317_)
  );
  al_mux2l _3183_ (
    .a(_0480_),
    .b(_0474_),
    .s(_0945_),
    .y(_1318_)
  );
  al_aoi21ftt _3184_ (
    .a(_1011_),
    .b(_1317_),
    .c(_1318_),
    .y(_1319_)
  );
  al_and2 _3185_ (
    .a(\DFF_300.Q ),
    .b(_1319_),
    .y(_1320_)
  );
  al_or2 _3186_ (
    .a(\DFF_300.Q ),
    .b(_1319_),
    .y(_1321_)
  );
  al_nand2ft _3187_ (
    .a(_1320_),
    .b(_1321_),
    .y(_1322_)
  );
  al_ao21 _3188_ (
    .a(_0513_),
    .b(_1322_),
    .c(_0951_),
    .y(\DFF_300.D )
  );
  al_and3 _3189_ (
    .a(\DFF_367.Q ),
    .b(_0536_),
    .c(\DFF_37.D ),
    .y(_1323_)
  );
  al_ao21 _3190_ (
    .a(\DFF_181.Q ),
    .b(_0977_),
    .c(_1323_),
    .y(\DFF_181.D )
  );
  al_nand2 _3191_ (
    .a(\DFF_195.Q ),
    .b(_1111_),
    .y(_1324_)
  );
  al_ao21ftf _3192_ (
    .a(_1111_),
    .b(\DFF_324.Q ),
    .c(_1324_),
    .y(\DFF_195.D )
  );
  al_or3fft _3193_ (
    .a(\DFF_488.Q ),
    .b(_0800_),
    .c(_0954_),
    .y(_1325_)
  );
  al_ao21ftf _3194_ (
    .a(_1171_),
    .b(_0954_),
    .c(_1325_),
    .y(\DFF_488.D )
  );
  al_inv _3195_ (
    .a(\DFF_60.Q ),
    .y(_1326_)
  );
  al_or3fft _3196_ (
    .a(\DFF_521.Q ),
    .b(_0800_),
    .c(_0954_),
    .y(_1327_)
  );
  al_ao21ftf _3197_ (
    .a(_1326_),
    .b(_0954_),
    .c(_1327_),
    .y(\DFF_521.D )
  );
  al_nand2ft _3198_ (
    .a(\DFF_276.Q ),
    .b(\DFF_162.Q ),
    .y(_1328_)
  );
  al_ao21ttf _3199_ (
    .a(\DFF_276.Q ),
    .b(\DFF_465.Q ),
    .c(_1328_),
    .y(g6955)
  );
  al_or3 _3200_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_82.Q ),
    .y(_1329_)
  );
  al_mux2h _3201_ (
    .a(\DFF_87.Q ),
    .b(_0635_),
    .s(_1329_),
    .y(\DFF_87.D )
  );
  al_or3ftt _3202_ (
    .a(_1028_),
    .b(_0685_),
    .c(_0696_),
    .y(_1330_)
  );
  al_or2 _3203_ (
    .a(\DFF_60.Q ),
    .b(_1028_),
    .y(_1331_)
  );
  al_and3 _3204_ (
    .a(_1069_),
    .b(_1331_),
    .c(_1330_),
    .y(_1332_)
  );
  al_and2 _3205_ (
    .a(\DFF_450.Q ),
    .b(_1332_),
    .y(_1333_)
  );
  al_or2 _3206_ (
    .a(\DFF_450.Q ),
    .b(_1332_),
    .y(_1334_)
  );
  al_and2ft _3207_ (
    .a(_1333_),
    .b(_1334_),
    .y(_1335_)
  );
  al_ao21 _3208_ (
    .a(_1335_),
    .b(_1025_),
    .c(_1039_),
    .y(\DFF_450.D )
  );
  al_nand3 _3209_ (
    .a(\DFF_475.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1336_)
  );
  al_ao21ttf _3210_ (
    .a(\DFF_210.Q ),
    .b(_0355_),
    .c(_1336_),
    .y(\DFF_475.D )
  );
  al_ao21 _3211_ (
    .a(\DFF_323.Q ),
    .b(\DFF_320.Q ),
    .c(\DFF_388.Q ),
    .y(_1337_)
  );
  al_mux2h _3212_ (
    .a(\DFF_332.Q ),
    .b(_0966_),
    .s(_1337_),
    .y(\DFF_388.D )
  );
  al_nand3 _3213_ (
    .a(\DFF_210.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1338_)
  );
  al_ao21ttf _3214_ (
    .a(\DFF_522.Q ),
    .b(_0355_),
    .c(_1338_),
    .y(\DFF_210.D )
  );
  al_nand3 _3215_ (
    .a(_0635_),
    .b(_0601_),
    .c(_0806_),
    .y(_1339_)
  );
  al_aoi21ftf _3216_ (
    .a(\DFF_249.Q ),
    .b(_0841_),
    .c(_1339_),
    .y(\DFF_249.D )
  );
  al_nand2 _3217_ (
    .a(\DFF_227.Q ),
    .b(_0455_),
    .y(\DFF_227.D )
  );
  al_oai21ftf _3218_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_479.Q ),
    .y(\DFF_479.D )
  );
  al_nor3fft _3219_ (
    .a(\DFF_231.Q ),
    .b(\DFF_0.Q ),
    .c(_0443_),
    .y(_1340_)
  );
  al_ao21 _3220_ (
    .a(\DFF_355.Q ),
    .b(_0839_),
    .c(_1340_),
    .y(\DFF_355.D )
  );
  al_ao21 _3221_ (
    .a(\DFF_323.Q ),
    .b(\DFF_320.Q ),
    .c(\DFF_78.Q ),
    .y(_1341_)
  );
  al_mux2h _3222_ (
    .a(\DFF_104.Q ),
    .b(_0966_),
    .s(_1341_),
    .y(\DFF_78.D )
  );
  al_nand3ftt _3223_ (
    .a(\DFF_42.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1342_)
  );
  al_mux2h _3224_ (
    .a(\DFF_519.Q ),
    .b(_0961_),
    .s(_1342_),
    .y(\DFF_42.D )
  );
  al_nand2ft _3225_ (
    .a(\DFF_276.Q ),
    .b(\DFF_280.Q ),
    .y(_1343_)
  );
  al_ao21ttf _3226_ (
    .a(\DFF_276.Q ),
    .b(\DFF_206.Q ),
    .c(_1343_),
    .y(g6942)
  );
  al_nand2ft _3227_ (
    .a(\DFF_358.Q ),
    .b(\DFF_310.Q ),
    .y(_1344_)
  );
  al_nand2 _3228_ (
    .a(\DFF_362.Q ),
    .b(\DFF_358.Q ),
    .y(_1345_)
  );
  al_aoi21ttf _3229_ (
    .a(\DFF_135.Q ),
    .b(\DFF_261.Q ),
    .c(_1345_),
    .y(_1346_)
  );
  al_nand3fft _3230_ (
    .a(\DFF_72.Q ),
    .b(_0677_),
    .c(_1346_),
    .y(_1347_)
  );
  al_ao21ftf _3231_ (
    .a(_0689_),
    .b(_1344_),
    .c(_1347_),
    .y(_1348_)
  );
  al_nor3fft _3232_ (
    .a(\DFF_43.Q ),
    .b(\DFF_270.Q ),
    .c(_1348_),
    .y(_1349_)
  );
  al_and2 _3233_ (
    .a(\DFF_43.Q ),
    .b(\DFF_270.Q ),
    .y(_1350_)
  );
  al_or3fft _3234_ (
    .a(_1344_),
    .b(_1346_),
    .c(_1037_),
    .y(_1351_)
  );
  al_mux2h _3235_ (
    .a(_0762_),
    .b(_1351_),
    .s(\DFF_157.D ),
    .y(_1352_)
  );
  al_ao21ftf _3236_ (
    .a(_1350_),
    .b(_1348_),
    .c(_1352_),
    .y(_1353_)
  );
  al_mux2h _3237_ (
    .a(_1349_),
    .b(_1353_),
    .s(\DFF_360.Q ),
    .y(_1354_)
  );
  al_ao21ftf _3238_ (
    .a(\DFF_43.Q ),
    .b(_0681_),
    .c(_0800_),
    .y(_1355_)
  );
  al_ao21 _3239_ (
    .a(\DFF_99.Q ),
    .b(\DFF_387.Q ),
    .c(_0506_),
    .y(_1356_)
  );
  al_and2 _3240_ (
    .a(\DFF_127.Q ),
    .b(\DFF_389.Q ),
    .y(_1357_)
  );
  al_mux2h _3241_ (
    .a(_1100_),
    .b(_1357_),
    .s(\DFF_347.Q ),
    .y(_1358_)
  );
  al_and3ftt _3242_ (
    .a(_0800_),
    .b(_1356_),
    .c(_1358_),
    .y(_1359_)
  );
  al_mux2l _3243_ (
    .a(_1355_),
    .b(_1354_),
    .s(_1359_),
    .y(\DFF_360.D )
  );
  al_nand3ftt _3244_ (
    .a(\DFF_46.Q ),
    .b(g109),
    .c(_0589_),
    .y(_1360_)
  );
  al_mux2h _3245_ (
    .a(\DFF_490.Q ),
    .b(_0956_),
    .s(_1360_),
    .y(\DFF_46.D )
  );
  al_nand3 _3246_ (
    .a(\DFF_217.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1361_)
  );
  al_ao21ttf _3247_ (
    .a(\DFF_124.Q ),
    .b(_0355_),
    .c(_1361_),
    .y(\DFF_217.D )
  );
  al_nand3 _3248_ (
    .a(\DFF_329.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1362_)
  );
  al_ao21ttf _3249_ (
    .a(\DFF_151.Q ),
    .b(_0355_),
    .c(_1362_),
    .y(\DFF_329.D )
  );
  al_oai21ftf _3250_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_496.Q ),
    .y(\DFF_496.D )
  );
  al_nand3ftt _3251_ (
    .a(\DFF_425.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1363_)
  );
  al_mux2h _3252_ (
    .a(\DFF_235.Q ),
    .b(_0961_),
    .s(_1363_),
    .y(\DFF_425.D )
  );
  al_nand3ftt _3253_ (
    .a(\DFF_218.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1364_)
  );
  al_mux2h _3254_ (
    .a(\DFF_503.Q ),
    .b(_0961_),
    .s(_1364_),
    .y(\DFF_218.D )
  );
  al_nand2ft _3255_ (
    .a(\DFF_276.Q ),
    .b(\DFF_423.Q ),
    .y(_1365_)
  );
  al_ao21ttf _3256_ (
    .a(\DFF_276.Q ),
    .b(\DFF_26.Q ),
    .c(_1365_),
    .y(g6920)
  );
  al_nand2 _3257_ (
    .a(\DFF_448.Q ),
    .b(_1111_),
    .y(_1366_)
  );
  al_ao21ftf _3258_ (
    .a(_1111_),
    .b(\DFF_332.Q ),
    .c(_1366_),
    .y(\DFF_448.D )
  );
  al_ao21 _3259_ (
    .a(\DFF_323.Q ),
    .b(\DFF_320.Q ),
    .c(\DFF_200.Q ),
    .y(_1367_)
  );
  al_mux2h _3260_ (
    .a(\DFF_75.Q ),
    .b(_0966_),
    .s(_1367_),
    .y(\DFF_200.D )
  );
  al_mux2h _3261_ (
    .a(_0151_),
    .b(\DFF_22.D ),
    .s(_1042_),
    .y(_1368_)
  );
  al_ao21ftt _3262_ (
    .a(_0831_),
    .b(_1134_),
    .c(_1368_),
    .y(_1369_)
  );
  al_mux2l _3263_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .s(\DFF_524.Q ),
    .y(_1370_)
  );
  al_mux2l _3264_ (
    .a(_0841_),
    .b(_1369_),
    .s(_1370_),
    .y(\DFF_524.D )
  );
  al_or3 _3265_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_16.Q ),
    .y(_1371_)
  );
  al_mux2h _3266_ (
    .a(\DFF_167.Q ),
    .b(_0635_),
    .s(_1371_),
    .y(\DFF_167.D )
  );
  al_nand3ftt _3267_ (
    .a(\DFF_229.Q ),
    .b(g109),
    .c(_0589_),
    .y(_1372_)
  );
  al_mux2h _3268_ (
    .a(\DFF_296.Q ),
    .b(_0956_),
    .s(_1372_),
    .y(\DFF_229.D )
  );
  al_nand3 _3269_ (
    .a(\DFF_205.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1373_)
  );
  al_ao21ttf _3270_ (
    .a(\DFF_379.Q ),
    .b(_0355_),
    .c(_1373_),
    .y(\DFF_205.D )
  );
  al_or3 _3271_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_376.Q ),
    .y(_1374_)
  );
  al_mux2h _3272_ (
    .a(\DFF_413.Q ),
    .b(_0635_),
    .s(_1374_),
    .y(\DFF_413.D )
  );
  al_nand3 _3273_ (
    .a(_0635_),
    .b(_0708_),
    .c(_0725_),
    .y(_1375_)
  );
  al_aoi21ftf _3274_ (
    .a(\DFF_404.Q ),
    .b(_0841_),
    .c(_1375_),
    .y(\DFF_404.D )
  );
  al_ao21ftf _3275_ (
    .a(_0635_),
    .b(\DFF_50.Q ),
    .c(_1206_),
    .y(\DFF_50.D )
  );
  al_ao21 _3276_ (
    .a(_0481_),
    .b(_0475_),
    .c(_0945_),
    .y(_1376_)
  );
  al_aoi21ftf _3277_ (
    .a(_1272_),
    .b(_1317_),
    .c(_1376_),
    .y(_1377_)
  );
  al_and2 _3278_ (
    .a(_0465_),
    .b(_1377_),
    .y(_1378_)
  );
  al_or2 _3279_ (
    .a(_0465_),
    .b(_1377_),
    .y(_1379_)
  );
  al_nand3ftt _3280_ (
    .a(_1378_),
    .b(_1379_),
    .c(_0513_),
    .y(_1380_)
  );
  al_nand2ft _3281_ (
    .a(_0951_),
    .b(_1380_),
    .y(\DFF_212.D )
  );
  al_oa21ftf _3282_ (
    .a(\DFF_372.Q ),
    .b(g1696),
    .c(\DFF_423.Q ),
    .y(_1381_)
  );
  al_mux2l _3283_ (
    .a(_1133_),
    .b(_1369_),
    .s(_1381_),
    .y(\DFF_423.D )
  );
  al_nand2 _3284_ (
    .a(\DFF_342.Q ),
    .b(_1111_),
    .y(_1382_)
  );
  al_ao21ftf _3285_ (
    .a(_1111_),
    .b(\DFF_523.Q ),
    .c(_1382_),
    .y(\DFF_342.D )
  );
  al_or3fft _3286_ (
    .a(\DFF_427.Q ),
    .b(_0800_),
    .c(_0954_),
    .y(_1383_)
  );
  al_ao21ttf _3287_ (
    .a(\DFF_48.Q ),
    .b(_0954_),
    .c(_1383_),
    .y(\DFF_427.D )
  );
  al_nand3ftt _3288_ (
    .a(\DFF_130.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1384_)
  );
  al_mux2h _3289_ (
    .a(\DFF_237.Q ),
    .b(_0961_),
    .s(_1384_),
    .y(\DFF_130.D )
  );
  al_nand3 _3290_ (
    .a(\DFF_492.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1385_)
  );
  al_ao21ttf _3291_ (
    .a(\DFF_512.Q ),
    .b(_0355_),
    .c(_1385_),
    .y(\DFF_492.D )
  );
  al_nand3ftt _3292_ (
    .a(\DFF_176.Q ),
    .b(g109),
    .c(_0589_),
    .y(_1386_)
  );
  al_mux2h _3293_ (
    .a(\DFF_337.Q ),
    .b(_0956_),
    .s(_1386_),
    .y(\DFF_176.D )
  );
  al_nand3 _3294_ (
    .a(\DFF_430.Q ),
    .b(_0354_),
    .c(_0568_),
    .y(_1387_)
  );
  al_ao21ftf _3295_ (
    .a(_0931_),
    .b(_0355_),
    .c(_1387_),
    .y(\DFF_430.D )
  );
  al_or2 _3296_ (
    .a(\DFF_395.Q ),
    .b(_0684_),
    .y(_1388_)
  );
  al_nand2 _3297_ (
    .a(\DFF_395.Q ),
    .b(_0684_),
    .y(_1389_)
  );
  al_ao21ttf _3298_ (
    .a(_1389_),
    .b(_1388_),
    .c(_1028_),
    .y(_1390_)
  );
  al_or2ft _3299_ (
    .a(\DFF_488.Q ),
    .b(_1028_),
    .y(_1391_)
  );
  al_ao21ttf _3300_ (
    .a(_1391_),
    .b(_1390_),
    .c(_1069_),
    .y(_1392_)
  );
  al_or2 _3301_ (
    .a(_0695_),
    .b(_1392_),
    .y(_1393_)
  );
  al_and2 _3302_ (
    .a(_0695_),
    .b(_1392_),
    .y(_1394_)
  );
  al_and2ft _3303_ (
    .a(_1394_),
    .b(_1393_),
    .y(_1395_)
  );
  al_ao21 _3304_ (
    .a(_1395_),
    .b(_1025_),
    .c(_1039_),
    .y(\DFF_381.D )
  );
  al_nand2ft _3305_ (
    .a(g85),
    .b(g90),
    .y(_1396_)
  );
  al_ao21ttf _3306_ (
    .a(g85),
    .b(\DFF_439.Q ),
    .c(_1396_),
    .y(\DFF_439.D )
  );
  al_nand3ftt _3307_ (
    .a(\DFF_17.Q ),
    .b(g109),
    .c(_0656_),
    .y(_1397_)
  );
  al_mux2h _3308_ (
    .a(\DFF_494.Q ),
    .b(_0961_),
    .s(_1397_),
    .y(\DFF_17.D )
  );
  al_nand3ftt _3309_ (
    .a(\DFF_251.Q ),
    .b(g109),
    .c(_0589_),
    .y(_1398_)
  );
  al_mux2h _3310_ (
    .a(\DFF_444.Q ),
    .b(_0956_),
    .s(_1398_),
    .y(\DFF_251.D )
  );
  al_ao21ftt _3311_ (
    .a(_0472_),
    .b(\DFF_1.Q ),
    .c(_1116_),
    .y(_1399_)
  );
  al_nor2 _3312_ (
    .a(_1304_),
    .b(_0944_),
    .y(_1400_)
  );
  al_aoi21ftt _3313_ (
    .a(_0945_),
    .b(_1399_),
    .c(_1400_),
    .y(_1401_)
  );
  al_and2 _3314_ (
    .a(_0469_),
    .b(_1401_),
    .y(_1402_)
  );
  al_or2 _3315_ (
    .a(_0469_),
    .b(_1401_),
    .y(_1403_)
  );
  al_and2ft _3316_ (
    .a(_1402_),
    .b(_1403_),
    .y(_1404_)
  );
  al_ao21 _3317_ (
    .a(_1404_),
    .b(_0513_),
    .c(_0951_),
    .y(\DFF_354.D )
  );
  al_nand3ftt _3318_ (
    .a(\DFF_390.Q ),
    .b(g109),
    .c(_0589_),
    .y(_1405_)
  );
  al_mux2h _3319_ (
    .a(\DFF_190.Q ),
    .b(_0956_),
    .s(_1405_),
    .y(\DFF_390.D )
  );
  al_or3fft _3320_ (
    .a(\DFF_15.Q ),
    .b(_0800_),
    .c(_0954_),
    .y(_1406_)
  );
  al_ao21ttf _3321_ (
    .a(\DFF_281.Q ),
    .b(_0954_),
    .c(_1406_),
    .y(\DFF_15.D )
  );
  al_nand3ftt _3322_ (
    .a(\DFF_133.Q ),
    .b(g109),
    .c(_0589_),
    .y(_1407_)
  );
  al_mux2h _3323_ (
    .a(\DFF_102.Q ),
    .b(_0956_),
    .s(_1407_),
    .y(\DFF_133.D )
  );
  al_or3 _3324_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_170.Q ),
    .y(_1408_)
  );
  al_mux2h _3325_ (
    .a(\DFF_115.Q ),
    .b(_0635_),
    .s(_1408_),
    .y(\DFF_115.D )
  );
  al_ao21ftf _3326_ (
    .a(_0667_),
    .b(\DFF_196.Q ),
    .c(_0670_),
    .y(\DFF_196.D )
  );
  al_oa21ftt _3327_ (
    .a(\DFF_372.Q ),
    .b(g1696),
    .c(\DFF_94.Q ),
    .y(_1409_)
  );
  al_ao21 _3328_ (
    .a(\DFF_70.Q ),
    .b(_0958_),
    .c(_1409_),
    .y(\DFF_94.D )
  );
  al_nor3fft _3329_ (
    .a(\DFF_442.Q ),
    .b(\DFF_0.Q ),
    .c(_0443_),
    .y(_1410_)
  );
  al_ao21 _3330_ (
    .a(\DFF_58.Q ),
    .b(_0839_),
    .c(_1410_),
    .y(\DFF_58.D )
  );
  al_ao21 _3331_ (
    .a(\DFF_323.Q ),
    .b(\DFF_320.Q ),
    .c(\DFF_9.Q ),
    .y(_1411_)
  );
  al_mux2h _3332_ (
    .a(\DFF_523.Q ),
    .b(_0966_),
    .s(_1411_),
    .y(\DFF_9.D )
  );
  al_or3 _3333_ (
    .a(g1696),
    .b(\DFF_372.Q ),
    .c(\DFF_56.Q ),
    .y(_1412_)
  );
  al_mux2h _3334_ (
    .a(\DFF_108.Q ),
    .b(_0635_),
    .s(_1412_),
    .y(\DFF_108.D )
  );
  al_oa21ftf _3335_ (
    .a(g750),
    .b(\DFF_431.Q ),
    .c(\DFF_440.Q ),
    .y(_1413_)
  );
  al_aoi21 _3336_ (
    .a(_0006_),
    .b(_0887_),
    .c(_1413_),
    .y(\DFF_440.D )
  );
  al_nor3fft _3337_ (
    .a(\DFF_480.Q ),
    .b(\DFF_0.Q ),
    .c(_0443_),
    .y(_1414_)
  );
  al_ao21 _3338_ (
    .a(\DFF_510.Q ),
    .b(_0839_),
    .c(_1414_),
    .y(\DFF_510.D )
  );
  al_and2 _3339_ (
    .a(\DFF_54.Q ),
    .b(_0450_),
    .y(_1415_)
  );
  al_or2 _3340_ (
    .a(\DFF_54.Q ),
    .b(_0450_),
    .y(_1416_)
  );
  al_nand2ft _3341_ (
    .a(_1415_),
    .b(_1416_),
    .y(\DFF_269.D )
  );
  al_buf _3342_ (
    .a(\DFF_479.Q ),
    .y(g8982)
  );
  al_buf _3343_ (
    .a(\DFF_287.Q ),
    .y(g8980)
  );
  al_buf _3344_ (
    .a(\DFF_363.Q ),
    .y(g8986)
  );
  al_buf _3345_ (
    .a(\DFF_63.Q ),
    .y(g8977)
  );
  al_buf _3346_ (
    .a(\DFF_224.Q ),
    .y(g8983)
  );
  al_buf _3347_ (
    .a(\DFF_49.Q ),
    .y(g8985)
  );
  al_or3 _3348_ (
    .a(g41),
    .b(g31),
    .c(g30),
    .y(g9961)
  );
  al_buf _3349_ (
    .a(\DFF_91.Q ),
    .y(g8979)
  );
  al_buf _3350_ (
    .a(\DFF_513.Q ),
    .y(g8981)
  );
  al_buf _3351_ (
    .a(\DFF_533.Q ),
    .y(g8984)
  );
  al_buf _3352_ (
    .a(\DFF_496.Q ),
    .y(g8976)
  );
  al_buf _3353_ (
    .a(\DFF_213.Q ),
    .y(g8978)
  );
  al_dffl _3354_ (
    .clk(CK),
    .d(\DFF_0.D ),
    .q(\DFF_0.Q )
  );
  al_dffl _3355_ (
    .clk(CK),
    .d(\DFF_1.D ),
    .q(\DFF_1.Q )
  );
  al_dffl _3356_ (
    .clk(CK),
    .d(\DFF_270.Q ),
    .q(\DFF_2.Q )
  );
  al_dffl _3357_ (
    .clk(CK),
    .d(\DFF_3.D ),
    .q(\DFF_3.Q )
  );
  al_dffl _3358_ (
    .clk(CK),
    .d(\DFF_4.D ),
    .q(\DFF_4.Q )
  );
  al_dffl _3359_ (
    .clk(CK),
    .d(\DFF_5.D ),
    .q(\DFF_5.Q )
  );
  al_dffl _3360_ (
    .clk(CK),
    .d(\DFF_6.D ),
    .q(\DFF_6.Q )
  );
  al_dffl _3361_ (
    .clk(CK),
    .d(\DFF_7.D ),
    .q(\DFF_7.Q )
  );
  al_dffl _3362_ (
    .clk(CK),
    .d(\DFF_9.D ),
    .q(\DFF_9.Q )
  );
  al_dffl _3363_ (
    .clk(CK),
    .d(\DFF_10.D ),
    .q(\DFF_10.Q )
  );
  al_dffl _3364_ (
    .clk(CK),
    .d(\DFF_11.D ),
    .q(\DFF_11.Q )
  );
  al_dffl _3365_ (
    .clk(CK),
    .d(\DFF_12.D ),
    .q(\DFF_12.Q )
  );
  al_dffl _3366_ (
    .clk(CK),
    .d(\DFF_13.D ),
    .q(\DFF_13.Q )
  );
  al_dffl _3367_ (
    .clk(CK),
    .d(\DFF_14.D ),
    .q(\DFF_14.Q )
  );
  al_dffl _3368_ (
    .clk(CK),
    .d(\DFF_15.D ),
    .q(\DFF_15.Q )
  );
  al_dffl _3369_ (
    .clk(CK),
    .d(\DFF_16.D ),
    .q(\DFF_16.Q )
  );
  al_dffl _3370_ (
    .clk(CK),
    .d(\DFF_17.D ),
    .q(\DFF_17.Q )
  );
  al_dffl _3371_ (
    .clk(CK),
    .d(\DFF_18.D ),
    .q(\DFF_18.Q )
  );
  al_dffl _3372_ (
    .clk(CK),
    .d(\DFF_19.D ),
    .q(\DFF_19.Q )
  );
  al_dffl _3373_ (
    .clk(CK),
    .d(\DFF_20.D ),
    .q(\DFF_20.Q )
  );
  al_dffl _3374_ (
    .clk(CK),
    .d(\DFF_21.D ),
    .q(\DFF_21.Q )
  );
  al_dffl _3375_ (
    .clk(CK),
    .d(\DFF_22.D ),
    .q(\DFF_22.Q )
  );
  al_dffl _3376_ (
    .clk(CK),
    .d(\DFF_23.D ),
    .q(\DFF_23.Q )
  );
  al_dffl _3377_ (
    .clk(CK),
    .d(\DFF_24.D ),
    .q(\DFF_24.Q )
  );
  al_dffl _3378_ (
    .clk(CK),
    .d(\DFF_21.Q ),
    .q(\DFF_25.Q )
  );
  al_dffl _3379_ (
    .clk(CK),
    .d(\DFF_26.D ),
    .q(\DFF_26.Q )
  );
  al_dffl _3380_ (
    .clk(CK),
    .d(\DFF_27.D ),
    .q(\DFF_27.Q )
  );
  al_dffl _3381_ (
    .clk(CK),
    .d(\DFF_28.D ),
    .q(\DFF_28.Q )
  );
  al_dffl _3382_ (
    .clk(CK),
    .d(\DFF_29.D ),
    .q(\DFF_29.Q )
  );
  al_dffl _3383_ (
    .clk(CK),
    .d(\DFF_30.D ),
    .q(\DFF_30.Q )
  );
  al_dffl _3384_ (
    .clk(CK),
    .d(\DFF_31.D ),
    .q(\DFF_31.Q )
  );
  al_dffl _3385_ (
    .clk(CK),
    .d(\DFF_32.D ),
    .q(\DFF_32.Q )
  );
  al_dffl _3386_ (
    .clk(CK),
    .d(\DFF_33.D ),
    .q(\DFF_33.Q )
  );
  al_dffl _3387_ (
    .clk(CK),
    .d(\DFF_34.D ),
    .q(\DFF_34.Q )
  );
  al_dffl _3388_ (
    .clk(CK),
    .d(\DFF_35.D ),
    .q(\DFF_35.Q )
  );
  al_dffl _3389_ (
    .clk(CK),
    .d(\DFF_36.D ),
    .q(\DFF_36.Q )
  );
  al_dffl _3390_ (
    .clk(CK),
    .d(\DFF_37.D ),
    .q(\DFF_37.Q )
  );
  al_dffl _3391_ (
    .clk(CK),
    .d(\DFF_38.D ),
    .q(\DFF_38.Q )
  );
  al_dffl _3392_ (
    .clk(CK),
    .d(\DFF_39.D ),
    .q(\DFF_39.Q )
  );
  al_dffl _3393_ (
    .clk(CK),
    .d(\DFF_500.Q ),
    .q(\DFF_41.Q )
  );
  al_dffl _3394_ (
    .clk(CK),
    .d(\DFF_42.D ),
    .q(\DFF_42.Q )
  );
  al_dffl _3395_ (
    .clk(CK),
    .d(\DFF_43.D ),
    .q(\DFF_43.Q )
  );
  al_dffl _3396_ (
    .clk(CK),
    .d(\DFF_44.D ),
    .q(\DFF_44.Q )
  );
  al_dffl _3397_ (
    .clk(CK),
    .d(\DFF_45.D ),
    .q(\DFF_45.Q )
  );
  al_dffl _3398_ (
    .clk(CK),
    .d(\DFF_46.D ),
    .q(\DFF_46.Q )
  );
  al_dffl _3399_ (
    .clk(CK),
    .d(\DFF_47.D ),
    .q(\DFF_47.Q )
  );
  al_dffl _3400_ (
    .clk(CK),
    .d(\DFF_48.D ),
    .q(\DFF_48.Q )
  );
  al_dffl _3401_ (
    .clk(CK),
    .d(\DFF_49.D ),
    .q(\DFF_49.Q )
  );
  al_dffl _3402_ (
    .clk(CK),
    .d(\DFF_50.D ),
    .q(\DFF_50.Q )
  );
  al_dffl _3403_ (
    .clk(CK),
    .d(\DFF_51.D ),
    .q(\DFF_51.Q )
  );
  al_dffl _3404_ (
    .clk(CK),
    .d(\DFF_52.D ),
    .q(\DFF_52.Q )
  );
  al_dffl _3405_ (
    .clk(CK),
    .d(\DFF_53.D ),
    .q(\DFF_53.Q )
  );
  al_dffl _3406_ (
    .clk(CK),
    .d(\DFF_174.Q ),
    .q(\DFF_54.Q )
  );
  al_dffl _3407_ (
    .clk(CK),
    .d(\DFF_227.Q ),
    .q(\DFF_55.Q )
  );
  al_dffl _3408_ (
    .clk(CK),
    .d(\DFF_56.D ),
    .q(\DFF_56.Q )
  );
  al_dffl _3409_ (
    .clk(CK),
    .d(\DFF_57.D ),
    .q(\DFF_57.Q )
  );
  al_dffl _3410_ (
    .clk(CK),
    .d(\DFF_58.D ),
    .q(\DFF_58.Q )
  );
  al_dffl _3411_ (
    .clk(CK),
    .d(\DFF_59.D ),
    .q(\DFF_59.Q )
  );
  al_dffl _3412_ (
    .clk(CK),
    .d(\DFF_60.D ),
    .q(\DFF_60.Q )
  );
  al_dffl _3413_ (
    .clk(CK),
    .d(\DFF_61.D ),
    .q(\DFF_61.Q )
  );
  al_dffl _3414_ (
    .clk(CK),
    .d(\DFF_63.D ),
    .q(\DFF_63.Q )
  );
  al_dffl _3415_ (
    .clk(CK),
    .d(\DFF_64.D ),
    .q(\DFF_64.Q )
  );
  al_dffl _3416_ (
    .clk(CK),
    .d(\DFF_443.Q ),
    .q(\DFF_65.Q )
  );
  al_dffl _3417_ (
    .clk(CK),
    .d(\DFF_66.D ),
    .q(\DFF_66.Q )
  );
  al_dffl _3418_ (
    .clk(CK),
    .d(\DFF_67.D ),
    .q(\DFF_67.Q )
  );
  al_dffl _3419_ (
    .clk(CK),
    .d(\DFF_69.D ),
    .q(\DFF_69.Q )
  );
  al_dffl _3420_ (
    .clk(CK),
    .d(\DFF_70.D ),
    .q(\DFF_70.Q )
  );
  al_dffl _3421_ (
    .clk(CK),
    .d(\DFF_71.D ),
    .q(\DFF_71.Q )
  );
  al_dffl _3422_ (
    .clk(CK),
    .d(\DFF_72.D ),
    .q(\DFF_72.Q )
  );
  al_dffl _3423_ (
    .clk(CK),
    .d(\DFF_73.D ),
    .q(\DFF_73.Q )
  );
  al_dffl _3424_ (
    .clk(CK),
    .d(\DFF_74.D ),
    .q(\DFF_74.Q )
  );
  al_dffl _3425_ (
    .clk(CK),
    .d(\DFF_75.D ),
    .q(\DFF_75.Q )
  );
  al_dffl _3426_ (
    .clk(CK),
    .d(\DFF_76.D ),
    .q(\DFF_76.Q )
  );
  al_dffl _3427_ (
    .clk(CK),
    .d(\DFF_77.D ),
    .q(\DFF_77.Q )
  );
  al_dffl _3428_ (
    .clk(CK),
    .d(\DFF_78.D ),
    .q(\DFF_78.Q )
  );
  al_dffl _3429_ (
    .clk(CK),
    .d(\DFF_79.D ),
    .q(\DFF_79.Q )
  );
  al_dffl _3430_ (
    .clk(CK),
    .d(\DFF_81.D ),
    .q(\DFF_81.Q )
  );
  al_dffl _3431_ (
    .clk(CK),
    .d(\DFF_82.D ),
    .q(\DFF_82.Q )
  );
  al_dffl _3432_ (
    .clk(CK),
    .d(\DFF_83.D ),
    .q(\DFF_83.Q )
  );
  al_dffl _3433_ (
    .clk(CK),
    .d(\DFF_85.D ),
    .q(\DFF_85.Q )
  );
  al_dffl _3434_ (
    .clk(CK),
    .d(\DFF_86.D ),
    .q(\DFF_86.Q )
  );
  al_dffl _3435_ (
    .clk(CK),
    .d(\DFF_87.D ),
    .q(\DFF_87.Q )
  );
  al_dffl _3436_ (
    .clk(CK),
    .d(\DFF_88.D ),
    .q(\DFF_88.Q )
  );
  al_dffl _3437_ (
    .clk(CK),
    .d(\DFF_304.Q ),
    .q(\DFF_89.Q )
  );
  al_dffl _3438_ (
    .clk(CK),
    .d(\DFF_90.D ),
    .q(\DFF_90.Q )
  );
  al_dffl _3439_ (
    .clk(CK),
    .d(\DFF_91.D ),
    .q(\DFF_91.Q )
  );
  al_dffl _3440_ (
    .clk(CK),
    .d(\DFF_92.D ),
    .q(\DFF_92.Q )
  );
  al_dffl _3441_ (
    .clk(CK),
    .d(\DFF_53.Q ),
    .q(\DFF_93.Q )
  );
  al_dffl _3442_ (
    .clk(CK),
    .d(\DFF_94.D ),
    .q(\DFF_94.Q )
  );
  al_dffl _3443_ (
    .clk(CK),
    .d(\DFF_95.D ),
    .q(\DFF_95.Q )
  );
  al_dffl _3444_ (
    .clk(CK),
    .d(\DFF_96.D ),
    .q(\DFF_96.Q )
  );
  al_dffl _3445_ (
    .clk(CK),
    .d(\DFF_97.D ),
    .q(\DFF_97.Q )
  );
  al_dffl _3446_ (
    .clk(CK),
    .d(\DFF_98.D ),
    .q(\DFF_98.Q )
  );
  al_dffl _3447_ (
    .clk(CK),
    .d(\DFF_99.D ),
    .q(\DFF_99.Q )
  );
  al_dffl _3448_ (
    .clk(CK),
    .d(\DFF_101.D ),
    .q(\DFF_101.Q )
  );
  al_dffl _3449_ (
    .clk(CK),
    .d(\DFF_102.D ),
    .q(\DFF_102.Q )
  );
  al_dffl _3450_ (
    .clk(CK),
    .d(\DFF_103.D ),
    .q(\DFF_103.Q )
  );
  al_dffl _3451_ (
    .clk(CK),
    .d(\DFF_104.D ),
    .q(\DFF_104.Q )
  );
  al_dffl _3452_ (
    .clk(CK),
    .d(\DFF_105.D ),
    .q(\DFF_105.Q )
  );
  al_dffl _3453_ (
    .clk(CK),
    .d(\DFF_106.D ),
    .q(\DFF_106.Q )
  );
  al_dffl _3454_ (
    .clk(CK),
    .d(\DFF_108.D ),
    .q(\DFF_108.Q )
  );
  al_dffl _3455_ (
    .clk(CK),
    .d(\DFF_109.D ),
    .q(\DFF_109.Q )
  );
  al_dffl _3456_ (
    .clk(CK),
    .d(\DFF_110.D ),
    .q(\DFF_110.Q )
  );
  al_dffl _3457_ (
    .clk(CK),
    .d(\DFF_111.D ),
    .q(\DFF_111.Q )
  );
  al_dffl _3458_ (
    .clk(CK),
    .d(\DFF_112.D ),
    .q(\DFF_112.Q )
  );
  al_dffl _3459_ (
    .clk(CK),
    .d(\DFF_113.D ),
    .q(\DFF_113.Q )
  );
  al_dffl _3460_ (
    .clk(CK),
    .d(\DFF_114.D ),
    .q(\DFF_114.Q )
  );
  al_dffl _3461_ (
    .clk(CK),
    .d(\DFF_115.D ),
    .q(\DFF_115.Q )
  );
  al_dffl _3462_ (
    .clk(CK),
    .d(\DFF_116.D ),
    .q(\DFF_116.Q )
  );
  al_dffl _3463_ (
    .clk(CK),
    .d(\DFF_117.D ),
    .q(\DFF_117.Q )
  );
  al_dffl _3464_ (
    .clk(CK),
    .d(\DFF_118.D ),
    .q(\DFF_118.Q )
  );
  al_dffl _3465_ (
    .clk(CK),
    .d(\DFF_119.D ),
    .q(\DFF_119.Q )
  );
  al_dffl _3466_ (
    .clk(CK),
    .d(\DFF_120.D ),
    .q(\DFF_120.Q )
  );
  al_dffl _3467_ (
    .clk(CK),
    .d(\DFF_291.D ),
    .q(\DFF_291.Q )
  );
  al_dffl _3468_ (
    .clk(CK),
    .d(\DFF_291.Q ),
    .q(\DFF_121.Q )
  );
  al_dffl _3469_ (
    .clk(CK),
    .d(\DFF_122.D ),
    .q(\DFF_122.Q )
  );
  al_dffl _3470_ (
    .clk(CK),
    .d(\DFF_123.D ),
    .q(\DFF_123.Q )
  );
  al_dffl _3471_ (
    .clk(CK),
    .d(\DFF_124.D ),
    .q(\DFF_124.Q )
  );
  al_dffl _3472_ (
    .clk(CK),
    .d(\DFF_125.D ),
    .q(\DFF_125.Q )
  );
  al_dffl _3473_ (
    .clk(CK),
    .d(\DFF_526.D ),
    .q(\DFF_526.Q )
  );
  al_dffl _3474_ (
    .clk(CK),
    .d(\DFF_526.Q ),
    .q(\DFF_126.Q )
  );
  al_dffl _3475_ (
    .clk(CK),
    .d(\DFF_127.D ),
    .q(\DFF_127.Q )
  );
  al_dffl _3476_ (
    .clk(CK),
    .d(\DFF_128.D ),
    .q(\DFF_128.Q )
  );
  al_dffl _3477_ (
    .clk(CK),
    .d(\DFF_130.D ),
    .q(\DFF_130.Q )
  );
  al_dffl _3478_ (
    .clk(CK),
    .d(\DFF_131.D ),
    .q(\DFF_131.Q )
  );
  al_dffl _3479_ (
    .clk(CK),
    .d(\DFF_132.D ),
    .q(\DFF_132.Q )
  );
  al_dffl _3480_ (
    .clk(CK),
    .d(\DFF_133.D ),
    .q(\DFF_133.Q )
  );
  al_dffl _3481_ (
    .clk(CK),
    .d(\DFF_134.D ),
    .q(\DFF_134.Q )
  );
  al_dffl _3482_ (
    .clk(CK),
    .d(\DFF_135.D ),
    .q(\DFF_135.Q )
  );
  al_dffl _3483_ (
    .clk(CK),
    .d(\DFF_136.D ),
    .q(\DFF_136.Q )
  );
  al_dffl _3484_ (
    .clk(CK),
    .d(\DFF_137.D ),
    .q(\DFF_137.Q )
  );
  al_dffl _3485_ (
    .clk(CK),
    .d(\DFF_138.D ),
    .q(\DFF_138.Q )
  );
  al_dffl _3486_ (
    .clk(CK),
    .d(\DFF_139.D ),
    .q(\DFF_139.Q )
  );
  al_dffl _3487_ (
    .clk(CK),
    .d(\DFF_140.D ),
    .q(\DFF_140.Q )
  );
  al_dffl _3488_ (
    .clk(CK),
    .d(\DFF_141.D ),
    .q(\DFF_141.Q )
  );
  al_dffl _3489_ (
    .clk(CK),
    .d(\DFF_142.D ),
    .q(\DFF_142.Q )
  );
  al_dffl _3490_ (
    .clk(CK),
    .d(\DFF_143.D ),
    .q(\DFF_143.Q )
  );
  al_dffl _3491_ (
    .clk(CK),
    .d(\DFF_145.D ),
    .q(\DFF_145.Q )
  );
  al_dffl _3492_ (
    .clk(CK),
    .d(\DFF_146.D ),
    .q(\DFF_146.Q )
  );
  al_dffl _3493_ (
    .clk(CK),
    .d(\DFF_147.D ),
    .q(\DFF_147.Q )
  );
  al_dffl _3494_ (
    .clk(CK),
    .d(\DFF_148.D ),
    .q(\DFF_148.Q )
  );
  al_dffl _3495_ (
    .clk(CK),
    .d(\DFF_149.D ),
    .q(\DFF_149.Q )
  );
  al_dffl _3496_ (
    .clk(CK),
    .d(\DFF_151.D ),
    .q(\DFF_151.Q )
  );
  al_dffl _3497_ (
    .clk(CK),
    .d(\DFF_152.D ),
    .q(\DFF_152.Q )
  );
  al_dffl _3498_ (
    .clk(CK),
    .d(\DFF_153.D ),
    .q(\DFF_153.Q )
  );
  al_dffl _3499_ (
    .clk(CK),
    .d(\DFF_155.D ),
    .q(\DFF_155.Q )
  );
  al_dffl _3500_ (
    .clk(CK),
    .d(g83),
    .q(\DFF_462.Q )
  );
  al_dffl _3501_ (
    .clk(CK),
    .d(\DFF_462.Q ),
    .q(\DFF_156.Q )
  );
  al_dffl _3502_ (
    .clk(CK),
    .d(\DFF_157.D ),
    .q(\DFF_157.Q )
  );
  al_dffl _3503_ (
    .clk(CK),
    .d(\DFF_158.D ),
    .q(\DFF_158.Q )
  );
  al_dffl _3504_ (
    .clk(CK),
    .d(\DFF_159.D ),
    .q(\DFF_159.Q )
  );
  al_dffl _3505_ (
    .clk(CK),
    .d(\DFF_160.D ),
    .q(\DFF_160.Q )
  );
  al_dffl _3506_ (
    .clk(CK),
    .d(\DFF_161.D ),
    .q(\DFF_161.Q )
  );
  al_dffl _3507_ (
    .clk(CK),
    .d(\DFF_162.D ),
    .q(\DFF_162.Q )
  );
  al_dffl _3508_ (
    .clk(CK),
    .d(\DFF_163.D ),
    .q(\DFF_163.Q )
  );
  al_dffl _3509_ (
    .clk(CK),
    .d(\DFF_164.D ),
    .q(\DFF_164.Q )
  );
  al_dffl _3510_ (
    .clk(CK),
    .d(\DFF_165.D ),
    .q(\DFF_165.Q )
  );
  al_dffl _3511_ (
    .clk(CK),
    .d(\DFF_166.D ),
    .q(\DFF_166.Q )
  );
  al_dffl _3512_ (
    .clk(CK),
    .d(\DFF_167.D ),
    .q(\DFF_167.Q )
  );
  al_dffl _3513_ (
    .clk(CK),
    .d(\DFF_168.D ),
    .q(\DFF_168.Q )
  );
  al_dffl _3514_ (
    .clk(CK),
    .d(\DFF_169.D ),
    .q(\DFF_169.Q )
  );
  al_dffl _3515_ (
    .clk(CK),
    .d(\DFF_170.D ),
    .q(\DFF_170.Q )
  );
  al_dffl _3516_ (
    .clk(CK),
    .d(\DFF_171.D ),
    .q(\DFF_171.Q )
  );
  al_dffl _3517_ (
    .clk(CK),
    .d(\DFF_172.D ),
    .q(\DFF_172.Q )
  );
  al_dffl _3518_ (
    .clk(CK),
    .d(\DFF_173.D ),
    .q(\DFF_173.Q )
  );
  al_dffl _3519_ (
    .clk(CK),
    .d(\DFF_174.D ),
    .q(\DFF_174.Q )
  );
  al_dffl _3520_ (
    .clk(CK),
    .d(\DFF_222.Q ),
    .q(\DFF_175.Q )
  );
  al_dffl _3521_ (
    .clk(CK),
    .d(\DFF_176.D ),
    .q(\DFF_176.Q )
  );
  al_dffl _3522_ (
    .clk(CK),
    .d(\DFF_177.D ),
    .q(\DFF_177.Q )
  );
  al_dffl _3523_ (
    .clk(CK),
    .d(\DFF_178.D ),
    .q(\DFF_178.Q )
  );
  al_dffl _3524_ (
    .clk(CK),
    .d(\DFF_179.D ),
    .q(\DFF_179.Q )
  );
  al_dffl _3525_ (
    .clk(CK),
    .d(\DFF_180.D ),
    .q(\DFF_180.Q )
  );
  al_dffl _3526_ (
    .clk(CK),
    .d(\DFF_181.D ),
    .q(\DFF_181.Q )
  );
  al_dffl _3527_ (
    .clk(CK),
    .d(\DFF_182.D ),
    .q(\DFF_182.Q )
  );
  al_dffl _3528_ (
    .clk(CK),
    .d(\DFF_246.Q ),
    .q(\DFF_183.Q )
  );
  al_dffl _3529_ (
    .clk(CK),
    .d(\DFF_184.D ),
    .q(\DFF_184.Q )
  );
  al_dffl _3530_ (
    .clk(CK),
    .d(\DFF_185.D ),
    .q(\DFF_185.Q )
  );
  al_dffl _3531_ (
    .clk(CK),
    .d(\DFF_186.D ),
    .q(\DFF_186.Q )
  );
  al_dffl _3532_ (
    .clk(CK),
    .d(g103),
    .q(\DFF_187.Q )
  );
  al_dffl _3533_ (
    .clk(CK),
    .d(\DFF_398.D ),
    .q(\DFF_398.Q )
  );
  al_dffl _3534_ (
    .clk(CK),
    .d(\DFF_398.Q ),
    .q(\DFF_188.Q )
  );
  al_dffl _3535_ (
    .clk(CK),
    .d(\DFF_189.D ),
    .q(\DFF_189.Q )
  );
  al_dffl _3536_ (
    .clk(CK),
    .d(\DFF_190.D ),
    .q(\DFF_190.Q )
  );
  al_dffl _3537_ (
    .clk(CK),
    .d(\DFF_191.D ),
    .q(\DFF_191.Q )
  );
  al_dffl _3538_ (
    .clk(CK),
    .d(\DFF_192.D ),
    .q(\DFF_192.Q )
  );
  al_dffl _3539_ (
    .clk(CK),
    .d(\DFF_193.D ),
    .q(\DFF_193.Q )
  );
  al_dffl _3540_ (
    .clk(CK),
    .d(\DFF_328.D ),
    .q(\DFF_328.Q )
  );
  al_dffl _3541_ (
    .clk(CK),
    .d(\DFF_328.Q ),
    .q(\DFF_194.Q )
  );
  al_dffl _3542_ (
    .clk(CK),
    .d(\DFF_195.D ),
    .q(\DFF_195.Q )
  );
  al_dffl _3543_ (
    .clk(CK),
    .d(\DFF_196.D ),
    .q(\DFF_196.Q )
  );
  al_dffl _3544_ (
    .clk(CK),
    .d(\DFF_197.D ),
    .q(\DFF_197.Q )
  );
  al_dffl _3545_ (
    .clk(CK),
    .d(\DFF_198.D ),
    .q(\DFF_198.Q )
  );
  al_dffl _3546_ (
    .clk(CK),
    .d(\DFF_199.D ),
    .q(\DFF_199.Q )
  );
  al_dffl _3547_ (
    .clk(CK),
    .d(\DFF_200.D ),
    .q(\DFF_200.Q )
  );
  al_dffl _3548_ (
    .clk(CK),
    .d(\DFF_201.D ),
    .q(\DFF_201.Q )
  );
  al_dffl _3549_ (
    .clk(CK),
    .d(\DFF_202.D ),
    .q(\DFF_202.Q )
  );
  al_dffl _3550_ (
    .clk(CK),
    .d(\DFF_203.D ),
    .q(\DFF_203.Q )
  );
  al_dffl _3551_ (
    .clk(CK),
    .d(\DFF_204.D ),
    .q(\DFF_204.Q )
  );
  al_dffl _3552_ (
    .clk(CK),
    .d(\DFF_205.D ),
    .q(\DFF_205.Q )
  );
  al_dffl _3553_ (
    .clk(CK),
    .d(\DFF_206.D ),
    .q(\DFF_206.Q )
  );
  al_dffl _3554_ (
    .clk(CK),
    .d(\DFF_207.D ),
    .q(\DFF_207.Q )
  );
  al_dffl _3555_ (
    .clk(CK),
    .d(\DFF_208.D ),
    .q(\DFF_208.Q )
  );
  al_dffl _3556_ (
    .clk(CK),
    .d(\DFF_209.D ),
    .q(\DFF_209.Q )
  );
  al_dffl _3557_ (
    .clk(CK),
    .d(\DFF_210.D ),
    .q(\DFF_210.Q )
  );
  al_dffl _3558_ (
    .clk(CK),
    .d(\DFF_211.D ),
    .q(\DFF_211.Q )
  );
  al_dffl _3559_ (
    .clk(CK),
    .d(\DFF_212.D ),
    .q(\DFF_212.Q )
  );
  al_dffl _3560_ (
    .clk(CK),
    .d(\DFF_213.D ),
    .q(\DFF_213.Q )
  );
  al_dffl _3561_ (
    .clk(CK),
    .d(\DFF_214.D ),
    .q(\DFF_214.Q )
  );
  al_dffl _3562_ (
    .clk(CK),
    .d(\DFF_226.D ),
    .q(\DFF_226.Q )
  );
  al_dffl _3563_ (
    .clk(CK),
    .d(\DFF_226.Q ),
    .q(\DFF_215.Q )
  );
  al_dffl _3564_ (
    .clk(CK),
    .d(\DFF_216.D ),
    .q(\DFF_216.Q )
  );
  al_dffl _3565_ (
    .clk(CK),
    .d(\DFF_217.D ),
    .q(\DFF_217.Q )
  );
  al_dffl _3566_ (
    .clk(CK),
    .d(\DFF_218.D ),
    .q(\DFF_218.Q )
  );
  al_dffl _3567_ (
    .clk(CK),
    .d(\DFF_220.D ),
    .q(\DFF_220.Q )
  );
  al_dffl _3568_ (
    .clk(CK),
    .d(\DFF_221.D ),
    .q(\DFF_221.Q )
  );
  al_dffl _3569_ (
    .clk(CK),
    .d(\DFF_222.D ),
    .q(\DFF_222.Q )
  );
  al_dffl _3570_ (
    .clk(CK),
    .d(\DFF_223.D ),
    .q(\DFF_223.Q )
  );
  al_dffl _3571_ (
    .clk(CK),
    .d(\DFF_224.D ),
    .q(\DFF_224.Q )
  );
  al_dffl _3572_ (
    .clk(CK),
    .d(\DFF_356.Q ),
    .q(\DFF_225.Q )
  );
  al_dffl _3573_ (
    .clk(CK),
    .d(\DFF_227.D ),
    .q(\DFF_227.Q )
  );
  al_dffl _3574_ (
    .clk(CK),
    .d(\DFF_228.D ),
    .q(\DFF_228.Q )
  );
  al_dffl _3575_ (
    .clk(CK),
    .d(\DFF_229.D ),
    .q(\DFF_229.Q )
  );
  al_dffl _3576_ (
    .clk(CK),
    .d(\DFF_230.D ),
    .q(\DFF_230.Q )
  );
  al_dffl _3577_ (
    .clk(CK),
    .d(\DFF_231.D ),
    .q(\DFF_231.Q )
  );
  al_dffl _3578_ (
    .clk(CK),
    .d(\DFF_232.D ),
    .q(\DFF_232.Q )
  );
  al_dffl _3579_ (
    .clk(CK),
    .d(\DFF_318.Q ),
    .q(\DFF_233.Q )
  );
  al_dffl _3580_ (
    .clk(CK),
    .d(\DFF_234.D ),
    .q(\DFF_234.Q )
  );
  al_dffl _3581_ (
    .clk(CK),
    .d(\DFF_235.D ),
    .q(\DFF_235.Q )
  );
  al_dffl _3582_ (
    .clk(CK),
    .d(\DFF_236.D ),
    .q(\DFF_236.Q )
  );
  al_dffl _3583_ (
    .clk(CK),
    .d(\DFF_237.D ),
    .q(\DFF_237.Q )
  );
  al_dffl _3584_ (
    .clk(CK),
    .d(\DFF_238.D ),
    .q(\DFF_238.Q )
  );
  al_dffl _3585_ (
    .clk(CK),
    .d(\DFF_244.Q ),
    .q(\DFF_239.Q )
  );
  al_dffl _3586_ (
    .clk(CK),
    .d(\DFF_240.D ),
    .q(\DFF_240.Q )
  );
  al_dffl _3587_ (
    .clk(CK),
    .d(\DFF_241.D ),
    .q(\DFF_241.Q )
  );
  al_dffl _3588_ (
    .clk(CK),
    .d(\DFF_242.D ),
    .q(\DFF_242.Q )
  );
  al_dffl _3589_ (
    .clk(CK),
    .d(\DFF_243.D ),
    .q(\DFF_243.Q )
  );
  al_dffl _3590_ (
    .clk(CK),
    .d(\DFF_244.D ),
    .q(\DFF_244.Q )
  );
  al_dffl _3591_ (
    .clk(CK),
    .d(\DFF_245.D ),
    .q(\DFF_245.Q )
  );
  al_dffl _3592_ (
    .clk(CK),
    .d(\DFF_246.D ),
    .q(\DFF_246.Q )
  );
  al_dffl _3593_ (
    .clk(CK),
    .d(\DFF_247.D ),
    .q(\DFF_247.Q )
  );
  al_dffl _3594_ (
    .clk(CK),
    .d(\DFF_347.Q ),
    .q(\DFF_248.Q )
  );
  al_dffl _3595_ (
    .clk(CK),
    .d(\DFF_249.D ),
    .q(\DFF_249.Q )
  );
  al_dffl _3596_ (
    .clk(CK),
    .d(\DFF_250.D ),
    .q(\DFF_250.Q )
  );
  al_dffl _3597_ (
    .clk(CK),
    .d(\DFF_251.D ),
    .q(\DFF_251.Q )
  );
  al_dffl _3598_ (
    .clk(CK),
    .d(\DFF_252.D ),
    .q(\DFF_252.Q )
  );
  al_dffl _3599_ (
    .clk(CK),
    .d(\DFF_253.D ),
    .q(\DFF_253.Q )
  );
  al_dffl _3600_ (
    .clk(CK),
    .d(\DFF_254.D ),
    .q(\DFF_254.Q )
  );
  al_dffl _3601_ (
    .clk(CK),
    .d(\DFF_255.D ),
    .q(\DFF_255.Q )
  );
  al_dffl _3602_ (
    .clk(CK),
    .d(\DFF_256.D ),
    .q(\DFF_256.Q )
  );
  al_dffl _3603_ (
    .clk(CK),
    .d(\DFF_258.D ),
    .q(\DFF_258.Q )
  );
  al_dffl _3604_ (
    .clk(CK),
    .d(\DFF_259.D ),
    .q(\DFF_259.Q )
  );
  al_dffl _3605_ (
    .clk(CK),
    .d(\DFF_260.D ),
    .q(\DFF_260.Q )
  );
  al_dffl _3606_ (
    .clk(CK),
    .d(\DFF_261.D ),
    .q(\DFF_261.Q )
  );
  al_dffl _3607_ (
    .clk(CK),
    .d(\DFF_262.D ),
    .q(\DFF_262.Q )
  );
  al_dffl _3608_ (
    .clk(CK),
    .d(\DFF_263.D ),
    .q(\DFF_263.Q )
  );
  al_dffl _3609_ (
    .clk(CK),
    .d(\DFF_264.D ),
    .q(\DFF_264.Q )
  );
  al_dffl _3610_ (
    .clk(CK),
    .d(\DFF_397.Q ),
    .q(\DFF_265.Q )
  );
  al_dffl _3611_ (
    .clk(CK),
    .d(\DFF_266.D ),
    .q(\DFF_266.Q )
  );
  al_dffl _3612_ (
    .clk(CK),
    .d(\DFF_360.Q ),
    .q(\DFF_267.Q )
  );
  al_dffl _3613_ (
    .clk(CK),
    .d(\DFF_268.D ),
    .q(\DFF_268.Q )
  );
  al_dffl _3614_ (
    .clk(CK),
    .d(\DFF_269.D ),
    .q(\DFF_269.Q )
  );
  al_dffl _3615_ (
    .clk(CK),
    .d(\DFF_270.D ),
    .q(\DFF_270.Q )
  );
  al_dffl _3616_ (
    .clk(CK),
    .d(\DFF_271.D ),
    .q(\DFF_271.Q )
  );
  al_dffl _3617_ (
    .clk(CK),
    .d(\DFF_272.D ),
    .q(\DFF_272.Q )
  );
  al_dffl _3618_ (
    .clk(CK),
    .d(\DFF_273.D ),
    .q(\DFF_273.Q )
  );
  al_dffl _3619_ (
    .clk(CK),
    .d(\DFF_274.D ),
    .q(\DFF_274.Q )
  );
  al_dffl _3620_ (
    .clk(CK),
    .d(\DFF_275.D ),
    .q(\DFF_275.Q )
  );
  al_dffl _3621_ (
    .clk(CK),
    .d(\DFF_276.D ),
    .q(\DFF_276.Q )
  );
  al_dffl _3622_ (
    .clk(CK),
    .d(\DFF_277.D ),
    .q(\DFF_277.Q )
  );
  al_dffl _3623_ (
    .clk(CK),
    .d(\DFF_278.D ),
    .q(\DFF_278.Q )
  );
  al_dffl _3624_ (
    .clk(CK),
    .d(\DFF_279.D ),
    .q(\DFF_279.Q )
  );
  al_dffl _3625_ (
    .clk(CK),
    .d(\DFF_280.D ),
    .q(\DFF_280.Q )
  );
  al_dffl _3626_ (
    .clk(CK),
    .d(\DFF_281.D ),
    .q(\DFF_281.Q )
  );
  al_dffl _3627_ (
    .clk(CK),
    .d(\DFF_282.D ),
    .q(\DFF_282.Q )
  );
  al_dffl _3628_ (
    .clk(CK),
    .d(\DFF_283.D ),
    .q(\DFF_283.Q )
  );
  al_dffl _3629_ (
    .clk(CK),
    .d(\DFF_284.D ),
    .q(\DFF_284.Q )
  );
  al_dffl _3630_ (
    .clk(CK),
    .d(\DFF_285.D ),
    .q(\DFF_285.Q )
  );
  al_dffl _3631_ (
    .clk(CK),
    .d(\DFF_286.D ),
    .q(\DFF_286.Q )
  );
  al_dffl _3632_ (
    .clk(CK),
    .d(\DFF_287.D ),
    .q(\DFF_287.Q )
  );
  al_dffl _3633_ (
    .clk(CK),
    .d(\DFF_288.D ),
    .q(\DFF_288.Q )
  );
  al_dffl _3634_ (
    .clk(CK),
    .d(\DFF_289.D ),
    .q(\DFF_289.Q )
  );
  al_dffl _3635_ (
    .clk(CK),
    .d(\DFF_290.D ),
    .q(\DFF_290.Q )
  );
  al_dffl _3636_ (
    .clk(CK),
    .d(\DFF_292.D ),
    .q(\DFF_292.Q )
  );
  al_dffl _3637_ (
    .clk(CK),
    .d(\DFF_293.D ),
    .q(\DFF_293.Q )
  );
  al_dffl _3638_ (
    .clk(CK),
    .d(\DFF_294.D ),
    .q(\DFF_294.Q )
  );
  al_dffl _3639_ (
    .clk(CK),
    .d(\DFF_296.D ),
    .q(\DFF_296.Q )
  );
  al_dffl _3640_ (
    .clk(CK),
    .d(\DFF_297.D ),
    .q(\DFF_297.Q )
  );
  al_dffl _3641_ (
    .clk(CK),
    .d(\DFF_298.D ),
    .q(\DFF_298.Q )
  );
  al_dffl _3642_ (
    .clk(CK),
    .d(\DFF_137.Q ),
    .q(\DFF_299.Q )
  );
  al_dffl _3643_ (
    .clk(CK),
    .d(\DFF_300.D ),
    .q(\DFF_300.Q )
  );
  al_dffl _3644_ (
    .clk(CK),
    .d(\DFF_301.D ),
    .q(\DFF_301.Q )
  );
  al_dffl _3645_ (
    .clk(CK),
    .d(\DFF_302.D ),
    .q(\DFF_302.Q )
  );
  al_dffl _3646_ (
    .clk(CK),
    .d(\DFF_303.D ),
    .q(\DFF_303.Q )
  );
  al_dffl _3647_ (
    .clk(CK),
    .d(\DFF_156.Q ),
    .q(\DFF_304.Q )
  );
  al_dffl _3648_ (
    .clk(CK),
    .d(\DFF_305.D ),
    .q(\DFF_305.Q )
  );
  al_dffl _3649_ (
    .clk(CK),
    .d(\DFF_306.D ),
    .q(\DFF_306.Q )
  );
  al_dffl _3650_ (
    .clk(CK),
    .d(\DFF_307.D ),
    .q(\DFF_307.Q )
  );
  al_dffl _3651_ (
    .clk(CK),
    .d(\DFF_308.D ),
    .q(\DFF_308.Q )
  );
  al_dffl _3652_ (
    .clk(CK),
    .d(\DFF_389.Q ),
    .q(\DFF_309.Q )
  );
  al_dffl _3653_ (
    .clk(CK),
    .d(\DFF_310.D ),
    .q(\DFF_310.Q )
  );
  al_dffl _3654_ (
    .clk(CK),
    .d(\DFF_311.D ),
    .q(\DFF_311.Q )
  );
  al_dffl _3655_ (
    .clk(CK),
    .d(\DFF_312.D ),
    .q(\DFF_312.Q )
  );
  al_dffl _3656_ (
    .clk(CK),
    .d(\DFF_313.D ),
    .q(\DFF_313.Q )
  );
  al_dffl _3657_ (
    .clk(CK),
    .d(\DFF_314.D ),
    .q(\DFF_314.Q )
  );
  al_dffl _3658_ (
    .clk(CK),
    .d(\DFF_315.D ),
    .q(\DFF_315.Q )
  );
  al_dffl _3659_ (
    .clk(CK),
    .d(\DFF_316.D ),
    .q(\DFF_316.Q )
  );
  al_dffl _3660_ (
    .clk(CK),
    .d(\DFF_317.D ),
    .q(\DFF_317.Q )
  );
  al_dffl _3661_ (
    .clk(CK),
    .d(\DFF_318.D ),
    .q(\DFF_318.Q )
  );
  al_dffl _3662_ (
    .clk(CK),
    .d(\DFF_319.D ),
    .q(\DFF_319.Q )
  );
  al_dffl _3663_ (
    .clk(CK),
    .d(\DFF_320.D ),
    .q(\DFF_320.Q )
  );
  al_dffl _3664_ (
    .clk(CK),
    .d(\DFF_321.D ),
    .q(\DFF_321.Q )
  );
  al_dffl _3665_ (
    .clk(CK),
    .d(\DFF_322.D ),
    .q(\DFF_322.Q )
  );
  al_dffl _3666_ (
    .clk(CK),
    .d(\DFF_323.D ),
    .q(\DFF_323.Q )
  );
  al_dffl _3667_ (
    .clk(CK),
    .d(\DFF_324.D ),
    .q(\DFF_324.Q )
  );
  al_dffl _3668_ (
    .clk(CK),
    .d(\DFF_325.D ),
    .q(\DFF_325.Q )
  );
  al_dffl _3669_ (
    .clk(CK),
    .d(\DFF_326.D ),
    .q(\DFF_326.Q )
  );
  al_dffl _3670_ (
    .clk(CK),
    .d(\DFF_327.D ),
    .q(\DFF_327.Q )
  );
  al_dffl _3671_ (
    .clk(CK),
    .d(\DFF_329.D ),
    .q(\DFF_329.Q )
  );
  al_dffl _3672_ (
    .clk(CK),
    .d(\DFF_330.D ),
    .q(\DFF_330.Q )
  );
  al_dffl _3673_ (
    .clk(CK),
    .d(\DFF_331.D ),
    .q(\DFF_331.Q )
  );
  al_dffl _3674_ (
    .clk(CK),
    .d(\DFF_332.D ),
    .q(\DFF_332.Q )
  );
  al_dffl _3675_ (
    .clk(CK),
    .d(\DFF_333.D ),
    .q(\DFF_333.Q )
  );
  al_dffl _3676_ (
    .clk(CK),
    .d(\DFF_334.D ),
    .q(\DFF_334.Q )
  );
  al_dffl _3677_ (
    .clk(CK),
    .d(\DFF_335.D ),
    .q(\DFF_335.Q )
  );
  al_dffl _3678_ (
    .clk(CK),
    .d(\DFF_336.D ),
    .q(\DFF_336.Q )
  );
  al_dffl _3679_ (
    .clk(CK),
    .d(\DFF_337.D ),
    .q(\DFF_337.Q )
  );
  al_dffl _3680_ (
    .clk(CK),
    .d(\DFF_429.Q ),
    .q(\DFF_338.Q )
  );
  al_dffl _3681_ (
    .clk(CK),
    .d(\DFF_339.D ),
    .q(\DFF_339.Q )
  );
  al_dffl _3682_ (
    .clk(CK),
    .d(\DFF_340.D ),
    .q(\DFF_340.Q )
  );
  al_dffl _3683_ (
    .clk(CK),
    .d(\DFF_342.D ),
    .q(\DFF_342.Q )
  );
  al_dffl _3684_ (
    .clk(CK),
    .d(\DFF_184.Q ),
    .q(\DFF_343.Q )
  );
  al_dffl _3685_ (
    .clk(CK),
    .d(\DFF_344.D ),
    .q(\DFF_344.Q )
  );
  al_dffl _3686_ (
    .clk(CK),
    .d(\DFF_345.D ),
    .q(\DFF_345.Q )
  );
  al_dffl _3687_ (
    .clk(CK),
    .d(\DFF_346.D ),
    .q(\DFF_346.Q )
  );
  al_dffl _3688_ (
    .clk(CK),
    .d(\DFF_347.D ),
    .q(\DFF_347.Q )
  );
  al_dffl _3689_ (
    .clk(CK),
    .d(\DFF_348.D ),
    .q(\DFF_348.Q )
  );
  al_dffl _3690_ (
    .clk(CK),
    .d(\DFF_349.D ),
    .q(\DFF_349.Q )
  );
  al_dffl _3691_ (
    .clk(CK),
    .d(\DFF_350.D ),
    .q(\DFF_350.Q )
  );
  al_dffl _3692_ (
    .clk(CK),
    .d(\DFF_351.D ),
    .q(\DFF_351.Q )
  );
  al_dffl _3693_ (
    .clk(CK),
    .d(\DFF_352.D ),
    .q(\DFF_352.Q )
  );
  al_dffl _3694_ (
    .clk(CK),
    .d(\DFF_353.D ),
    .q(\DFF_353.Q )
  );
  al_dffl _3695_ (
    .clk(CK),
    .d(\DFF_354.D ),
    .q(\DFF_354.Q )
  );
  al_dffl _3696_ (
    .clk(CK),
    .d(\DFF_355.D ),
    .q(\DFF_355.Q )
  );
  al_dffl _3697_ (
    .clk(CK),
    .d(\DFF_356.D ),
    .q(\DFF_356.Q )
  );
  al_dffl _3698_ (
    .clk(CK),
    .d(\DFF_357.D ),
    .q(\DFF_357.Q )
  );
  al_dffl _3699_ (
    .clk(CK),
    .d(\DFF_358.D ),
    .q(\DFF_358.Q )
  );
  al_dffl _3700_ (
    .clk(CK),
    .d(\DFF_359.D ),
    .q(\DFF_359.Q )
  );
  al_dffl _3701_ (
    .clk(CK),
    .d(\DFF_360.D ),
    .q(\DFF_360.Q )
  );
  al_dffl _3702_ (
    .clk(CK),
    .d(\DFF_361.D ),
    .q(\DFF_361.Q )
  );
  al_dffl _3703_ (
    .clk(CK),
    .d(\DFF_362.D ),
    .q(\DFF_362.Q )
  );
  al_dffl _3704_ (
    .clk(CK),
    .d(\DFF_363.D ),
    .q(\DFF_363.Q )
  );
  al_dffl _3705_ (
    .clk(CK),
    .d(\DFF_364.D ),
    .q(\DFF_364.Q )
  );
  al_dffl _3706_ (
    .clk(CK),
    .d(\DFF_365.D ),
    .q(\DFF_365.Q )
  );
  al_dffl _3707_ (
    .clk(CK),
    .d(\DFF_366.D ),
    .q(\DFF_366.Q )
  );
  al_dffl _3708_ (
    .clk(CK),
    .d(\DFF_99.Q ),
    .q(\DFF_367.Q )
  );
  al_dffl _3709_ (
    .clk(CK),
    .d(\DFF_368.D ),
    .q(\DFF_368.Q )
  );
  al_dffl _3710_ (
    .clk(CK),
    .d(\DFF_369.D ),
    .q(\DFF_369.Q )
  );
  al_dffl _3711_ (
    .clk(CK),
    .d(\DFF_370.D ),
    .q(\DFF_370.Q )
  );
  al_dffl _3712_ (
    .clk(CK),
    .d(\DFF_371.D ),
    .q(\DFF_371.Q )
  );
  al_dffl _3713_ (
    .clk(CK),
    .d(\DFF_372.D ),
    .q(\DFF_372.Q )
  );
  al_dffl _3714_ (
    .clk(CK),
    .d(\DFF_373.D ),
    .q(\DFF_373.Q )
  );
  al_dffl _3715_ (
    .clk(CK),
    .d(\DFF_374.D ),
    .q(\DFF_374.Q )
  );
  al_dffl _3716_ (
    .clk(CK),
    .d(\DFF_376.D ),
    .q(\DFF_376.Q )
  );
  al_dffl _3717_ (
    .clk(CK),
    .d(\DFF_378.D ),
    .q(\DFF_378.Q )
  );
  al_dffl _3718_ (
    .clk(CK),
    .d(\DFF_379.D ),
    .q(\DFF_379.Q )
  );
  al_dffl _3719_ (
    .clk(CK),
    .d(\DFF_380.D ),
    .q(\DFF_380.Q )
  );
  al_dffl _3720_ (
    .clk(CK),
    .d(\DFF_381.D ),
    .q(\DFF_381.Q )
  );
  al_dffl _3721_ (
    .clk(CK),
    .d(\DFF_382.D ),
    .q(\DFF_382.Q )
  );
  al_dffl _3722_ (
    .clk(CK),
    .d(\DFF_383.D ),
    .q(\DFF_383.Q )
  );
  al_dffl _3723_ (
    .clk(CK),
    .d(\DFF_384.D ),
    .q(\DFF_384.Q )
  );
  al_dffl _3724_ (
    .clk(CK),
    .d(\DFF_385.D ),
    .q(\DFF_385.Q )
  );
  al_dffl _3725_ (
    .clk(CK),
    .d(\DFF_386.D ),
    .q(\DFF_386.Q )
  );
  al_dffl _3726_ (
    .clk(CK),
    .d(\DFF_387.D ),
    .q(\DFF_387.Q )
  );
  al_dffl _3727_ (
    .clk(CK),
    .d(\DFF_388.D ),
    .q(\DFF_388.Q )
  );
  al_dffl _3728_ (
    .clk(CK),
    .d(\DFF_389.D ),
    .q(\DFF_389.Q )
  );
  al_dffl _3729_ (
    .clk(CK),
    .d(\DFF_390.D ),
    .q(\DFF_390.Q )
  );
  al_dffl _3730_ (
    .clk(CK),
    .d(\DFF_391.D ),
    .q(\DFF_391.Q )
  );
  al_dffl _3731_ (
    .clk(CK),
    .d(\DFF_392.D ),
    .q(\DFF_392.Q )
  );
  al_dffl _3732_ (
    .clk(CK),
    .d(\DFF_393.D ),
    .q(\DFF_393.Q )
  );
  al_dffl _3733_ (
    .clk(CK),
    .d(\DFF_394.D ),
    .q(\DFF_394.Q )
  );
  al_dffl _3734_ (
    .clk(CK),
    .d(\DFF_395.D ),
    .q(\DFF_395.Q )
  );
  al_dffl _3735_ (
    .clk(CK),
    .d(\DFF_396.D ),
    .q(\DFF_396.Q )
  );
  al_dffl _3736_ (
    .clk(CK),
    .d(\DFF_397.D ),
    .q(\DFF_397.Q )
  );
  al_dffl _3737_ (
    .clk(CK),
    .d(\DFF_399.D ),
    .q(\DFF_399.Q )
  );
  al_dffl _3738_ (
    .clk(CK),
    .d(\DFF_400.D ),
    .q(\DFF_400.Q )
  );
  al_dffl _3739_ (
    .clk(CK),
    .d(\DFF_401.D ),
    .q(\DFF_401.Q )
  );
  al_dffl _3740_ (
    .clk(CK),
    .d(\DFF_402.D ),
    .q(\DFF_402.Q )
  );
  al_dffl _3741_ (
    .clk(CK),
    .d(\DFF_403.D ),
    .q(\DFF_403.Q )
  );
  al_dffl _3742_ (
    .clk(CK),
    .d(\DFF_404.D ),
    .q(\DFF_404.Q )
  );
  al_dffl _3743_ (
    .clk(CK),
    .d(\DFF_387.Q ),
    .q(\DFF_405.Q )
  );
  al_dffl _3744_ (
    .clk(CK),
    .d(\DFF_406.D ),
    .q(\DFF_406.Q )
  );
  al_dffl _3745_ (
    .clk(CK),
    .d(\DFF_407.D ),
    .q(\DFF_407.Q )
  );
  al_dffl _3746_ (
    .clk(CK),
    .d(\DFF_408.D ),
    .q(\DFF_408.Q )
  );
  al_dffl _3747_ (
    .clk(CK),
    .d(\DFF_409.D ),
    .q(\DFF_409.Q )
  );
  al_dffl _3748_ (
    .clk(CK),
    .d(\DFF_410.D ),
    .q(\DFF_410.Q )
  );
  al_dffl _3749_ (
    .clk(CK),
    .d(g29),
    .q(\DFF_411.Q )
  );
  al_dffl _3750_ (
    .clk(CK),
    .d(\DFF_127.Q ),
    .q(\DFF_412.Q )
  );
  al_dffl _3751_ (
    .clk(CK),
    .d(\DFF_413.D ),
    .q(\DFF_413.Q )
  );
  al_dffl _3752_ (
    .clk(CK),
    .d(\DFF_414.D ),
    .q(\DFF_414.Q )
  );
  al_dffl _3753_ (
    .clk(CK),
    .d(\DFF_415.D ),
    .q(\DFF_415.Q )
  );
  al_dffl _3754_ (
    .clk(CK),
    .d(\DFF_416.D ),
    .q(\DFF_416.Q )
  );
  al_dffl _3755_ (
    .clk(CK),
    .d(\DFF_417.D ),
    .q(\DFF_417.Q )
  );
  al_dffl _3756_ (
    .clk(CK),
    .d(\DFF_418.D ),
    .q(\DFF_418.Q )
  );
  al_dffl _3757_ (
    .clk(CK),
    .d(\DFF_419.D ),
    .q(\DFF_419.Q )
  );
  al_dffl _3758_ (
    .clk(CK),
    .d(\DFF_420.D ),
    .q(\DFF_420.Q )
  );
  al_dffl _3759_ (
    .clk(CK),
    .d(\DFF_421.D ),
    .q(\DFF_421.Q )
  );
  al_dffl _3760_ (
    .clk(CK),
    .d(\DFF_422.D ),
    .q(\DFF_422.Q )
  );
  al_dffl _3761_ (
    .clk(CK),
    .d(\DFF_423.D ),
    .q(\DFF_423.Q )
  );
  al_dffl _3762_ (
    .clk(CK),
    .d(\DFF_424.D ),
    .q(\DFF_424.Q )
  );
  al_dffl _3763_ (
    .clk(CK),
    .d(\DFF_425.D ),
    .q(\DFF_425.Q )
  );
  al_dffl _3764_ (
    .clk(CK),
    .d(\DFF_426.D ),
    .q(\DFF_426.Q )
  );
  al_dffl _3765_ (
    .clk(CK),
    .d(\DFF_427.D ),
    .q(\DFF_427.Q )
  );
  al_dffl _3766_ (
    .clk(CK),
    .d(\DFF_428.D ),
    .q(\DFF_428.Q )
  );
  al_dffl _3767_ (
    .clk(CK),
    .d(\DFF_429.D ),
    .q(\DFF_429.Q )
  );
  al_dffl _3768_ (
    .clk(CK),
    .d(\DFF_430.D ),
    .q(\DFF_430.Q )
  );
  al_dffl _3769_ (
    .clk(CK),
    .d(\DFF_431.D ),
    .q(\DFF_431.Q )
  );
  al_dffl _3770_ (
    .clk(CK),
    .d(\DFF_432.D ),
    .q(\DFF_432.Q )
  );
  al_dffl _3771_ (
    .clk(CK),
    .d(\DFF_393.Q ),
    .q(\DFF_433.Q )
  );
  al_dffl _3772_ (
    .clk(CK),
    .d(\DFF_434.D ),
    .q(\DFF_434.Q )
  );
  al_dffl _3773_ (
    .clk(CK),
    .d(\DFF_435.D ),
    .q(\DFF_435.Q )
  );
  al_dffl _3774_ (
    .clk(CK),
    .d(\DFF_71.Q ),
    .q(\DFF_436.Q )
  );
  al_dffl _3775_ (
    .clk(CK),
    .d(\DFF_437.D ),
    .q(\DFF_437.Q )
  );
  al_dffl _3776_ (
    .clk(CK),
    .d(\DFF_438.D ),
    .q(\DFF_438.Q )
  );
  al_dffl _3777_ (
    .clk(CK),
    .d(\DFF_439.D ),
    .q(\DFF_439.Q )
  );
  al_dffl _3778_ (
    .clk(CK),
    .d(\DFF_440.D ),
    .q(\DFF_440.Q )
  );
  al_dffl _3779_ (
    .clk(CK),
    .d(\DFF_357.Q ),
    .q(\DFF_441.Q )
  );
  al_dffl _3780_ (
    .clk(CK),
    .d(\DFF_442.D ),
    .q(\DFF_442.Q )
  );
  al_dffl _3781_ (
    .clk(CK),
    .d(\DFF_443.D ),
    .q(\DFF_443.Q )
  );
  al_dffl _3782_ (
    .clk(CK),
    .d(\DFF_444.D ),
    .q(\DFF_444.Q )
  );
  al_dffl _3783_ (
    .clk(CK),
    .d(\DFF_311.Q ),
    .q(\DFF_445.Q )
  );
  al_dffl _3784_ (
    .clk(CK),
    .d(\DFF_446.D ),
    .q(\DFF_446.Q )
  );
  al_dffl _3785_ (
    .clk(CK),
    .d(\DFF_447.D ),
    .q(\DFF_447.Q )
  );
  al_dffl _3786_ (
    .clk(CK),
    .d(\DFF_448.D ),
    .q(\DFF_448.Q )
  );
  al_dffl _3787_ (
    .clk(CK),
    .d(\DFF_449.D ),
    .q(\DFF_449.Q )
  );
  al_dffl _3788_ (
    .clk(CK),
    .d(\DFF_450.D ),
    .q(\DFF_450.Q )
  );
  al_dffl _3789_ (
    .clk(CK),
    .d(g28),
    .q(\DFF_451.Q )
  );
  al_dffl _3790_ (
    .clk(CK),
    .d(\DFF_452.D ),
    .q(\DFF_452.Q )
  );
  al_dffl _3791_ (
    .clk(CK),
    .d(\DFF_453.D ),
    .q(\DFF_453.Q )
  );
  al_dffl _3792_ (
    .clk(CK),
    .d(\DFF_454.D ),
    .q(\DFF_454.Q )
  );
  al_dffl _3793_ (
    .clk(CK),
    .d(\DFF_455.D ),
    .q(\DFF_455.Q )
  );
  al_dffl _3794_ (
    .clk(CK),
    .d(\DFF_456.D ),
    .q(\DFF_456.Q )
  );
  al_dffl _3795_ (
    .clk(CK),
    .d(\DFF_457.D ),
    .q(\DFF_457.Q )
  );
  al_dffl _3796_ (
    .clk(CK),
    .d(\DFF_458.D ),
    .q(\DFF_458.Q )
  );
  al_dffl _3797_ (
    .clk(CK),
    .d(\DFF_459.D ),
    .q(\DFF_459.Q )
  );
  al_dffl _3798_ (
    .clk(CK),
    .d(\DFF_460.D ),
    .q(\DFF_460.Q )
  );
  al_dffl _3799_ (
    .clk(CK),
    .d(\DFF_461.D ),
    .q(\DFF_461.Q )
  );
  al_dffl _3800_ (
    .clk(CK),
    .d(\DFF_463.D ),
    .q(\DFF_463.Q )
  );
  al_dffl _3801_ (
    .clk(CK),
    .d(g101),
    .q(\DFF_464.Q )
  );
  al_dffl _3802_ (
    .clk(CK),
    .d(\DFF_465.D ),
    .q(\DFF_465.Q )
  );
  al_dffl _3803_ (
    .clk(CK),
    .d(\DFF_466.D ),
    .q(\DFF_466.Q )
  );
  al_dffl _3804_ (
    .clk(CK),
    .d(\DFF_193.Q ),
    .q(\DFF_467.Q )
  );
  al_dffl _3805_ (
    .clk(CK),
    .d(\DFF_468.D ),
    .q(\DFF_468.Q )
  );
  al_dffl _3806_ (
    .clk(CK),
    .d(\DFF_470.D ),
    .q(\DFF_470.Q )
  );
  al_dffl _3807_ (
    .clk(CK),
    .d(\DFF_471.D ),
    .q(\DFF_471.Q )
  );
  al_dffl _3808_ (
    .clk(CK),
    .d(\DFF_472.D ),
    .q(\DFF_472.Q )
  );
  al_dffl _3809_ (
    .clk(CK),
    .d(\DFF_473.D ),
    .q(\DFF_473.Q )
  );
  al_dffl _3810_ (
    .clk(CK),
    .d(\DFF_474.D ),
    .q(\DFF_474.Q )
  );
  al_dffl _3811_ (
    .clk(CK),
    .d(\DFF_475.D ),
    .q(\DFF_475.Q )
  );
  al_dffl _3812_ (
    .clk(CK),
    .d(g104),
    .q(\DFF_476.Q )
  );
  al_dffl _3813_ (
    .clk(CK),
    .d(\DFF_477.D ),
    .q(\DFF_477.Q )
  );
  al_dffl _3814_ (
    .clk(CK),
    .d(\DFF_446.Q ),
    .q(\DFF_478.Q )
  );
  al_dffl _3815_ (
    .clk(CK),
    .d(\DFF_479.D ),
    .q(\DFF_479.Q )
  );
  al_dffl _3816_ (
    .clk(CK),
    .d(\DFF_480.D ),
    .q(\DFF_480.Q )
  );
  al_dffl _3817_ (
    .clk(CK),
    .d(\DFF_481.D ),
    .q(\DFF_481.Q )
  );
  al_dffl _3818_ (
    .clk(CK),
    .d(\DFF_482.D ),
    .q(\DFF_482.Q )
  );
  al_dffl _3819_ (
    .clk(CK),
    .d(\DFF_483.D ),
    .q(\DFF_483.Q )
  );
  al_dffl _3820_ (
    .clk(CK),
    .d(\DFF_484.D ),
    .q(\DFF_484.Q )
  );
  al_dffl _3821_ (
    .clk(CK),
    .d(\DFF_485.D ),
    .q(\DFF_485.Q )
  );
  al_dffl _3822_ (
    .clk(CK),
    .d(\DFF_486.D ),
    .q(\DFF_486.Q )
  );
  al_dffl _3823_ (
    .clk(CK),
    .d(\DFF_487.D ),
    .q(\DFF_487.Q )
  );
  al_dffl _3824_ (
    .clk(CK),
    .d(\DFF_488.D ),
    .q(\DFF_488.Q )
  );
  al_dffl _3825_ (
    .clk(CK),
    .d(\DFF_489.D ),
    .q(\DFF_489.Q )
  );
  al_dffl _3826_ (
    .clk(CK),
    .d(\DFF_490.D ),
    .q(\DFF_490.Q )
  );
  al_dffl _3827_ (
    .clk(CK),
    .d(\DFF_491.D ),
    .q(\DFF_491.Q )
  );
  al_dffl _3828_ (
    .clk(CK),
    .d(\DFF_492.D ),
    .q(\DFF_492.Q )
  );
  al_dffl _3829_ (
    .clk(CK),
    .d(\DFF_493.D ),
    .q(\DFF_493.Q )
  );
  al_dffl _3830_ (
    .clk(CK),
    .d(\DFF_494.D ),
    .q(\DFF_494.Q )
  );
  al_dffl _3831_ (
    .clk(CK),
    .d(\DFF_495.D ),
    .q(\DFF_495.Q )
  );
  al_dffl _3832_ (
    .clk(CK),
    .d(\DFF_496.D ),
    .q(\DFF_496.Q )
  );
  al_dffl _3833_ (
    .clk(CK),
    .d(\DFF_497.D ),
    .q(\DFF_497.Q )
  );
  al_dffl _3834_ (
    .clk(CK),
    .d(\DFF_498.D ),
    .q(\DFF_498.Q )
  );
  al_dffl _3835_ (
    .clk(CK),
    .d(\DFF_499.D ),
    .q(\DFF_499.Q )
  );
  al_dffl _3836_ (
    .clk(CK),
    .d(\DFF_500.D ),
    .q(\DFF_500.Q )
  );
  al_dffl _3837_ (
    .clk(CK),
    .d(\DFF_501.D ),
    .q(\DFF_501.Q )
  );
  al_dffl _3838_ (
    .clk(CK),
    .d(g102),
    .q(\DFF_502.Q )
  );
  al_dffl _3839_ (
    .clk(CK),
    .d(\DFF_503.D ),
    .q(\DFF_503.Q )
  );
  al_dffl _3840_ (
    .clk(CK),
    .d(\DFF_504.D ),
    .q(\DFF_504.Q )
  );
  al_dffl _3841_ (
    .clk(CK),
    .d(\DFF_505.D ),
    .q(\DFF_505.Q )
  );
  al_dffl _3842_ (
    .clk(CK),
    .d(\DFF_506.D ),
    .q(\DFF_506.Q )
  );
  al_dffl _3843_ (
    .clk(CK),
    .d(\DFF_507.D ),
    .q(\DFF_507.Q )
  );
  al_dffl _3844_ (
    .clk(CK),
    .d(\DFF_508.D ),
    .q(\DFF_508.Q )
  );
  al_dffl _3845_ (
    .clk(CK),
    .d(\DFF_509.D ),
    .q(\DFF_509.Q )
  );
  al_dffl _3846_ (
    .clk(CK),
    .d(\DFF_510.D ),
    .q(\DFF_510.Q )
  );
  al_dffl _3847_ (
    .clk(CK),
    .d(\DFF_511.D ),
    .q(\DFF_511.Q )
  );
  al_dffl _3848_ (
    .clk(CK),
    .d(\DFF_512.D ),
    .q(\DFF_512.Q )
  );
  al_dffl _3849_ (
    .clk(CK),
    .d(\DFF_513.D ),
    .q(\DFF_513.Q )
  );
  al_dffl _3850_ (
    .clk(CK),
    .d(\DFF_514.D ),
    .q(\DFF_514.Q )
  );
  al_dffl _3851_ (
    .clk(CK),
    .d(\DFF_515.D ),
    .q(\DFF_515.Q )
  );
  al_dffl _3852_ (
    .clk(CK),
    .d(\DFF_516.D ),
    .q(\DFF_516.Q )
  );
  al_dffl _3853_ (
    .clk(CK),
    .d(\DFF_517.D ),
    .q(\DFF_517.Q )
  );
  al_dffl _3854_ (
    .clk(CK),
    .d(\DFF_518.D ),
    .q(\DFF_518.Q )
  );
  al_dffl _3855_ (
    .clk(CK),
    .d(\DFF_519.D ),
    .q(\DFF_519.Q )
  );
  al_dffl _3856_ (
    .clk(CK),
    .d(\DFF_520.D ),
    .q(\DFF_520.Q )
  );
  al_dffl _3857_ (
    .clk(CK),
    .d(\DFF_521.D ),
    .q(\DFF_521.Q )
  );
  al_dffl _3858_ (
    .clk(CK),
    .d(\DFF_522.D ),
    .q(\DFF_522.Q )
  );
  al_dffl _3859_ (
    .clk(CK),
    .d(\DFF_523.D ),
    .q(\DFF_523.Q )
  );
  al_dffl _3860_ (
    .clk(CK),
    .d(\DFF_524.D ),
    .q(\DFF_524.Q )
  );
  al_dffl _3861_ (
    .clk(CK),
    .d(\DFF_525.D ),
    .q(\DFF_525.Q )
  );
  al_dffl _3862_ (
    .clk(CK),
    .d(\DFF_527.D ),
    .q(\DFF_527.Q )
  );
  al_dffl _3863_ (
    .clk(CK),
    .d(\DFF_528.D ),
    .q(\DFF_528.Q )
  );
  al_dffl _3864_ (
    .clk(CK),
    .d(\DFF_529.D ),
    .q(\DFF_529.Q )
  );
  al_dffl _3865_ (
    .clk(CK),
    .d(\DFF_530.D ),
    .q(\DFF_530.Q )
  );
  al_dffl _3866_ (
    .clk(CK),
    .d(\DFF_531.D ),
    .q(\DFF_531.Q )
  );
  al_dffl _3867_ (
    .clk(CK),
    .d(\DFF_532.D ),
    .q(\DFF_532.Q )
  );
  al_dffl _3868_ (
    .clk(CK),
    .d(\DFF_533.D ),
    .q(\DFF_533.Q )
  );
  assign \DFF_0.CK  = CK;
  assign \DFF_1.CK  = CK;
  assign \DFF_10.CK  = CK;
  assign \DFF_100.CK  = CK;
  assign \DFF_100.D  = g29;
  assign \DFF_100.Q  = \DFF_411.Q ;
  assign \DFF_101.CK  = CK;
  assign \DFF_102.CK  = CK;
  assign \DFF_103.CK  = CK;
  assign \DFF_104.CK  = CK;
  assign \DFF_105.CK  = CK;
  assign \DFF_106.CK  = CK;
  assign \DFF_107.CK  = CK;
  assign \DFF_108.CK  = CK;
  assign \DFF_109.CK  = CK;
  assign \DFF_11.CK  = CK;
  assign \DFF_110.CK  = CK;
  assign \DFF_111.CK  = CK;
  assign \DFF_112.CK  = CK;
  assign \DFF_113.CK  = CK;
  assign \DFF_114.CK  = CK;
  assign \DFF_115.CK  = CK;
  assign \DFF_116.CK  = CK;
  assign \DFF_117.CK  = CK;
  assign \DFF_118.CK  = CK;
  assign \DFF_119.CK  = CK;
  assign \DFF_12.CK  = CK;
  assign \DFF_120.CK  = CK;
  assign \DFF_121.CK  = CK;
  assign \DFF_121.D  = \DFF_291.Q ;
  assign \DFF_122.CK  = CK;
  assign \DFF_123.CK  = CK;
  assign \DFF_124.CK  = CK;
  assign \DFF_125.CK  = CK;
  assign \DFF_126.CK  = CK;
  assign \DFF_126.D  = \DFF_526.Q ;
  assign \DFF_127.CK  = CK;
  assign \DFF_128.CK  = CK;
  assign \DFF_129.CK  = CK;
  assign \DFF_129.D  = g102;
  assign \DFF_129.Q  = \DFF_502.Q ;
  assign \DFF_13.CK  = CK;
  assign \DFF_130.CK  = CK;
  assign \DFF_131.CK  = CK;
  assign \DFF_132.CK  = CK;
  assign \DFF_133.CK  = CK;
  assign \DFF_134.CK  = CK;
  assign \DFF_135.CK  = CK;
  assign \DFF_136.CK  = CK;
  assign \DFF_137.CK  = CK;
  assign \DFF_138.CK  = CK;
  assign \DFF_139.CK  = CK;
  assign \DFF_14.CK  = CK;
  assign \DFF_140.CK  = CK;
  assign \DFF_141.CK  = CK;
  assign \DFF_142.CK  = CK;
  assign \DFF_143.CK  = CK;
  assign \DFF_144.CK  = CK;
  assign \DFF_145.CK  = CK;
  assign \DFF_146.CK  = CK;
  assign \DFF_147.CK  = CK;
  assign \DFF_148.CK  = CK;
  assign \DFF_149.CK  = CK;
  assign \DFF_15.CK  = CK;
  assign \DFF_150.CK  = CK;
  assign \DFF_150.D  = g28;
  assign \DFF_150.Q  = \DFF_451.Q ;
  assign \DFF_151.CK  = CK;
  assign \DFF_152.CK  = CK;
  assign \DFF_153.CK  = CK;
  assign \DFF_154.CK  = CK;
  assign \DFF_154.D  = g103;
  assign \DFF_154.Q  = \DFF_187.Q ;
  assign \DFF_155.CK  = CK;
  assign \DFF_156.CK  = CK;
  assign \DFF_156.D  = \DFF_462.Q ;
  assign \DFF_157.CK  = CK;
  assign \DFF_158.CK  = CK;
  assign \DFF_159.CK  = CK;
  assign \DFF_16.CK  = CK;
  assign \DFF_160.CK  = CK;
  assign \DFF_161.CK  = CK;
  assign \DFF_162.CK  = CK;
  assign \DFF_163.CK  = CK;
  assign \DFF_164.CK  = CK;
  assign \DFF_165.CK  = CK;
  assign \DFF_166.CK  = CK;
  assign \DFF_167.CK  = CK;
  assign \DFF_168.CK  = CK;
  assign \DFF_169.CK  = CK;
  assign \DFF_17.CK  = CK;
  assign \DFF_170.CK  = CK;
  assign \DFF_171.CK  = CK;
  assign \DFF_172.CK  = CK;
  assign \DFF_173.CK  = CK;
  assign \DFF_174.CK  = CK;
  assign \DFF_175.CK  = CK;
  assign \DFF_175.D  = \DFF_222.Q ;
  assign \DFF_176.CK  = CK;
  assign \DFF_177.CK  = CK;
  assign \DFF_178.CK  = CK;
  assign \DFF_179.CK  = CK;
  assign \DFF_18.CK  = CK;
  assign \DFF_180.CK  = CK;
  assign \DFF_181.CK  = CK;
  assign \DFF_182.CK  = CK;
  assign \DFF_183.CK  = CK;
  assign \DFF_183.D  = \DFF_246.Q ;
  assign \DFF_184.CK  = CK;
  assign \DFF_185.CK  = CK;
  assign \DFF_186.CK  = CK;
  assign \DFF_187.CK  = CK;
  assign \DFF_187.D  = g103;
  assign \DFF_188.CK  = CK;
  assign \DFF_188.D  = \DFF_398.Q ;
  assign \DFF_189.CK  = CK;
  assign \DFF_19.CK  = CK;
  assign \DFF_190.CK  = CK;
  assign \DFF_191.CK  = CK;
  assign \DFF_192.CK  = CK;
  assign \DFF_193.CK  = CK;
  assign \DFF_194.CK  = CK;
  assign \DFF_194.D  = \DFF_328.Q ;
  assign \DFF_195.CK  = CK;
  assign \DFF_196.CK  = CK;
  assign \DFF_197.CK  = CK;
  assign \DFF_198.CK  = CK;
  assign \DFF_199.CK  = CK;
  assign \DFF_2.CK  = CK;
  assign \DFF_2.D  = \DFF_270.Q ;
  assign \DFF_20.CK  = CK;
  assign \DFF_200.CK  = CK;
  assign \DFF_201.CK  = CK;
  assign \DFF_202.CK  = CK;
  assign \DFF_203.CK  = CK;
  assign \DFF_204.CK  = CK;
  assign \DFF_205.CK  = CK;
  assign \DFF_206.CK  = CK;
  assign \DFF_207.CK  = CK;
  assign \DFF_208.CK  = CK;
  assign \DFF_209.CK  = CK;
  assign \DFF_21.CK  = CK;
  assign \DFF_210.CK  = CK;
  assign \DFF_211.CK  = CK;
  assign \DFF_212.CK  = CK;
  assign \DFF_213.CK  = CK;
  assign \DFF_214.CK  = CK;
  assign \DFF_215.CK  = CK;
  assign \DFF_215.D  = \DFF_226.Q ;
  assign \DFF_216.CK  = CK;
  assign \DFF_217.CK  = CK;
  assign \DFF_218.CK  = CK;
  assign \DFF_219.CK  = CK;
  assign \DFF_22.CK  = CK;
  assign \DFF_220.CK  = CK;
  assign \DFF_221.CK  = CK;
  assign \DFF_222.CK  = CK;
  assign \DFF_223.CK  = CK;
  assign \DFF_224.CK  = CK;
  assign \DFF_225.CK  = CK;
  assign \DFF_225.D  = \DFF_356.Q ;
  assign \DFF_226.CK  = CK;
  assign \DFF_227.CK  = CK;
  assign \DFF_228.CK  = CK;
  assign \DFF_229.CK  = CK;
  assign \DFF_23.CK  = CK;
  assign \DFF_230.CK  = CK;
  assign \DFF_231.CK  = CK;
  assign \DFF_232.CK  = CK;
  assign \DFF_233.CK  = CK;
  assign \DFF_233.D  = \DFF_318.Q ;
  assign \DFF_234.CK  = CK;
  assign \DFF_235.CK  = CK;
  assign \DFF_236.CK  = CK;
  assign \DFF_237.CK  = CK;
  assign \DFF_238.CK  = CK;
  assign \DFF_239.CK  = CK;
  assign \DFF_239.D  = \DFF_244.Q ;
  assign \DFF_24.CK  = CK;
  assign \DFF_240.CK  = CK;
  assign \DFF_241.CK  = CK;
  assign \DFF_242.CK  = CK;
  assign \DFF_243.CK  = CK;
  assign \DFF_244.CK  = CK;
  assign \DFF_245.CK  = CK;
  assign \DFF_246.CK  = CK;
  assign \DFF_247.CK  = CK;
  assign \DFF_248.CK  = CK;
  assign \DFF_248.D  = \DFF_347.Q ;
  assign \DFF_249.CK  = CK;
  assign \DFF_25.CK  = CK;
  assign \DFF_25.D  = \DFF_21.Q ;
  assign \DFF_250.CK  = CK;
  assign \DFF_251.CK  = CK;
  assign \DFF_252.CK  = CK;
  assign \DFF_253.CK  = CK;
  assign \DFF_254.CK  = CK;
  assign \DFF_255.CK  = CK;
  assign \DFF_256.CK  = CK;
  assign \DFF_257.CK  = CK;
  assign \DFF_258.CK  = CK;
  assign \DFF_259.CK  = CK;
  assign \DFF_26.CK  = CK;
  assign \DFF_260.CK  = CK;
  assign \DFF_261.CK  = CK;
  assign \DFF_262.CK  = CK;
  assign \DFF_263.CK  = CK;
  assign \DFF_264.CK  = CK;
  assign \DFF_265.CK  = CK;
  assign \DFF_265.D  = \DFF_397.Q ;
  assign \DFF_266.CK  = CK;
  assign \DFF_267.CK  = CK;
  assign \DFF_267.D  = \DFF_360.Q ;
  assign \DFF_268.CK  = CK;
  assign \DFF_269.CK  = CK;
  assign \DFF_27.CK  = CK;
  assign \DFF_270.CK  = CK;
  assign \DFF_271.CK  = CK;
  assign \DFF_272.CK  = CK;
  assign \DFF_273.CK  = CK;
  assign \DFF_274.CK  = CK;
  assign \DFF_275.CK  = CK;
  assign \DFF_276.CK  = CK;
  assign \DFF_277.CK  = CK;
  assign \DFF_278.CK  = CK;
  assign \DFF_279.CK  = CK;
  assign \DFF_28.CK  = CK;
  assign \DFF_280.CK  = CK;
  assign \DFF_281.CK  = CK;
  assign \DFF_282.CK  = CK;
  assign \DFF_283.CK  = CK;
  assign \DFF_284.CK  = CK;
  assign \DFF_285.CK  = CK;
  assign \DFF_286.CK  = CK;
  assign \DFF_287.CK  = CK;
  assign \DFF_288.CK  = CK;
  assign \DFF_289.CK  = CK;
  assign \DFF_29.CK  = CK;
  assign \DFF_290.CK  = CK;
  assign \DFF_291.CK  = CK;
  assign \DFF_292.CK  = CK;
  assign \DFF_293.CK  = CK;
  assign \DFF_294.CK  = CK;
  assign \DFF_295.CK  = CK;
  assign \DFF_295.D  = g83;
  assign \DFF_295.Q  = \DFF_462.Q ;
  assign \DFF_296.CK  = CK;
  assign \DFF_297.CK  = CK;
  assign \DFF_298.CK  = CK;
  assign \DFF_299.CK  = CK;
  assign \DFF_299.D  = \DFF_137.Q ;
  assign \DFF_3.CK  = CK;
  assign \DFF_30.CK  = CK;
  assign \DFF_300.CK  = CK;
  assign \DFF_301.CK  = CK;
  assign \DFF_302.CK  = CK;
  assign \DFF_303.CK  = CK;
  assign \DFF_304.CK  = CK;
  assign \DFF_304.D  = \DFF_156.Q ;
  assign \DFF_305.CK  = CK;
  assign \DFF_306.CK  = CK;
  assign \DFF_307.CK  = CK;
  assign \DFF_308.CK  = CK;
  assign \DFF_309.CK  = CK;
  assign \DFF_309.D  = \DFF_389.Q ;
  assign \DFF_31.CK  = CK;
  assign \DFF_310.CK  = CK;
  assign \DFF_311.CK  = CK;
  assign \DFF_312.CK  = CK;
  assign \DFF_313.CK  = CK;
  assign \DFF_314.CK  = CK;
  assign \DFF_315.CK  = CK;
  assign \DFF_316.CK  = CK;
  assign \DFF_317.CK  = CK;
  assign \DFF_318.CK  = CK;
  assign \DFF_319.CK  = CK;
  assign \DFF_32.CK  = CK;
  assign \DFF_320.CK  = CK;
  assign \DFF_321.CK  = CK;
  assign \DFF_322.CK  = CK;
  assign \DFF_323.CK  = CK;
  assign \DFF_324.CK  = CK;
  assign \DFF_325.CK  = CK;
  assign \DFF_326.CK  = CK;
  assign \DFF_327.CK  = CK;
  assign \DFF_328.CK  = CK;
  assign \DFF_329.CK  = CK;
  assign \DFF_33.CK  = CK;
  assign \DFF_330.CK  = CK;
  assign \DFF_331.CK  = CK;
  assign \DFF_332.CK  = CK;
  assign \DFF_333.CK  = CK;
  assign \DFF_334.CK  = CK;
  assign \DFF_335.CK  = CK;
  assign \DFF_336.CK  = CK;
  assign \DFF_337.CK  = CK;
  assign \DFF_338.CK  = CK;
  assign \DFF_338.D  = \DFF_429.Q ;
  assign \DFF_339.CK  = CK;
  assign \DFF_34.CK  = CK;
  assign \DFF_340.CK  = CK;
  assign \DFF_341.CK  = CK;
  assign \DFF_342.CK  = CK;
  assign \DFF_343.CK  = CK;
  assign \DFF_343.D  = \DFF_184.Q ;
  assign \DFF_344.CK  = CK;
  assign \DFF_345.CK  = CK;
  assign \DFF_346.CK  = CK;
  assign \DFF_347.CK  = CK;
  assign \DFF_348.CK  = CK;
  assign \DFF_349.CK  = CK;
  assign \DFF_35.CK  = CK;
  assign \DFF_350.CK  = CK;
  assign \DFF_351.CK  = CK;
  assign \DFF_352.CK  = CK;
  assign \DFF_353.CK  = CK;
  assign \DFF_354.CK  = CK;
  assign \DFF_355.CK  = CK;
  assign \DFF_356.CK  = CK;
  assign \DFF_357.CK  = CK;
  assign \DFF_358.CK  = CK;
  assign \DFF_359.CK  = CK;
  assign \DFF_36.CK  = CK;
  assign \DFF_360.CK  = CK;
  assign \DFF_361.CK  = CK;
  assign \DFF_362.CK  = CK;
  assign \DFF_363.CK  = CK;
  assign \DFF_364.CK  = CK;
  assign \DFF_365.CK  = CK;
  assign \DFF_366.CK  = CK;
  assign \DFF_367.CK  = CK;
  assign \DFF_367.D  = \DFF_99.Q ;
  assign \DFF_368.CK  = CK;
  assign \DFF_369.CK  = CK;
  assign \DFF_37.CK  = CK;
  assign \DFF_370.CK  = CK;
  assign \DFF_371.CK  = CK;
  assign \DFF_372.CK  = CK;
  assign \DFF_373.CK  = CK;
  assign \DFF_374.CK  = CK;
  assign \DFF_375.CK  = CK;
  assign \DFF_376.CK  = CK;
  assign \DFF_377.CK  = CK;
  assign \DFF_377.D  = g101;
  assign \DFF_377.Q  = \DFF_464.Q ;
  assign \DFF_378.CK  = CK;
  assign \DFF_379.CK  = CK;
  assign \DFF_38.CK  = CK;
  assign \DFF_380.CK  = CK;
  assign \DFF_381.CK  = CK;
  assign \DFF_382.CK  = CK;
  assign \DFF_383.CK  = CK;
  assign \DFF_384.CK  = CK;
  assign \DFF_385.CK  = CK;
  assign \DFF_386.CK  = CK;
  assign \DFF_387.CK  = CK;
  assign \DFF_388.CK  = CK;
  assign \DFF_389.CK  = CK;
  assign \DFF_39.CK  = CK;
  assign \DFF_390.CK  = CK;
  assign \DFF_391.CK  = CK;
  assign \DFF_392.CK  = CK;
  assign \DFF_393.CK  = CK;
  assign \DFF_394.CK  = CK;
  assign \DFF_395.CK  = CK;
  assign \DFF_396.CK  = CK;
  assign \DFF_397.CK  = CK;
  assign \DFF_398.CK  = CK;
  assign \DFF_399.CK  = CK;
  assign \DFF_4.CK  = CK;
  assign \DFF_40.CK  = CK;
  assign \DFF_400.CK  = CK;
  assign \DFF_401.CK  = CK;
  assign \DFF_402.CK  = CK;
  assign \DFF_403.CK  = CK;
  assign \DFF_404.CK  = CK;
  assign \DFF_405.CK  = CK;
  assign \DFF_405.D  = \DFF_387.Q ;
  assign \DFF_406.CK  = CK;
  assign \DFF_407.CK  = CK;
  assign \DFF_408.CK  = CK;
  assign \DFF_409.CK  = CK;
  assign \DFF_41.CK  = CK;
  assign \DFF_41.D  = \DFF_500.Q ;
  assign \DFF_410.CK  = CK;
  assign \DFF_411.CK  = CK;
  assign \DFF_411.D  = g29;
  assign \DFF_412.CK  = CK;
  assign \DFF_412.D  = \DFF_127.Q ;
  assign \DFF_413.CK  = CK;
  assign \DFF_414.CK  = CK;
  assign \DFF_415.CK  = CK;
  assign \DFF_416.CK  = CK;
  assign \DFF_417.CK  = CK;
  assign \DFF_418.CK  = CK;
  assign \DFF_419.CK  = CK;
  assign \DFF_42.CK  = CK;
  assign \DFF_420.CK  = CK;
  assign \DFF_421.CK  = CK;
  assign \DFF_422.CK  = CK;
  assign \DFF_423.CK  = CK;
  assign \DFF_424.CK  = CK;
  assign \DFF_425.CK  = CK;
  assign \DFF_426.CK  = CK;
  assign \DFF_427.CK  = CK;
  assign \DFF_428.CK  = CK;
  assign \DFF_429.CK  = CK;
  assign \DFF_43.CK  = CK;
  assign \DFF_430.CK  = CK;
  assign \DFF_431.CK  = CK;
  assign \DFF_432.CK  = CK;
  assign \DFF_433.CK  = CK;
  assign \DFF_433.D  = \DFF_393.Q ;
  assign \DFF_434.CK  = CK;
  assign \DFF_435.CK  = CK;
  assign \DFF_436.CK  = CK;
  assign \DFF_436.D  = \DFF_71.Q ;
  assign \DFF_437.CK  = CK;
  assign \DFF_438.CK  = CK;
  assign \DFF_439.CK  = CK;
  assign \DFF_44.CK  = CK;
  assign \DFF_440.CK  = CK;
  assign \DFF_441.CK  = CK;
  assign \DFF_441.D  = \DFF_357.Q ;
  assign \DFF_442.CK  = CK;
  assign \DFF_443.CK  = CK;
  assign \DFF_444.CK  = CK;
  assign \DFF_445.CK  = CK;
  assign \DFF_445.D  = \DFF_311.Q ;
  assign \DFF_446.CK  = CK;
  assign \DFF_447.CK  = CK;
  assign \DFF_448.CK  = CK;
  assign \DFF_449.CK  = CK;
  assign \DFF_45.CK  = CK;
  assign \DFF_450.CK  = CK;
  assign \DFF_451.CK  = CK;
  assign \DFF_451.D  = g28;
  assign \DFF_452.CK  = CK;
  assign \DFF_453.CK  = CK;
  assign \DFF_454.CK  = CK;
  assign \DFF_455.CK  = CK;
  assign \DFF_456.CK  = CK;
  assign \DFF_457.CK  = CK;
  assign \DFF_458.CK  = CK;
  assign \DFF_459.CK  = CK;
  assign \DFF_46.CK  = CK;
  assign \DFF_460.CK  = CK;
  assign \DFF_461.CK  = CK;
  assign \DFF_462.CK  = CK;
  assign \DFF_462.D  = g83;
  assign \DFF_463.CK  = CK;
  assign \DFF_464.CK  = CK;
  assign \DFF_464.D  = g101;
  assign \DFF_465.CK  = CK;
  assign \DFF_466.CK  = CK;
  assign \DFF_467.CK  = CK;
  assign \DFF_467.D  = \DFF_193.Q ;
  assign \DFF_468.CK  = CK;
  assign \DFF_469.CK  = CK;
  assign \DFF_47.CK  = CK;
  assign \DFF_470.CK  = CK;
  assign \DFF_471.CK  = CK;
  assign \DFF_472.CK  = CK;
  assign \DFF_473.CK  = CK;
  assign \DFF_474.CK  = CK;
  assign \DFF_475.CK  = CK;
  assign \DFF_476.CK  = CK;
  assign \DFF_476.D  = g104;
  assign \DFF_477.CK  = CK;
  assign \DFF_478.CK  = CK;
  assign \DFF_478.D  = \DFF_446.Q ;
  assign \DFF_479.CK  = CK;
  assign \DFF_48.CK  = CK;
  assign \DFF_480.CK  = CK;
  assign \DFF_481.CK  = CK;
  assign \DFF_482.CK  = CK;
  assign \DFF_483.CK  = CK;
  assign \DFF_484.CK  = CK;
  assign \DFF_485.CK  = CK;
  assign \DFF_486.CK  = CK;
  assign \DFF_487.CK  = CK;
  assign \DFF_488.CK  = CK;
  assign \DFF_489.CK  = CK;
  assign \DFF_49.CK  = CK;
  assign \DFF_490.CK  = CK;
  assign \DFF_491.CK  = CK;
  assign \DFF_492.CK  = CK;
  assign \DFF_493.CK  = CK;
  assign \DFF_494.CK  = CK;
  assign \DFF_495.CK  = CK;
  assign \DFF_496.CK  = CK;
  assign \DFF_497.CK  = CK;
  assign \DFF_498.CK  = CK;
  assign \DFF_499.CK  = CK;
  assign \DFF_5.CK  = CK;
  assign \DFF_50.CK  = CK;
  assign \DFF_500.CK  = CK;
  assign \DFF_501.CK  = CK;
  assign \DFF_502.CK  = CK;
  assign \DFF_502.D  = g102;
  assign \DFF_503.CK  = CK;
  assign \DFF_504.CK  = CK;
  assign \DFF_505.CK  = CK;
  assign \DFF_506.CK  = CK;
  assign \DFF_507.CK  = CK;
  assign \DFF_508.CK  = CK;
  assign \DFF_509.CK  = CK;
  assign \DFF_51.CK  = CK;
  assign \DFF_510.CK  = CK;
  assign \DFF_511.CK  = CK;
  assign \DFF_512.CK  = CK;
  assign \DFF_513.CK  = CK;
  assign \DFF_514.CK  = CK;
  assign \DFF_515.CK  = CK;
  assign \DFF_516.CK  = CK;
  assign \DFF_517.CK  = CK;
  assign \DFF_518.CK  = CK;
  assign \DFF_519.CK  = CK;
  assign \DFF_52.CK  = CK;
  assign \DFF_520.CK  = CK;
  assign \DFF_521.CK  = CK;
  assign \DFF_522.CK  = CK;
  assign \DFF_523.CK  = CK;
  assign \DFF_524.CK  = CK;
  assign \DFF_525.CK  = CK;
  assign \DFF_526.CK  = CK;
  assign \DFF_527.CK  = CK;
  assign \DFF_528.CK  = CK;
  assign \DFF_529.CK  = CK;
  assign \DFF_53.CK  = CK;
  assign \DFF_530.CK  = CK;
  assign \DFF_531.CK  = CK;
  assign \DFF_532.CK  = CK;
  assign \DFF_533.CK  = CK;
  assign \DFF_54.CK  = CK;
  assign \DFF_54.D  = \DFF_174.Q ;
  assign \DFF_55.CK  = CK;
  assign \DFF_55.D  = \DFF_227.Q ;
  assign \DFF_56.CK  = CK;
  assign \DFF_57.CK  = CK;
  assign \DFF_58.CK  = CK;
  assign \DFF_59.CK  = CK;
  assign \DFF_6.CK  = CK;
  assign \DFF_60.CK  = CK;
  assign \DFF_61.CK  = CK;
  assign \DFF_62.CK  = CK;
  assign \DFF_62.D  = g104;
  assign \DFF_62.Q  = \DFF_476.Q ;
  assign \DFF_63.CK  = CK;
  assign \DFF_64.CK  = CK;
  assign \DFF_65.CK  = CK;
  assign \DFF_65.D  = \DFF_443.Q ;
  assign \DFF_66.CK  = CK;
  assign \DFF_67.CK  = CK;
  assign \DFF_68.CK  = CK;
  assign \DFF_68.D  = \DFF_462.Q ;
  assign \DFF_68.Q  = \DFF_156.Q ;
  assign \DFF_69.CK  = CK;
  assign \DFF_7.CK  = CK;
  assign \DFF_70.CK  = CK;
  assign \DFF_71.CK  = CK;
  assign \DFF_72.CK  = CK;
  assign \DFF_73.CK  = CK;
  assign \DFF_74.CK  = CK;
  assign \DFF_75.CK  = CK;
  assign \DFF_76.CK  = CK;
  assign \DFF_77.CK  = CK;
  assign \DFF_78.CK  = CK;
  assign \DFF_79.CK  = CK;
  assign \DFF_8.CK  = CK;
  assign \DFF_80.CK  = CK;
  assign \DFF_80.D  = \DFF_156.Q ;
  assign \DFF_80.Q  = \DFF_304.Q ;
  assign \DFF_81.CK  = CK;
  assign \DFF_82.CK  = CK;
  assign \DFF_83.CK  = CK;
  assign \DFF_84.CK  = CK;
  assign \DFF_85.CK  = CK;
  assign \DFF_86.CK  = CK;
  assign \DFF_87.CK  = CK;
  assign \DFF_88.CK  = CK;
  assign \DFF_89.CK  = CK;
  assign \DFF_89.D  = \DFF_304.Q ;
  assign \DFF_9.CK  = CK;
  assign \DFF_90.CK  = CK;
  assign \DFF_91.CK  = CK;
  assign \DFF_92.CK  = CK;
  assign \DFF_93.CK  = CK;
  assign \DFF_93.D  = \DFF_53.Q ;
  assign \DFF_94.CK  = CK;
  assign \DFF_95.CK  = CK;
  assign \DFF_96.CK  = CK;
  assign \DFF_97.CK  = CK;
  assign \DFF_98.CK  = CK;
  assign \DFF_99.CK  = CK;
  assign I10015 = g27;
  assign I10698 = g82;
  assign I11397 = g82;
  assign I11989 = \DFF_233.Q ;
  assign I12655 = g41;
  assign I12690 = \DFF_233.Q ;
  assign I13117 = \DFF_233.Q ;
  assign I13185 = \DFF_233.Q ;
  assign I16387 = g11206;
  assign I5254 = \DFF_275.D ;
  assign I5336 = \DFF_275.D ;
  assign I5801 = \DFF_112.Q ;
  assign I5815 = \DFF_227.Q ;
  assign I5827 = g877;
  assign I5830 = \DFF_335.Q ;
  assign I5847 = \DFF_37.Q ;
  assign I5850 = g881;
  assign I5913 = g42;
  assign I5922 = g30;
  assign I5926 = g43;
  assign I5935 = g31;
  assign I5940 = g44;
  assign I5946 = g82;
  assign I5952 = \DFF_360.Q ;
  assign I5957 = g45;
  assign I5963 = g89;
  assign I5970 = g46;
  assign I5976 = g90;
  assign I5986 = g47;
  assign I5992 = g83;
  assign I5995 = g91;
  assign I5998 = g101;
  assign I6007 = g48;
  assign I6013 = g92;
  assign I6016 = g102;
  assign I6028 = g84;
  assign I6031 = g93;
  assign I6034 = g103;
  assign I6040 = g41;
  assign I6046 = g85;
  assign I6049 = g94;
  assign I6052 = g104;
  assign I6061 = \DFF_233.Q ;
  assign I6065 = g86;
  assign I6068 = g95;
  assign I6074 = g28;
  assign I6085 = g87;
  assign I6088 = g96;
  assign I6102 = g88;
  assign I6118 = g99;
  assign I6133 = g100;
  assign I6163 = g23;
  assign I6217 = g29;
  assign I6233 = \DFF_77.Q ;
  assign I6260 = g1696;
  assign I6264 = \DFF_311.Q ;
  assign I6343 = g109;
  assign I6360 = \DFF_174.Q ;
  assign I6367 = \DFF_420.Q ;
  assign I6373 = \DFF_113.Q ;
  assign I6461 = \DFF_174.Q ;
  assign I6474 = \DFF_269.Q ;
  assign I6498 = g23;
  assign I6507 = \DFF_384.Q ;
  assign I6513 = \DFF_242.Q ;
  assign I6520 = \DFF_113.Q ;
  assign I6523 = \DFF_228.Q ;
  assign I6531 = \DFF_113.Q ;
  assign I6535 = \DFF_92.Q ;
  assign I6538 = \DFF_350.Q ;
  assign I6543 = \DFF_113.Q ;
  assign I6549 = \DFF_116.Q ;
  assign I6553 = \DFF_113.Q ;
  assign I6560 = \DFF_22.Q ;
  assign I6569 = \DFF_113.Q ;
  assign I6572 = \DFF_319.Q ;
  assign I6580 = \DFF_113.Q ;
  assign I6590 = \DFF_113.Q ;
  assign I6601 = \DFF_113.Q ;
  assign I6616 = \DFF_113.Q ;
  assign I6679 = \DFF_233.Q ;
  assign I6690 = \DFF_112.Q ;
  assign I6694 = \DFF_227.Q ;
  assign I6738 = g109;
  assign I6812 = \DFF_174.Q ;
  assign I6856 = g1700;
  assign I6894 = g42;
  assign I6901 = g30;
  assign I6904 = g43;
  assign I6911 = g31;
  assign I6914 = g44;
  assign I6917 = g82;
  assign I6921 = g45;
  assign I6924 = g89;
  assign I6929 = g46;
  assign I6932 = g90;
  assign I6938 = g47;
  assign I6941 = g83;
  assign I6944 = g91;
  assign I6947 = g101;
  assign I6952 = g48;
  assign I6955 = g92;
  assign I6958 = g102;
  assign I6965 = g84;
  assign I6968 = g93;
  assign I6971 = g103;
  assign I6976 = g41;
  assign I6979 = g85;
  assign I6982 = g94;
  assign I6985 = g104;
  assign I6996 = g86;
  assign I6999 = g95;
  assign I7002 = g28;
  assign I7006 = g87;
  assign I7009 = g96;
  assign I7014 = g88;
  assign I7022 = g99;
  assign I7029 = g100;
  assign I7061 = g1696;
  assign I7076 = g29;
  assign I7086 = \DFF_174.Q ;
  assign I7096 = \DFF_113.Q ;
  assign I7104 = \DFF_113.Q ;
  assign I7112 = \DFF_113.Q ;
  assign I7311 = \DFF_168.Q ;
  assign I7468 = g1700;
  assign I7478 = g109;
  assign I7509 = g109;
  assign I7625 = \DFF_168.Q ;
  assign I7633 = \DFF_233.Q ;
  assign I7636 = \DFF_384.Q ;
  assign I7639 = g42;
  assign I7648 = g30;
  assign I7651 = \DFF_242.Q ;
  assign I7654 = g43;
  assign I7659 = g31;
  assign I7662 = \DFF_228.Q ;
  assign I7665 = g44;
  assign I7668 = g82;
  assign I7671 = \DFF_92.Q ;
  assign I7674 = \DFF_350.Q ;
  assign I7677 = g45;
  assign I7680 = g89;
  assign I7691 = \DFF_116.Q ;
  assign I7694 = g46;
  assign I7697 = g90;
  assign I7707 = \DFF_22.Q ;
  assign I7710 = g47;
  assign I7713 = g83;
  assign I7716 = g91;
  assign I7719 = g101;
  assign I7726 = \DFF_319.Q ;
  assign I7729 = g48;
  assign I7732 = g92;
  assign I7735 = g102;
  assign I7743 = g84;
  assign I7746 = g93;
  assign I7749 = g103;
  assign I7757 = g41;
  assign I7760 = g85;
  assign I7763 = g94;
  assign I7766 = g104;
  assign I7776 = g86;
  assign I7779 = g95;
  assign I7782 = g28;
  assign I7790 = g87;
  assign I7793 = g96;
  assign I7800 = g88;
  assign I7810 = g99;
  assign I7820 = g100;
  assign I7906 = g29;
  assign I8031 = g109;
  assign I8164 = g109;
  assign I8192 = g109;
  assign I8211 = g109;
  assign I8231 = g27;
  assign I8311 = g109;
  assign I8324 = g109;
  assign I8337 = \DFF_233.Q ;
  assign I8351 = g109;
  assign I8358 = g109;
  assign I8418 = g109;
  assign I9040 = g109;
  assign I9084 = g27;
  assign I9424 = \DFF_233.Q ;
  assign I9427 = \DFF_233.Q ;
  assign g1 = \DFF_528.Q ;
  assign g1003 = \DFF_414.Q ;
  assign g1007 = \DFF_108.Q ;
  assign g1011 = \DFF_167.Q ;
  assign g1015 = \DFF_115.Q ;
  assign g1019 = \DFF_87.Q ;
  assign g1023 = \DFF_192.Q ;
  assign g1027 = \DFF_413.Q ;
  assign g1032 = \DFF_234.Q ;
  assign g10336 = g10377;
  assign g10339 = g10379;
  assign g1035 = \DFF_274.Q ;
  assign g10378 = g10377;
  assign g1038 = \DFF_298.Q ;
  assign g10380 = g10379;
  assign g10402 = g10455;
  assign g10405 = g10457;
  assign g10408 = g10459;
  assign g1041 = \DFF_160.Q ;
  assign g10411 = g10461;
  assign g10414 = g10463;
  assign g10417 = g10465;
  assign g1044 = \DFF_35.Q ;
  assign g10456 = g10455;
  assign g10458 = g10457;
  assign g10460 = g10459;
  assign g10462 = g10461;
  assign g10464 = g10463;
  assign g10466 = g10465;
  assign g1047 = \DFF_422.Q ;
  assign g105 = \DFF_161.Q ;
  assign g1050 = \DFF_527.Q ;
  assign g10515 = g10628;
  assign g1053 = \DFF_236.Q ;
  assign g10531 = g10377;
  assign g10532 = g10379;
  assign g1056 = \DFF_439.Q ;
  assign g10575 = g10455;
  assign g10576 = g10457;
  assign g10577 = g10459;
  assign g10578 = g10461;
  assign g10579 = g10463;
  assign g10580 = g10465;
  assign g10583 = g11206;
  assign g10589 = g10628;
  assign g1059 = \DFF_110.Q ;
  assign g1062 = \DFF_305.Q ;
  assign g1065 = \DFF_348.Q ;
  assign g10663 = \DFF_22.D ;
  assign g10664 = \DFF_319.D ;
  assign g1068 = \DFF_376.Q ;
  assign g10707 = \DFF_96.D ;
  assign g1071 = \DFF_292.Q ;
  assign g10711 = \DFF_321.D ;
  assign g10712 = g10801;
  assign g10717 = \DFF_524.D ;
  assign g10718 = \DFF_166.D ;
  assign g10719 = \DFF_168.D ;
  assign g10720 = \DFF_384.D ;
  assign g10721 = \DFF_242.D ;
  assign g10722 = \DFF_228.D ;
  assign g10724 = \DFF_350.D ;
  assign g10726 = \DFF_116.D ;
  assign g10734 = \DFF_22.D ;
  assign g10735 = \DFF_319.D ;
  assign g1074 = \DFF_170.Q ;
  assign g10765 = \DFF_423.D ;
  assign g10767 = \DFF_285.D ;
  assign g1077 = \DFF_27.Q ;
  assign g10770 = \DFF_120.D ;
  assign g10771 = \DFF_530.D ;
  assign g10773 = \DFF_370.D ;
  assign g10774 = \DFF_22.D ;
  assign g10775 = \DFF_319.D ;
  assign g10776 = \DFF_465.D ;
  assign g10779 = g11163;
  assign g10780 = \DFF_507.D ;
  assign g10781 = \DFF_423.D ;
  assign g10782 = \DFF_23.D ;
  assign g10783 = \DFF_285.D ;
  assign g10784 = \DFF_421.D ;
  assign g10785 = \DFF_472.D ;
  assign g10786 = \DFF_120.D ;
  assign g10787 = \DFF_530.D ;
  assign g10788 = \DFF_37.D ;
  assign g10791 = \DFF_460.D ;
  assign g10792 = \DFF_370.D ;
  assign g10793 = \DFF_50.D ;
  assign g10794 = \DFF_96.D ;
  assign g10795 = \DFF_186.D ;
  assign g10796 = \DFF_321.D ;
  assign g10797 = \DFF_260.D ;
  assign g10798 = \DFF_208.D ;
  assign g10799 = \DFF_288.D ;
  assign g108 = \DFF_335.Q ;
  assign g1080 = \DFF_173.Q ;
  assign g10800 = \DFF_211.D ;
  assign g10802 = g10801;
  assign g10803 = g11206;
  assign g10804 = \DFF_524.D ;
  assign g10806 = \DFF_166.D ;
  assign g10819 = \DFF_168.D ;
  assign g10821 = \DFF_384.D ;
  assign g10825 = \DFF_242.D ;
  assign g10826 = \DFF_228.D ;
  assign g1083 = \DFF_402.Q ;
  assign g10848 = \DFF_350.D ;
  assign g10850 = \DFF_116.D ;
  assign g10854 = g11206;
  assign g10855 = \DFF_159.D ;
  assign g10858 = \DFF_26.D ;
  assign g10859 = \DFF_45.D ;
  assign g1086 = \DFF_94.Q ;
  assign g10860 = \DFF_69.D ;
  assign g10861 = \DFF_280.D ;
  assign g10862 = \DFF_101.D ;
  assign g10863 = \DFF_504.D ;
  assign g10864 = \DFF_206.D ;
  assign g10865 = \DFF_162.D ;
  assign g10866 = \DFF_73.D ;
  assign g10867 = \DFF_168.D ;
  assign g10868 = \DFF_384.D ;
  assign g10869 = \DFF_242.D ;
  assign g10870 = \DFF_228.D ;
  assign g10871 = \DFF_350.D ;
  assign g10872 = \DFF_116.D ;
  assign g10874 = \DFF_423.D ;
  assign g10875 = \DFF_285.D ;
  assign g10876 = \DFF_524.D ;
  assign g10877 = \DFF_166.D ;
  assign g10878 = \DFF_120.D ;
  assign g10879 = \DFF_530.D ;
  assign g10880 = \DFF_370.D ;
  assign g10881 = \DFF_96.D ;
  assign g10882 = \DFF_321.D ;
  assign g10887 = \DFF_26.D ;
  assign g10888 = \DFF_45.D ;
  assign g10889 = \DFF_69.D ;
  assign g1089 = \DFF_290.Q ;
  assign g10890 = \DFF_280.D ;
  assign g10891 = \DFF_101.D ;
  assign g10892 = \DFF_504.D ;
  assign g10893 = \DFF_206.D ;
  assign g10894 = \DFF_162.D ;
  assign g10895 = \DFF_73.D ;
  assign g10896 = \DFF_465.D ;
  assign g10898 = \DFF_161.D ;
  assign g10900 = \DFF_460.D ;
  assign g10902 = \DFF_50.D ;
  assign g10904 = \DFF_186.D ;
  assign g10905 = \DFF_507.D ;
  assign g10906 = \DFF_260.D ;
  assign g10907 = \DFF_23.D ;
  assign g10908 = \DFF_208.D ;
  assign g10909 = \DFF_421.D ;
  assign g10910 = \DFF_288.D ;
  assign g10911 = \DFF_472.D ;
  assign g10912 = \DFF_211.D ;
  assign g10913 = \DFF_37.D ;
  assign g1092 = \DFF_16.Q ;
  assign g10936 = \DFF_420.D ;
  assign g1095 = \DFF_56.Q ;
  assign g10972 = g11163;
  assign g10973 = g11206;
  assign g1098 = \DFF_82.Q ;
  assign g110 = g109;
  assign g1101 = \DFF_158.Q ;
  assign g11014 = \DFF_159.D ;
  assign g11033 = \DFF_45.D ;
  assign g11034 = \DFF_280.D ;
  assign g11035 = \DFF_504.D ;
  assign g11036 = \DFF_162.D ;
  assign g11037 = \DFF_26.D ;
  assign g11038 = \DFF_69.D ;
  assign g11039 = \DFF_101.D ;
  assign g1104 = \DFF_31.Q ;
  assign g11040 = \DFF_206.D ;
  assign g11041 = \DFF_73.D ;
  assign g11042 = \DFF_465.D ;
  assign g11043 = \DFF_460.D ;
  assign g11044 = \DFF_159.D ;
  assign g11047 = \DFF_50.D ;
  assign g11048 = \DFF_186.D ;
  assign g11049 = \DFF_260.D ;
  assign g11050 = \DFF_208.D ;
  assign g11051 = \DFF_288.D ;
  assign g11052 = \DFF_211.D ;
  assign g1107 = \DFF_417.Q ;
  assign g11074 = g10801;
  assign g11076 = \DFF_161.D ;
  assign g11079 = \DFF_507.D ;
  assign g11080 = \DFF_23.D ;
  assign g11081 = \DFF_421.D ;
  assign g11082 = \DFF_472.D ;
  assign g11084 = g11163;
  assign g11086 = \DFF_37.D ;
  assign g11088 = g11206;
  assign g11096 = \DFF_420.D ;
  assign g1110 = \DFF_278.Q ;
  assign g1113 = \DFF_517.Q ;
  assign g1117 = \DFF_214.Q ;
  assign g11179 = \DFF_37.D ;
  assign g11180 = \DFF_161.D ;
  assign g11181 = \DFF_507.D ;
  assign g11182 = \DFF_23.D ;
  assign g11183 = \DFF_421.D ;
  assign g11184 = \DFF_472.D ;
  assign g11185 = \DFF_420.D ;
  assign g11207 = g11206;
  assign g1121 = \DFF_457.Q ;
  assign g1125 = \DFF_399.Q ;
  assign g11256 = \DFF_124.D ;
  assign g11257 = \DFF_3.D ;
  assign g11258 = \DFF_368.D ;
  assign g11259 = \DFF_171.D ;
  assign g11260 = \DFF_378.D ;
  assign g11261 = \DFF_512.D ;
  assign g11262 = \DFF_492.D ;
  assign g11263 = \DFF_217.D ;
  assign g11264 = \DFF_394.D ;
  assign g11265 = \DFF_114.D ;
  assign g11266 = \DFF_177.D ;
  assign g11267 = \DFF_419.D ;
  assign g11268 = \DFF_491.D ;
  assign g11269 = \DFF_204.D ;
  assign g11270 = \DFF_406.D ;
  assign g11286 = \DFF_92.D ;
  assign g1129 = \DFF_366.Q ;
  assign g11290 = \DFF_207.D ;
  assign g11291 = \DFF_409.D ;
  assign g11292 = \DFF_483.D ;
  assign g11293 = \DFF_311.D ;
  assign g11294 = \DFF_178.D ;
  assign g11298 = \DFF_312.D ;
  assign g113 = \DFF_71.Q ;
  assign g11300 = \DFF_454.D ;
  assign g11303 = \DFF_365.D ;
  assign g11305 = \DFF_317.D ;
  assign g11306 = \DFF_408.D ;
  assign g11308 = \DFF_106.D ;
  assign g11310 = \DFF_148.D ;
  assign g11312 = \DFF_181.D ;
  assign g11314 = \DFF_351.D ;
  assign g11320 = \DFF_19.D ;
  assign g11324 = \DFF_430.D ;
  assign g11325 = \DFF_205.D ;
  assign g11326 = \DFF_203.D ;
  assign g11327 = \DFF_522.D ;
  assign g11328 = \DFF_210.D ;
  assign g11329 = \DFF_475.D ;
  assign g1133 = \DFF_145.Q ;
  assign g11330 = \DFF_447.D ;
  assign g11331 = \DFF_151.D ;
  assign g11332 = \DFF_329.D ;
  assign g11333 = \DFF_51.D ;
  assign g11334 = \DFF_221.D ;
  assign g11335 = \DFF_459.D ;
  assign g11336 = \DFF_529.D ;
  assign g11337 = \DFF_245.D ;
  assign g11338 = \DFF_379.D ;
  assign g11340 = \DFF_264.D ;
  assign g11341 = \DFF_317.D ;
  assign g11342 = \DFF_408.D ;
  assign g11343 = \DFF_106.D ;
  assign g11344 = \DFF_148.D ;
  assign g11345 = \DFF_181.D ;
  assign g11346 = \DFF_351.D ;
  assign g11347 = \DFF_19.D ;
  assign g11349 = \DFF_294.D ;
  assign g11350 = g11206;
  assign g11351 = \DFF_178.D ;
  assign g11352 = \DFF_311.D ;
  assign g11353 = \DFF_92.D ;
  assign g1137 = \DFF_353.Q ;
  assign g11372 = \DFF_12.D ;
  assign g11376 = \DFF_255.D ;
  assign g11380 = \DFF_152.D ;
  assign g11388 = \DFF_207.D ;
  assign g11389 = \DFF_409.D ;
  assign g11390 = \DFF_483.D ;
  assign g11391 = \DFF_14.D ;
  assign g11392 = \DFF_52.D ;
  assign g11393 = \DFF_293.D ;
  assign g11394 = \DFF_312.D ;
  assign g11395 = \DFF_454.D ;
  assign g11396 = \DFF_365.D ;
  assign g11397 = \DFF_92.D ;
  assign g11398 = \DFF_312.D ;
  assign g11399 = \DFF_454.D ;
  assign g114 = \DFF_436.Q ;
  assign g11400 = \DFF_365.D ;
  assign g11401 = \DFF_317.D ;
  assign g11402 = \DFF_408.D ;
  assign g11403 = \DFF_106.D ;
  assign g11404 = \DFF_148.D ;
  assign g11405 = \DFF_181.D ;
  assign g11406 = \DFF_351.D ;
  assign g11408 = \DFF_311.D ;
  assign g11409 = \DFF_178.D ;
  assign g1141 = \DFF_468.Q ;
  assign g11410 = \DFF_207.D ;
  assign g11411 = \DFF_409.D ;
  assign g11412 = \DFF_483.D ;
  assign g11417 = \DFF_14.D ;
  assign g11419 = \DFF_52.D ;
  assign g11420 = \DFF_293.D ;
  assign g11421 = \DFF_264.D ;
  assign g11423 = \DFF_19.D ;
  assign g11424 = \DFF_294.D ;
  assign g11436 = \DFF_12.D ;
  assign g11437 = \DFF_255.D ;
  assign g11438 = \DFF_152.D ;
  assign g11439 = \DFF_19.D ;
  assign g11440 = \DFF_207.D ;
  assign g11441 = \DFF_409.D ;
  assign g11442 = \DFF_483.D ;
  assign g11443 = \DFF_480.D ;
  assign g11444 = \DFF_12.D ;
  assign g11445 = \DFF_255.D ;
  assign g11446 = \DFF_152.D ;
  assign g1145 = \DFF_416.Q ;
  assign g11450 = \DFF_14.D ;
  assign g11451 = \DFF_52.D ;
  assign g11453 = \DFF_293.D ;
  assign g11454 = \DFF_264.D ;
  assign g11457 = \DFF_294.D ;
  assign g11466 = \DFF_264.D ;
  assign g11467 = \DFF_12.D ;
  assign g11468 = \DFF_255.D ;
  assign g11469 = \DFF_152.D ;
  assign g11470 = \DFF_294.D ;
  assign g11471 = \DFF_14.D ;
  assign g11472 = \DFF_52.D ;
  assign g11473 = \DFF_293.D ;
  assign g11478 = \DFF_499.D ;
  assign g11481 = \DFF_440.D ;
  assign g11482 = \DFF_79.D ;
  assign g11483 = \DFF_70.D ;
  assign g11484 = \DFF_216.D ;
  assign g11485 = \DFF_283.D ;
  assign g11486 = \DFF_238.D ;
  assign g11487 = \DFF_308.D ;
  assign g11488 = \DFF_230.D ;
  assign g11489 = 1'b0;
  assign g1149 = \DFF_383.Q ;
  assign g11495 = \DFF_499.D ;
  assign g11497 = \DFF_440.D ;
  assign g11498 = \DFF_79.D ;
  assign g11499 = \DFF_70.D ;
  assign g115 = \DFF_473.Q ;
  assign g11500 = \DFF_216.D ;
  assign g11501 = \DFF_283.D ;
  assign g11502 = \DFF_238.D ;
  assign g11503 = \DFF_308.D ;
  assign g11504 = \DFF_230.D ;
  assign g11505 = \DFF_499.D ;
  assign g11506 = \DFF_440.D ;
  assign g11507 = \DFF_79.D ;
  assign g11508 = \DFF_70.D ;
  assign g11509 = \DFF_216.D ;
  assign g11510 = \DFF_283.D ;
  assign g11511 = \DFF_238.D ;
  assign g11512 = \DFF_308.D ;
  assign g11513 = \DFF_230.D ;
  assign g11514 = \DFF_143.D ;
  assign g1153 = \DFF_7.Q ;
  assign g11550 = \DFF_143.D ;
  assign g11561 = \DFF_335.D ;
  assign g1157 = \DFF_240.Q ;
  assign g11577 = \DFF_143.D ;
  assign g11578 = \DFF_335.D ;
  assign g11579 = \DFF_509.D ;
  assign g11593 = \DFF_335.D ;
  assign g11594 = \DFF_143.D ;
  assign g11598 = \DFF_509.D ;
  assign g1160 = \DFF_525.Q ;
  assign g11602 = \DFF_134.D ;
  assign g11603 = \DFF_481.D ;
  assign g11604 = \DFF_342.D ;
  assign g11605 = \DFF_448.D ;
  assign g11606 = \DFF_458.D ;
  assign g11607 = \DFF_325.D ;
  assign g11608 = \DFF_195.D ;
  assign g11609 = \DFF_432.D ;
  assign g11610 = \DFF_146.D ;
  assign g11611 = \DFF_509.D ;
  assign g11614 = \DFF_134.D ;
  assign g11616 = \DFF_481.D ;
  assign g11617 = \DFF_342.D ;
  assign g11618 = \DFF_448.D ;
  assign g11619 = \DFF_458.D ;
  assign g11620 = \DFF_325.D ;
  assign g11621 = \DFF_195.D ;
  assign g11622 = \DFF_432.D ;
  assign g11623 = \DFF_146.D ;
  assign g11625 = \DFF_266.D ;
  assign g11627 = \DFF_134.D ;
  assign g11628 = \DFF_481.D ;
  assign g11629 = \DFF_342.D ;
  assign g1163 = \DFF_232.Q ;
  assign g11630 = \DFF_448.D ;
  assign g11631 = \DFF_458.D ;
  assign g11632 = \DFF_325.D ;
  assign g11633 = \DFF_195.D ;
  assign g11634 = \DFF_432.D ;
  assign g11635 = \DFF_146.D ;
  assign g11636 = \DFF_344.D ;
  assign g11638 = \DFF_266.D ;
  assign g11639 = \DFF_470.D ;
  assign g11640 = \DFF_198.D ;
  assign g11641 = \DFF_506.D ;
  assign g11642 = \DFF_266.D ;
  assign g11643 = \DFF_470.D ;
  assign g11644 = \DFF_198.D ;
  assign g11645 = \DFF_506.D ;
  assign g11646 = \DFF_344.D ;
  assign g11647 = \DFF_263.D ;
  assign g11648 = \DFF_470.D ;
  assign g11649 = \DFF_198.D ;
  assign g11650 = \DFF_506.D ;
  assign g11651 = \DFF_344.D ;
  assign g11652 = \DFF_263.D ;
  assign g11653 = \DFF_263.D ;
  assign g11654 = \DFF_344.D ;
  assign g11655 = \DFF_470.D ;
  assign g11656 = \DFF_198.D ;
  assign g11657 = \DFF_506.D ;
  assign g1166 = \DFF_438.Q ;
  assign g119 = \DFF_380.Q ;
  assign g12 = \DFF_531.Q ;
  assign g1206 = \DFF_328.Q ;
  assign g1212 = \DFF_299.Q ;
  assign g1216 = \DFF_126.Q ;
  assign g1217 = \DFF_137.Q ;
  assign g1218 = \DFF_361.Q ;
  assign g1223 = \DFF_418.Q ;
  assign g1227 = \DFF_119.Q ;
  assign g123 = \DFF_4.Q ;
  assign g1231 = \DFF_28.Q ;
  assign g1235 = \DFF_510.Q ;
  assign g1240 = \DFF_202.Q ;
  assign g1245 = \DFF_334.Q ;
  assign g1250 = \DFF_231.Q ;
  assign g1255 = \DFF_355.Q ;
  assign g1260 = \DFF_442.Q ;
  assign g1265 = \DFF_58.Q ;
  assign g127 = \DFF_508.Q ;
  assign g1270 = \DFF_322.Q ;
  assign g1275 = \DFF_480.Q ;
  assign g1280 = \DFF_401.Q ;
  assign g1284 = \DFF_486.Q ;
  assign g1289 = \DFF_0.Q ;
  assign g1292 = \DFF_250.Q ;
  assign g1296 = \DFF_61.Q ;
  assign g1300 = \DFF_498.Q ;
  assign g1304 = \DFF_32.Q ;
  assign g1308 = \DFF_134.Q ;
  assign g131 = \DFF_444.Q ;
  assign g1311 = \DFF_481.Q ;
  assign g1314 = \DFF_342.Q ;
  assign g1317 = \DFF_215.Q ;
  assign g1318 = \DFF_448.Q ;
  assign g1321 = \DFF_458.Q ;
  assign g1324 = \DFF_325.Q ;
  assign g1327 = \DFF_195.Q ;
  assign g1330 = \DFF_432.Q ;
  assign g1333 = \DFF_146.Q ;
  assign g1336 = \DFF_344.Q ;
  assign g1341 = \DFF_470.Q ;
  assign g1346 = \DFF_198.Q ;
  assign g135 = \DFF_474.Q ;
  assign g1351 = \DFF_506.Q ;
  assign g1356 = \DFF_226.Q ;
  assign g1357 = \DFF_241.Q ;
  assign g1360 = \DFF_526.Q ;
  assign g1361 = \DFF_194.Q ;
  assign g1362 = \DFF_88.Q ;
  assign g1365 = \DFF_142.Q ;
  assign g1368 = \DFF_163.Q ;
  assign g1371 = \DFF_67.Q ;
  assign g1374 = \DFF_484.Q ;
  assign g1377 = \DFF_327.Q ;
  assign g1380 = \DFF_487.Q ;
  assign g1383 = \DFF_189.Q ;
  assign g1386 = \DFF_396.Q ;
  assign g1389 = \DFF_66.Q ;
  assign g139 = \DFF_382.Q ;
  assign g1393 = \DFF_452.Q ;
  assign g1394 = \DFF_289.Q ;
  assign g1397 = \DFF_153.Q ;
  assign g1400 = \DFF_182.Q ;
  assign g1403 = \DFF_415.Q ;
  assign g1407 = \DFF_109.Q ;
  assign g1411 = \DFF_169.Q ;
  assign g1415 = \DFF_118.Q ;
  assign g1419 = \DFF_90.Q ;
  assign g1424 = \DFF_24.Q ;
  assign g1428 = \DFF_128.Q ;
  assign g143 = \DFF_296.Q ;
  assign g1432 = \DFF_235.Q ;
  assign g1436 = \DFF_47.Q ;
  assign g1440 = \DFF_503.Q ;
  assign g1444 = \DFF_36.Q ;
  assign g1448 = \DFF_143.Q ;
  assign g1453 = \DFF_237.Q ;
  assign g1458 = \DFF_165.Q ;
  assign g1462 = \DFF_306.Q ;
  assign g1466 = \DFF_139.Q ;
  assign g1470 = \DFF_98.Q ;
  assign g1474 = \DFF_172.Q ;
  assign g1478 = \DFF_273.Q ;
  assign g148 = \DFF_337.Q ;
  assign g1482 = \DFF_277.Q ;
  assign g1486 = \DFF_95.Q ;
  assign g1490 = \DFF_437.Q ;
  assign g1494 = \DFF_519.Q ;
  assign g1499 = \DFF_34.Q ;
  assign g1504 = \DFF_97.Q ;
  assign g1508 = \DFF_201.Q ;
  assign g1512 = \DFF_435.Q ;
  assign g1515 = \DFF_494.Q ;
  assign g1520 = \DFF_315.Q ;
  assign g1524 = \DFF_391.Q ;
  assign g1528 = \DFF_505.Q ;
  assign g153 = \DFF_147.Q ;
  assign g1531 = \DFF_164.Q ;
  assign g1534 = \DFF_42.Q ;
  assign g1537 = \DFF_426.Q ;
  assign g1540 = \DFF_326.Q ;
  assign g1543 = \DFF_39.Q ;
  assign g1546 = \DFF_258.Q ;
  assign g1549 = \DFF_453.Q ;
  assign g1552 = \DFF_463.Q ;
  assign g1555 = \DFF_514.Q ;
  assign g1558 = \DFF_10.Q ;
  assign g1561 = \DFF_256.Q ;
  assign g1564 = \DFF_130.Q ;
  assign g1567 = \DFF_520.Q ;
  assign g1571 = \DFF_140.Q ;
  assign g1574 = \DFF_17.Q ;
  assign g1577 = \DFF_392.Q ;
  assign g158 = \DFF_190.Q ;
  assign g1580 = \DFF_20.Q ;
  assign g1583 = \DFF_254.Q ;
  assign g1586 = \DFF_466.Q ;
  assign g1589 = \DFF_138.Q ;
  assign g1592 = \DFF_371.Q ;
  assign g1595 = \DFF_425.Q ;
  assign g1598 = \DFF_456.Q ;
  assign g16 = \DFF_122.Q ;
  assign g1601 = \DFF_218.Q ;
  assign g1604 = \DFF_81.Q ;
  assign g1607 = \DFF_477.Q ;
  assign g1610 = \DFF_323.Q ;
  assign g1615 = \DFF_482.Q ;
  assign g1618 = \DFF_509.Q ;
  assign g162 = \DFF_490.Q ;
  assign g1621 = \DFF_516.Q ;
  assign g1624 = \DFF_374.Q ;
  assign g1627 = \DFF_249.Q ;
  assign g1630 = \DFF_495.Q ;
  assign g1633 = \DFF_199.Q ;
  assign g1636 = \DFF_404.Q ;
  assign g1639 = \DFF_74.Q ;
  assign g1642 = \DFF_421.Q ;
  assign g1645 = \DFF_472.Q ;
  assign g1648 = \DFF_507.Q ;
  assign g1651 = \DFF_23.Q ;
  assign g1654 = \DFF_423.Q ;
  assign g1657 = \DFF_285.Q ;
  assign g166 = \DFF_220.Q ;
  assign g1660 = \DFF_45.Q ;
  assign g1663 = \DFF_280.Q ;
  assign g1666 = \DFF_504.Q ;
  assign g1669 = \DFF_162.Q ;
  assign g1672 = \DFF_26.Q ;
  assign g1675 = \DFF_69.Q ;
  assign g1678 = \DFF_101.Q ;
  assign g1681 = \DFF_206.Q ;
  assign g1684 = \DFF_73.Q ;
  assign g1687 = \DFF_465.Q ;
  assign g1690 = \DFF_276.Q ;
  assign g17 = \DFF_262.Q ;
  assign g170 = \DFF_314.Q ;
  assign g1703 = \DFF_372.Q ;
  assign g1707 = \DFF_77.Q ;
  assign g1710 = \DFF_471.Q ;
  assign g1713 = \DFF_174.Q ;
  assign g1718 = \DFF_113.Q ;
  assign g1721 = \DFF_120.Q ;
  assign g1724 = \DFF_530.Q ;
  assign g1727 = \DFF_370.Q ;
  assign g1730 = \DFF_96.Q ;
  assign g1733 = \DFF_321.Q ;
  assign g1736 = \DFF_21.Q ;
  assign g1737 = \DFF_25.Q ;
  assign g1738 = \DFF_272.Q ;
  assign g174 = \DFF_102.Q ;
  assign g1741 = \DFF_131.Q ;
  assign g1744 = \DFF_9.Q ;
  assign g1747 = \DFF_388.Q ;
  assign g1750 = \DFF_501.Q ;
  assign g1753 = \DFF_200.Q ;
  assign g1756 = \DFF_410.Q ;
  assign g1759 = \DFF_78.Q ;
  assign g1762 = \DFF_282.Q ;
  assign g1765 = \DFF_320.Q ;
  assign g1766 = \DFF_103.Q ;
  assign g1771 = \DFF_268.Q ;
  assign g1776 = \DFF_523.Q ;
  assign g178 = \DFF_307.Q ;
  assign g1781 = \DFF_332.Q ;
  assign g1786 = \DFF_59.Q ;
  assign g1791 = \DFF_75.Q ;
  assign g1796 = \DFF_324.Q ;
  assign g1801 = \DFF_104.Q ;
  assign g1806 = \DFF_346.Q ;
  assign g1810 = \DFF_233.Q ;
  assign g1811 = \DFF_420.Q ;
  assign g1814 = \DFF_297.Q ;
  assign g182 = \DFF_364.Q ;
  assign g1822 = \DFF_302.Q ;
  assign g1828 = \DFF_369.Q ;
  assign g1834 = \DFF_455.Q ;
  assign g1840 = \DFF_223.Q ;
  assign g1845 = \DFF_352.Q ;
  assign g1848 = \DFF_385.Q ;
  assign g1849 = \DFF_330.Q ;
  assign g1850 = \DFF_252.Q ;
  assign g1853 = \DFF_489.Q ;
  assign g1854 = \DFF_311.Q ;
  assign g1857 = \DFF_178.Q ;
  assign g186 = \DFF_105.Q ;
  assign g1861 = \DFF_141.Q ;
  assign g1864 = \DFF_18.Q ;
  assign g1868 = \DFF_111.Q ;
  assign g1872 = \DFF_449.Q ;
  assign g1878 = \DFF_532.Q ;
  assign g1882 = \DFF_1.Q ;
  assign g1887 = \DFF_349.Q ;
  assign g1891 = \DFF_354.Q ;
  assign g1896 = \DFF_85.Q ;
  assign g1900 = \DFF_333.Q ;
  assign g1905 = \DFF_493.Q ;
  assign g1909 = \DFF_461.Q ;
  assign g1914 = \DFF_209.Q ;
  assign g1918 = \DFF_300.Q ;
  assign g192 = \DFF_284.Q ;
  assign g1923 = \DFF_339.Q ;
  assign g1927 = \DFF_44.Q ;
  assign g1932 = \DFF_373.Q ;
  assign g1936 = \DFF_212.Q ;
  assign g1941 = \DFF_313.Q ;
  assign g1945 = \DFF_271.Q ;
  assign g1950 = \DFF_155.Q ;
  assign g1955 = \DFF_462.Q ;
  assign g1956 = \DFF_156.Q ;
  assign g1957 = \DFF_304.Q ;
  assign g1958 = \DFF_318.Q ;
  assign g1959 = \DFF_275.Q ;
  assign g197 = \DFF_424.Q ;
  assign g2004 = \DFF_269.Q ;
  assign g201 = \DFF_400.Q ;
  assign g2044 = \DFF_318.Q ;
  assign g2056 = \DFF_464.Q ;
  assign g2068 = \DFF_502.Q ;
  assign g2069 = \DFF_397.Q ;
  assign g207 = \DFF_5.Q ;
  assign g2071 = \DFF_161.Q ;
  assign g2072 = \DFF_187.Q ;
  assign g2073 = \DFF_500.Q ;
  assign g2075 = \DFF_476.Q ;
  assign g2076 = \DFF_356.Q ;
  assign g2079 = \DFF_451.Q ;
  assign g2080 = \DFF_446.Q ;
  assign g2084 = \DFF_411.Q ;
  assign g2085 = \DFF_193.Q ;
  assign g2086 = \DFF_380.Q ;
  assign g2089 = \DFF_464.Q ;
  assign g2090 = \DFF_443.Q ;
  assign g2094 = \DFF_4.Q ;
  assign g2097 = \DFF_502.Q ;
  assign g2098 = \DFF_244.Q ;
  assign g2100 = \DFF_187.Q ;
  assign g2101 = \DFF_222.Q ;
  assign g2103 = \DFF_246.Q ;
  assign g2108 = g1170;
  assign g2110 = g1173;
  assign g2116 = g1176;
  assign g2119 = \DFF_243.Q ;
  assign g2121 = g1179;
  assign g2122 = g1182;
  assign g2123 = g1185;
  assign g2124 = \DFF_126.Q ;
  assign g2125 = g1188;
  assign g213 = \DFF_331.Q ;
  assign g2130 = g1961;
  assign g2131 = g1191;
  assign g2135 = \DFF_276.Q ;
  assign g2154 = \DFF_168.Q ;
  assign g2155 = g1194;
  assign g2156 = \DFF_384.Q ;
  assign g2158 = \DFF_242.Q ;
  assign g2159 = \DFF_228.Q ;
  assign g2162 = \DFF_311.Q ;
  assign g2163 = \DFF_92.Q ;
  assign g2164 = \DFF_350.Q ;
  assign g2165 = \DFF_116.Q ;
  assign g2166 = g1960;
  assign g2168 = \DFF_22.Q ;
  assign g2171 = \DFF_319.Q ;
  assign g2173 = \DFF_43.Q ;
  assign g2181 = \DFF_72.Q ;
  assign g219 = \DFF_125.Q ;
  assign g2190 = \DFF_237.Q ;
  assign g22 = g18;
  assign g2206 = \DFF_90.Q ;
  assign g2207 = \DFF_63.Q ;
  assign g2217 = \DFF_213.Q ;
  assign g2221 = \DFF_296.Q ;
  assign g2225 = \DFF_91.Q ;
  assign g2231 = \DFF_31.Q ;
  assign g2232 = \DFF_109.Q ;
  assign g2233 = \DFF_287.Q ;
  assign g2238 = \DFF_417.Q ;
  assign g2239 = \DFF_513.Q ;
  assign g2242 = g925;
  assign g2243 = \DFF_278.Q ;
  assign g2244 = \DFF_24.Q ;
  assign g2245 = g1700;
  assign g2246 = g5816;
  assign g2247 = \DFF_479.Q ;
  assign g225 = \DFF_132.Q ;
  assign g2252 = \DFF_224.Q ;
  assign g2255 = \DFF_169.Q ;
  assign g2256 = \DFF_533.Q ;
  assign g2258 = \DFF_496.Q ;
  assign g2259 = \DFF_49.Q ;
  assign g2267 = \DFF_363.Q ;
  assign g2269 = g872;
  assign g2270 = g873;
  assign g2296 = \DFF_156.Q ;
  assign g2298 = g1700;
  assign g2304 = \DFF_304.Q ;
  assign g231 = \DFF_185.Q ;
  assign g2322 = \DFF_178.Q ;
  assign g2329 = g886;
  assign g2334 = g889;
  assign g2335 = \DFF_158.Q ;
  assign g2337 = g892;
  assign g2339 = g895;
  assign g2341 = \DFF_360.Q ;
  assign g2342 = g898;
  assign g2344 = g901;
  assign g2346 = g904;
  assign g2348 = g907;
  assign g2349 = \DFF_159.Q ;
  assign g2350 = g910;
  assign g2351 = g913;
  assign g2352 = g916;
  assign g2355 = g18;
  assign g2356 = g18;
  assign g2363 = g919;
  assign g2368 = g922;
  assign g237 = \DFF_303.Q ;
  assign g2390 = \DFF_0.Q ;
  assign g2391 = \DFF_299.Q ;
  assign g2411 = \DFF_276.Q ;
  assign g2418 = \DFF_476.Q ;
  assign g243 = \DFF_33.Q ;
  assign g2431 = \DFF_451.Q ;
  assign g2432 = \DFF_270.Q ;
  assign g2436 = \DFF_411.Q ;
  assign g2454 = \DFF_441.Q ;
  assign g2462 = g109;
  assign g2478 = \DFF_320.D ;
  assign g248 = \DFF_76.Q ;
  assign g2480 = \DFF_188.Q ;
  assign g2482 = \DFF_174.Q ;
  assign g2502 = g1197;
  assign g2507 = g1200;
  assign g2509 = g1203;
  assign g2523 = \DFF_83.Q ;
  assign g2529 = \DFF_340.Q ;
  assign g253 = \DFF_397.Q ;
  assign g2530 = \DFF_460.Q ;
  assign g2537 = \DFF_13.Q ;
  assign g2539 = \DFF_50.Q ;
  assign g254 = \DFF_246.Q ;
  assign g2540 = \DFF_186.Q ;
  assign g2541 = \DFF_260.Q ;
  assign g2543 = \DFF_208.Q ;
  assign g2547 = g3327;
  assign g2548 = \DFF_288.Q ;
  assign g255 = \DFF_270.Q ;
  assign g2554 = \DFF_524.Q ;
  assign g256 = \DFF_500.Q ;
  assign g2560 = \DFF_166.Q ;
  assign g2569 = \DFF_211.Q ;
  assign g257 = \DFF_356.Q ;
  assign g2578 = g27;
  assign g2579 = \DFF_264.Q ;
  assign g258 = \DFF_446.Q ;
  assign g2586 = \DFF_12.Q ;
  assign g259 = \DFF_193.Q ;
  assign g2593 = \DFF_255.Q ;
  assign g260 = \DFF_443.Q ;
  assign g2601 = \DFF_464.Q ;
  assign g2602 = \DFF_476.Q ;
  assign g2603 = \DFF_451.Q ;
  assign g2604 = \DFF_411.Q ;
  assign g2605 = \DFF_502.Q ;
  assign g2606 = \DFF_187.Q ;
  assign g2607 = \DFF_476.Q ;
  assign g2608 = \DFF_451.Q ;
  assign g2609 = \DFF_411.Q ;
  assign g261 = \DFF_244.Q ;
  assign g2610 = \DFF_464.Q ;
  assign g2611 = \DFF_502.Q ;
  assign g2612 = \DFF_187.Q ;
  assign g2613 = \DFF_360.Q ;
  assign g2614 = \DFF_227.Q ;
  assign g2617 = \DFF_429.Q ;
  assign g262 = \DFF_222.Q ;
  assign g2620 = \DFF_389.Q ;
  assign g2623 = \DFF_127.Q ;
  assign g2626 = \DFF_393.Q ;
  assign g2629 = \DFF_184.Q ;
  assign g263 = \DFF_386.Q ;
  assign g2632 = \DFF_387.Q ;
  assign g2635 = \DFF_99.Q ;
  assign g2638 = \DFF_156.Q ;
  assign g2639 = \DFF_304.Q ;
  assign g2640 = \DFF_112.Q ;
  assign g2641 = \DFF_407.Q ;
  assign g2642 = \DFF_149.Q ;
  assign g2643 = \DFF_253.Q ;
  assign g2644 = \DFF_30.Q ;
  assign g2645 = \DFF_247.Q ;
  assign g2646 = \DFF_301.Q ;
  assign g2647 = \DFF_38.Q ;
  assign g2648 = \DFF_269.Q ;
  assign g2649 = \DFF_243.Q ;
  assign g2650 = \DFF_83.Q ;
  assign g2651 = \DFF_340.Q ;
  assign g2652 = \DFF_294.Q ;
  assign g2653 = \DFF_14.Q ;
  assign g2654 = \DFF_52.Q ;
  assign g2655 = \DFF_158.Q ;
  assign g266 = \DFF_485.Q ;
  assign g2662 = \DFF_31.Q ;
  assign g2669 = \DFF_417.Q ;
  assign g2677 = \DFF_103.Q ;
  assign g2683 = \DFF_268.Q ;
  assign g2689 = \DFF_523.Q ;
  assign g269 = \DFF_176.Q ;
  assign g2695 = \DFF_332.Q ;
  assign g2701 = \DFF_59.Q ;
  assign g2707 = \DFF_75.Q ;
  assign g2713 = \DFF_324.Q ;
  assign g2719 = \DFF_104.Q ;
  assign g272 = \DFF_345.Q ;
  assign g2725 = \DFF_344.Q ;
  assign g2726 = \DFF_470.Q ;
  assign g2727 = \DFF_198.Q ;
  assign g2728 = g1696;
  assign g2731 = \DFF_311.Q ;
  assign g2732 = \DFF_446.Q ;
  assign g2733 = g109;
  assign g2742 = \DFF_193.Q ;
  assign g2745 = g18;
  assign g2748 = \DFF_443.Q ;
  assign g275 = \DFF_390.Q ;
  assign g2750 = \DFF_244.Q ;
  assign g2751 = \DFF_222.Q ;
  assign g2752 = g1197;
  assign g2755 = \DFF_246.Q ;
  assign g2757 = g1200;
  assign g2758 = \DFF_270.Q ;
  assign g2759 = g1203;
  assign g2765 = \DFF_346.Q ;
  assign g2771 = \DFF_83.Q ;
  assign g2772 = \DFF_13.Q ;
  assign g2773 = \DFF_340.Q ;
  assign g2775 = \DFF_13.Q ;
  assign g2779 = \DFF_191.Q ;
  assign g278 = \DFF_46.Q ;
  assign g2791 = g4171;
  assign g2797 = \DFF_293.Q ;
  assign g2798 = \DFF_434.Q ;
  assign g2809 = \DFF_63.Q ;
  assign g281 = \DFF_133.Q ;
  assign g2814 = \DFF_213.Q ;
  assign g2817 = \DFF_460.Q ;
  assign g2821 = \DFF_91.Q ;
  assign g2824 = \DFF_50.Q ;
  assign g2829 = \DFF_287.Q ;
  assign g2833 = \DFF_186.Q ;
  assign g284 = \DFF_123.Q ;
  assign g2840 = \DFF_513.Q ;
  assign g2844 = \DFF_260.Q ;
  assign g2847 = \DFF_479.Q ;
  assign g2851 = \DFF_208.Q ;
  assign g2855 = \DFF_224.Q ;
  assign g2861 = \DFF_288.Q ;
  assign g2864 = \DFF_275.D ;
  assign g2868 = \DFF_533.Q ;
  assign g287 = \DFF_259.Q ;
  assign g2873 = \DFF_524.Q ;
  assign g2874 = \DFF_496.Q ;
  assign g2877 = \DFF_49.Q ;
  assign g2883 = \DFF_166.Q ;
  assign g2885 = \DFF_363.Q ;
  assign g2891 = \DFF_211.Q ;
  assign g290 = \DFF_251.Q ;
  assign g2902 = g5816;
  assign g2906 = g872;
  assign g2908 = \DFF_159.Q ;
  assign g2909 = g1170;
  assign g2914 = g873;
  assign g2915 = g1173;
  assign g2916 = \DFF_299.Q ;
  assign g293 = \DFF_197.Q ;
  assign g2937 = g1176;
  assign g2942 = g1179;
  assign g2949 = g1182;
  assign g2952 = \DFF_347.Q ;
  assign g2955 = \DFF_243.Q ;
  assign g2956 = g1185;
  assign g2958 = g3327;
  assign g296 = \DFF_279.Q ;
  assign g2960 = g1188;
  assign g2962 = g1191;
  assign g2964 = g1194;
  assign g2965 = g109;
  assign g2971 = \DFF_352.Q ;
  assign g2980 = g750;
  assign g2986 = \DFF_291.Q ;
  assign g299 = \DFF_511.Q ;
  assign g2994 = \DFF_431.Q ;
  assign g3007 = \DFF_53.Q ;
  assign g3012 = g109;
  assign g302 = \DFF_229.Q ;
  assign g3038 = \DFF_86.Q ;
  assign g3044 = g109;
  assign g305 = \DFF_265.Q ;
  assign g3067 = \DFF_174.Q ;
  assign g3069 = \DFF_328.Q ;
  assign g3076 = \DFF_31.Q ;
  assign g3077 = \DFF_278.Q ;
  assign g3088 = \DFF_417.Q ;
  assign g309 = \DFF_183.Q ;
  assign g3093 = g925;
  assign g3094 = \DFF_278.Q ;
  assign g3119 = g109;
  assign g312 = \DFF_2.Q ;
  assign g315 = \DFF_41.Q ;
  assign g3164 = g18;
  assign g318 = \DFF_225.Q ;
  assign g32 = \DFF_92.Q ;
  assign g3206 = \DFF_155.Q ;
  assign g321 = \DFF_478.Q ;
  assign g3213 = g886;
  assign g3214 = \DFF_320.D ;
  assign g3219 = g889;
  assign g3220 = \DFF_158.Q ;
  assign g3226 = g892;
  assign g3227 = g895;
  assign g3228 = g18;
  assign g324 = \DFF_467.Q ;
  assign g3252 = g898;
  assign g3253 = g901;
  assign g3255 = g904;
  assign g3256 = g109;
  assign g3260 = g907;
  assign g3262 = g910;
  assign g3266 = g913;
  assign g3267 = g916;
  assign g327 = \DFF_65.Q ;
  assign g3271 = g919;
  assign g3272 = \DFF_506.Q ;
  assign g3274 = g922;
  assign g3292 = \DFF_152.Q ;
  assign g33 = \DFF_168.Q ;
  assign g330 = \DFF_239.Q ;
  assign g3306 = \DFF_397.Q ;
  assign g3307 = g109;
  assign g3318 = \DFF_275.D ;
  assign g3321 = \DFF_500.Q ;
  assign g3323 = \DFF_372.Q ;
  assign g3326 = \DFF_356.Q ;
  assign g3328 = g27;
  assign g3329 = \DFF_320.D ;
  assign g333 = \DFF_175.Q ;
  assign g3331 = g916;
  assign g3334 = g919;
  assign g3344 = g922;
  assign g3353 = g109;
  assign g336 = \DFF_263.Q ;
  assign g3364 = g109;
  assign g3371 = g1961;
  assign g3372 = g109;
  assign g3373 = \DFF_227.Q ;
  assign g3379 = g109;
  assign g3380 = \DFF_429.Q ;
  assign g3381 = \DFF_291.D ;
  assign g3385 = g109;
  assign g3386 = g109;
  assign g3387 = \DFF_389.Q ;
  assign g339 = \DFF_499.Q ;
  assign g3390 = \DFF_420.Q ;
  assign g3391 = g18;
  assign g3392 = g109;
  assign g3393 = g109;
  assign g3394 = \DFF_127.Q ;
  assign g3397 = g18;
  assign g3398 = g18;
  assign g3399 = g6920;
  assign g34 = \DFF_384.Q ;
  assign g3404 = g109;
  assign g3405 = g109;
  assign g3406 = \DFF_393.Q ;
  assign g3407 = g5658;
  assign g3413 = g18;
  assign g3414 = g6926;
  assign g3415 = g109;
  assign g3416 = g109;
  assign g3417 = \DFF_184.Q ;
  assign g3418 = g5659;
  assign g342 = \DFF_230.Q ;
  assign g3424 = g18;
  assign g3425 = g6932;
  assign g3426 = g109;
  assign g3427 = g109;
  assign g3428 = \DFF_387.Q ;
  assign g3431 = g6942;
  assign g3432 = g109;
  assign g3433 = \DFF_99.Q ;
  assign g3435 = g6949;
  assign g3436 = g109;
  assign g3437 = \DFF_347.Q ;
  assign g3438 = g6955;
  assign g3439 = g109;
  assign g345 = \DFF_266.Q ;
  assign g3458 = g109;
  assign g3459 = g1197;
  assign g3461 = g1200;
  assign g3462 = \DFF_431.D ;
  assign g3473 = g1203;
  assign g3474 = g5816;
  assign g348 = \DFF_440.Q ;
  assign g35 = \DFF_242.Q ;
  assign g3506 = \DFF_53.D ;
  assign g351 = \DFF_79.Q ;
  assign g3524 = \DFF_122.D ;
  assign g3538 = \DFF_397.Q ;
  assign g354 = \DFF_70.Q ;
  assign g3545 = \DFF_500.Q ;
  assign g357 = \DFF_216.Q ;
  assign g3583 = \DFF_356.Q ;
  assign g36 = \DFF_228.Q ;
  assign g360 = \DFF_283.Q ;
  assign g3621 = g872;
  assign g3622 = \DFF_446.Q ;
  assign g3624 = g873;
  assign g3627 = \DFF_193.Q ;
  assign g363 = \DFF_238.Q ;
  assign g3630 = \DFF_443.Q ;
  assign g3632 = \DFF_244.Q ;
  assign g3633 = \DFF_222.Q ;
  assign g3636 = \DFF_246.Q ;
  assign g3637 = \DFF_270.Q ;
  assign g366 = \DFF_308.Q ;
  assign g3663 = g1170;
  assign g3682 = g109;
  assign g3683 = g1173;
  assign g369 = \DFF_19.Q ;
  assign g3693 = g109;
  assign g3694 = g1176;
  assign g3697 = \DFF_275.D ;
  assign g37 = \DFF_350.Q ;
  assign g3703 = g109;
  assign g3704 = g1179;
  assign g3705 = g109;
  assign g3707 = g109;
  assign g3708 = g1182;
  assign g3715 = g109;
  assign g3716 = g1185;
  assign g3719 = g109;
  assign g3720 = g1188;
  assign g3721 = g1191;
  assign g3726 = g1194;
  assign g3729 = \DFF_431.Q ;
  assign g3737 = \DFF_360.Q ;
  assign g374 = \DFF_207.Q ;
  assign g3761 = g4171;
  assign g378 = \DFF_409.Q ;
  assign g38 = \DFF_116.Q ;
  assign g3817 = \DFF_159.Q ;
  assign g382 = \DFF_483.Q ;
  assign g3828 = g109;
  assign g386 = \DFF_217.Q ;
  assign g3861 = g925;
  assign g3862 = g109;
  assign g3874 = g109;
  assign g3878 = g109;
  assign g39 = \DFF_22.Q ;
  assign g3905 = g109;
  assign g3909 = g109;
  assign g391 = \DFF_394.Q ;
  assign g3913 = g109;
  assign g3938 = \DFF_77.Q ;
  assign g3940 = g109;
  assign g3944 = g109;
  assign g3946 = g18;
  assign g396 = \DFF_114.Q ;
  assign g3975 = g109;
  assign g3980 = g109;
  assign g3982 = \DFF_311.Q ;
  assign g3988 = g109;
  assign g3990 = g109;
  assign g3995 = g109;
  assign g3996 = g109;
  assign g3997 = \DFF_112.Q ;
  assign g4 = \DFF_29.Q ;
  assign g40 = \DFF_319.Q ;
  assign g4002 = g109;
  assign g4003 = g109;
  assign g4004 = \DFF_407.Q ;
  assign g4005 = \DFF_227.Q ;
  assign g401 = \DFF_177.Q ;
  assign g4010 = g109;
  assign g4011 = \DFF_149.Q ;
  assign g4012 = \DFF_429.Q ;
  assign g4049 = g109;
  assign g4050 = \DFF_253.Q ;
  assign g4051 = \DFF_389.Q ;
  assign g4055 = g109;
  assign g4056 = \DFF_30.Q ;
  assign g4057 = \DFF_127.Q ;
  assign g406 = \DFF_419.Q ;
  assign g4060 = g109;
  assign g4061 = \DFF_247.Q ;
  assign g4062 = \DFF_393.Q ;
  assign g4066 = \DFF_301.Q ;
  assign g4067 = \DFF_184.Q ;
  assign g4076 = \DFF_77.D ;
  assign g4077 = \DFF_38.Q ;
  assign g4078 = \DFF_387.Q ;
  assign g4080 = g1960;
  assign g4081 = \DFF_434.Q ;
  assign g4082 = \DFF_99.Q ;
  assign g4083 = \DFF_347.Q ;
  assign g4087 = g886;
  assign g4089 = \DFF_471.D ;
  assign g4095 = \DFF_460.Q ;
  assign g4096 = g889;
  assign g4098 = \DFF_50.Q ;
  assign g4102 = g892;
  assign g4105 = \DFF_186.Q ;
  assign g411 = \DFF_491.Q ;
  assign g4113 = g895;
  assign g4114 = \DFF_328.D ;
  assign g4116 = \DFF_260.Q ;
  assign g4117 = \DFF_262.D ;
  assign g4121 = g898;
  assign g4124 = \DFF_208.Q ;
  assign g4125 = g901;
  assign g4127 = \DFF_288.Q ;
  assign g4140 = g904;
  assign g4142 = \DFF_524.Q ;
  assign g4156 = g907;
  assign g4159 = \DFF_166.Q ;
  assign g416 = \DFF_204.Q ;
  assign g4160 = g910;
  assign g4166 = \DFF_211.Q ;
  assign g4167 = g913;
  assign g4172 = \DFF_431.Q ;
  assign g4173 = \DFF_112.Q ;
  assign g4174 = \DFF_407.Q ;
  assign g4175 = \DFF_149.Q ;
  assign g4176 = \DFF_253.Q ;
  assign g4177 = \DFF_30.Q ;
  assign g4178 = \DFF_247.Q ;
  assign g4179 = \DFF_301.Q ;
  assign g4180 = \DFF_38.Q ;
  assign g4181 = \DFF_434.Q ;
  assign g4182 = \DFF_227.Q ;
  assign g4183 = \DFF_429.Q ;
  assign g4184 = \DFF_389.Q ;
  assign g4185 = \DFF_127.Q ;
  assign g4186 = \DFF_393.Q ;
  assign g4187 = \DFF_184.Q ;
  assign g4188 = \DFF_387.Q ;
  assign g4189 = \DFF_99.Q ;
  assign g4190 = \DFF_347.Q ;
  assign g4191 = g886;
  assign g4192 = g889;
  assign g4193 = g892;
  assign g4194 = g895;
  assign g4195 = g898;
  assign g4196 = g925;
  assign g4197 = g901;
  assign g4198 = g904;
  assign g4199 = g907;
  assign g4200 = g910;
  assign g4201 = g913;
  assign g4202 = g916;
  assign g4203 = g919;
  assign g4204 = g922;
  assign g4205 = g1170;
  assign g4206 = g1197;
  assign g4207 = g1200;
  assign g4208 = g1203;
  assign g4209 = g1173;
  assign g421 = \DFF_406.Q ;
  assign g4210 = g1176;
  assign g4211 = g1179;
  assign g4212 = g1182;
  assign g4213 = g1185;
  assign g4214 = g1188;
  assign g4215 = g1191;
  assign g4216 = g1194;
  assign g4217 = \DFF_275.D ;
  assign g4219 = \DFF_174.Q ;
  assign g4231 = \DFF_272.D ;
  assign g4232 = g1961;
  assign g4238 = \DFF_131.D ;
  assign g4239 = \DFF_9.D ;
  assign g4255 = \DFF_388.D ;
  assign g426 = \DFF_124.Q ;
  assign g4264 = \DFF_501.D ;
  assign g4268 = \DFF_460.Q ;
  assign g4271 = \DFF_113.Q ;
  assign g4274 = \DFF_200.D ;
  assign g4279 = \DFF_50.Q ;
  assign g4283 = \DFF_410.D ;
  assign g4287 = \DFF_186.Q ;
  assign g4293 = \DFF_78.D ;
  assign g4295 = g1960;
  assign g4296 = \DFF_260.Q ;
  assign g4309 = \DFF_282.D ;
  assign g431 = \DFF_492.Q ;
  assign g4310 = \DFF_208.Q ;
  assign g4317 = \DFF_288.Q ;
  assign g4322 = \DFF_524.Q ;
  assign g4325 = \DFF_438.D ;
  assign g4327 = \DFF_166.Q ;
  assign g4330 = \DFF_232.D ;
  assign g4331 = \DFF_211.Q ;
  assign g4334 = \DFF_525.D ;
  assign g4335 = \DFF_159.Q ;
  assign g4338 = \DFF_240.D ;
  assign g4340 = \DFF_7.D ;
  assign g4342 = \DFF_383.D ;
  assign g435 = \DFF_512.Q ;
  assign g4351 = \DFF_122.D ;
  assign g4352 = g5816;
  assign g440 = \DFF_378.Q ;
  assign g4414 = g5658;
  assign g4425 = g5659;
  assign g4437 = \DFF_113.Q ;
  assign g444 = \DFF_171.Q ;
  assign g4443 = \DFF_113.Q ;
  assign g4452 = \DFF_113.Q ;
  assign g4456 = \DFF_113.Q ;
  assign g4458 = g6920;
  assign g4462 = g6926;
  assign g4464 = g6932;
  assign g4465 = \DFF_214.D ;
  assign g4469 = g6942;
  assign g4471 = \DFF_457.D ;
  assign g4472 = g6949;
  assign g4473 = \DFF_399.D ;
  assign g4475 = g6955;
  assign g4477 = \DFF_366.D ;
  assign g448 = \DFF_368.Q ;
  assign g4480 = \DFF_145.D ;
  assign g4484 = \DFF_353.D ;
  assign g4485 = g109;
  assign g4490 = \DFF_468.D ;
  assign g4491 = g109;
  assign g4495 = \DFF_77.D ;
  assign g4496 = \DFF_227.Q ;
  assign g4498 = \DFF_416.D ;
  assign g4499 = g109;
  assign g4500 = \DFF_241.D ;
  assign g4504 = \DFF_429.Q ;
  assign g4506 = \DFF_517.D ;
  assign g4507 = g109;
  assign g4510 = \DFF_389.Q ;
  assign g4513 = g109;
  assign g452 = \DFF_3.Q ;
  assign g4520 = \DFF_127.Q ;
  assign g4523 = g109;
  assign g4526 = g873;
  assign g4533 = \DFF_393.Q ;
  assign g4541 = \DFF_184.Q ;
  assign g4549 = \DFF_387.Q ;
  assign g4555 = \DFF_99.Q ;
  assign g4556 = \DFF_0.D ;
  assign g456 = \DFF_264.Q ;
  assign g4562 = \DFF_347.Q ;
  assign g4577 = g872;
  assign g4589 = \DFF_431.D ;
  assign g4590 = \DFF_328.D ;
  assign g461 = \DFF_12.Q ;
  assign g4615 = \DFF_262.D ;
  assign g4637 = \DFF_53.D ;
  assign g466 = \DFF_255.Q ;
  assign g4674 = \DFF_471.D ;
  assign g4678 = g109;
  assign g4681 = g109;
  assign g471 = \DFF_152.Q ;
  assign g4711 = \DFF_291.D ;
  assign g4713 = g109;
  assign g4716 = g109;
  assign g4721 = g109;
  assign g4726 = g109;
  assign g4728 = \DFF_397.Q ;
  assign g4730 = g109;
  assign g4733 = \DFF_500.Q ;
  assign g4735 = g109;
  assign g4746 = \DFF_356.Q ;
  assign g4748 = g109;
  assign g4757 = \DFF_446.Q ;
  assign g476 = \DFF_379.Q ;
  assign g4762 = \DFF_193.Q ;
  assign g4767 = \DFF_443.Q ;
  assign g4773 = \DFF_244.Q ;
  assign g4781 = \DFF_222.Q ;
  assign g4785 = g18;
  assign g4786 = \DFF_246.Q ;
  assign g4789 = g18;
  assign g4790 = g18;
  assign g4791 = \DFF_270.Q ;
  assign g4802 = g18;
  assign g4805 = g18;
  assign g481 = \DFF_430.Q ;
  assign g486 = \DFF_151.Q ;
  assign g4887 = g1961;
  assign g4888 = g1960;
  assign g4890 = \DFF_136.D ;
  assign g4891 = \DFF_117.D ;
  assign g4892 = \DFF_157.D ;
  assign g4893 = \DFF_191.D ;
  assign g4894 = \DFF_262.D ;
  assign g4895 = \DFF_431.D ;
  assign g4896 = \DFF_53.D ;
  assign g4897 = \DFF_291.D ;
  assign g4898 = \DFF_328.D ;
  assign g49 = \DFF_496.Q ;
  assign g4901 = \DFF_471.D ;
  assign g4902 = \DFF_330.D ;
  assign g4903 = \DFF_252.D ;
  assign g4904 = \DFF_489.D ;
  assign g4905 = \DFF_352.D ;
  assign g4906 = \DFF_122.D ;
  assign g4907 = \DFF_77.D ;
  assign g4908 = g102;
  assign g491 = \DFF_329.Q ;
  assign g4915 = g103;
  assign g4933 = \DFF_113.Q ;
  assign g4934 = \DFF_122.D ;
  assign g4935 = g104;
  assign g4940 = \DFF_112.D ;
  assign g4942 = \DFF_113.Q ;
  assign g4944 = g28;
  assign g4951 = \DFF_113.Q ;
  assign g4954 = g29;
  assign g496 = \DFF_51.Q ;
  assign g4961 = \DFF_113.Q ;
  assign g4963 = g5816;
  assign g4970 = g84;
  assign g5007 = \DFF_272.D ;
  assign g501 = \DFF_221.Q ;
  assign g5011 = \DFF_131.D ;
  assign g5012 = \DFF_9.D ;
  assign g5027 = \DFF_388.D ;
  assign g5032 = \DFF_501.D ;
  assign g5033 = \DFF_200.D ;
  assign g5035 = \DFF_410.D ;
  assign g5037 = \DFF_78.D ;
  assign g5040 = \DFF_282.D ;
  assign g5047 = g42;
  assign g5050 = g6920;
  assign g5052 = g48;
  assign g506 = \DFF_459.Q ;
  assign g5063 = g43;
  assign g5066 = g6926;
  assign g5069 = g44;
  assign g5072 = g6932;
  assign g5075 = g96;
  assign g5078 = g45;
  assign g5081 = g6942;
  assign g5083 = \DFF_372.D ;
  assign g5085 = g46;
  assign g5088 = g6949;
  assign g5091 = g47;
  assign g5094 = g6955;
  assign g5101 = g872;
  assign g5102 = g872;
  assign g5105 = g873;
  assign g5106 = g873;
  assign g5107 = g100;
  assign g5109 = \DFF_438.D ;
  assign g511 = \DFF_529.Q ;
  assign g5111 = \DFF_232.D ;
  assign g5114 = \DFF_525.D ;
  assign g5120 = \DFF_240.D ;
  assign g5126 = \DFF_31.D ;
  assign g5127 = \DFF_7.D ;
  assign g5128 = g109;
  assign g5148 = \DFF_417.D ;
  assign g5149 = \DFF_383.D ;
  assign g5151 = g109;
  assign g516 = \DFF_245.Q ;
  assign g5173 = \DFF_278.D ;
  assign g5194 = \DFF_323.D ;
  assign g5195 = g99;
  assign g5197 = \DFF_347.Q ;
  assign g5198 = g5658;
  assign g52 = \DFF_63.Q ;
  assign g5205 = g31;
  assign g521 = \DFF_447.Q ;
  assign g5210 = g5659;
  assign g5218 = \DFF_174.Q ;
  assign g5236 = g30;
  assign g5241 = g83;
  assign g5245 = g82;
  assign g525 = \DFF_475.Q ;
  assign g5253 = \DFF_168.Q ;
  assign g5262 = \DFF_384.Q ;
  assign g5265 = \DFF_242.Q ;
  assign g5270 = \DFF_228.Q ;
  assign g5272 = \DFF_270.Q ;
  assign g5275 = \DFF_350.Q ;
  assign g5281 = g86;
  assign g5284 = \DFF_116.Q ;
  assign g5287 = g6842;
  assign g5288 = g87;
  assign g5291 = \DFF_22.Q ;
  assign g5296 = g88;
  assign g5299 = \DFF_319.Q ;
  assign g530 = \DFF_210.Q ;
  assign g5301 = g89;
  assign g5305 = g90;
  assign g5314 = g91;
  assign g5320 = g85;
  assign g534 = \DFF_522.Q ;
  assign g5344 = \DFF_214.D ;
  assign g5348 = \DFF_457.D ;
  assign g5353 = \DFF_399.D ;
  assign g5354 = g109;
  assign g538 = \DFF_203.Q ;
  assign g5390 = \DFF_158.D ;
  assign g5391 = \DFF_366.D ;
  assign g5392 = \DFF_21.D ;
  assign g5395 = \DFF_145.D ;
  assign g5396 = \DFF_174.D ;
  assign g5397 = \DFF_270.Q ;
  assign g5401 = \DFF_353.D ;
  assign g5402 = \DFF_0.D ;
  assign g5404 = \DFF_113.D ;
  assign g5415 = \DFF_468.D ;
  assign g5416 = \DFF_416.D ;
  assign g5417 = \DFF_241.D ;
  assign g5419 = \DFF_517.D ;
  assign g542 = \DFF_205.Q ;
  assign g5421 = \DFF_179.D ;
  assign g5445 = \DFF_531.D ;
  assign g546 = \DFF_460.Q ;
  assign g5471 = \DFF_92.Q ;
  assign g5486 = g92;
  assign g549 = \DFF_159.Q ;
  assign g5494 = g93;
  assign g55 = \DFF_213.Q ;
  assign g5504 = g94;
  assign g5509 = \DFF_262.D ;
  assign g5511 = \DFF_113.Q ;
  assign g5515 = g95;
  assign g5529 = \DFF_407.D ;
  assign g5536 = \DFF_149.D ;
  assign g554 = \DFF_50.Q ;
  assign g5543 = \DFF_389.D ;
  assign g5556 = \DFF_318.D ;
  assign g5567 = \DFF_397.Q ;
  assign g5568 = \DFF_500.Q ;
  assign g557 = \DFF_186.Q ;
  assign g5572 = \DFF_356.Q ;
  assign g5586 = \DFF_446.Q ;
  assign g5589 = \DFF_193.Q ;
  assign g5593 = \DFF_443.Q ;
  assign g5596 = \DFF_244.Q ;
  assign g560 = \DFF_260.Q ;
  assign g5603 = \DFF_222.Q ;
  assign g5615 = \DFF_246.Q ;
  assign g5620 = g41;
  assign g563 = \DFF_208.Q ;
  assign g5633 = g101;
  assign g5643 = \DFF_397.Q ;
  assign g5644 = \DFF_270.Q ;
  assign g5645 = \DFF_500.Q ;
  assign g5646 = \DFF_356.Q ;
  assign g5647 = \DFF_446.Q ;
  assign g5648 = \DFF_193.Q ;
  assign g5649 = \DFF_443.Q ;
  assign g5650 = \DFF_244.Q ;
  assign g5651 = \DFF_222.Q ;
  assign g5652 = \DFF_246.Q ;
  assign g5653 = \DFF_174.Q ;
  assign g5654 = \DFF_136.D ;
  assign g5655 = \DFF_117.D ;
  assign g5656 = \DFF_157.D ;
  assign g5657 = \DFF_191.D ;
  assign g566 = \DFF_288.Q ;
  assign g5660 = \DFF_0.D ;
  assign g5661 = \DFF_272.D ;
  assign g5662 = \DFF_131.D ;
  assign g5663 = \DFF_9.D ;
  assign g5664 = \DFF_388.D ;
  assign g5665 = \DFF_501.D ;
  assign g5666 = \DFF_200.D ;
  assign g5667 = \DFF_410.D ;
  assign g5668 = \DFF_78.D ;
  assign g5669 = \DFF_282.D ;
  assign g5670 = \DFF_330.D ;
  assign g5671 = \DFF_252.D ;
  assign g5672 = \DFF_489.D ;
  assign g5673 = \DFF_352.D ;
  assign g5676 = g103;
  assign g5677 = g102;
  assign g5679 = g30;
  assign g5682 = g104;
  assign g5683 = g103;
  assign g5685 = g42;
  assign g5688 = g28;
  assign g5689 = g104;
  assign g569 = \DFF_524.Q ;
  assign g5692 = g30;
  assign g5693 = g43;
  assign g5696 = g29;
  assign g5697 = g28;
  assign g5700 = g31;
  assign g5701 = g44;
  assign g5702 = g82;
  assign g5705 = g29;
  assign g5708 = g48;
  assign g5718 = g45;
  assign g5719 = g89;
  assign g572 = \DFF_166.Q ;
  assign g5723 = g46;
  assign g5724 = g90;
  assign g5727 = g47;
  assign g5728 = g83;
  assign g5729 = g91;
  assign g5730 = g101;
  assign g5734 = g48;
  assign g5735 = g92;
  assign g5736 = g102;
  assign g5741 = g84;
  assign g5742 = g93;
  assign g5743 = g103;
  assign g575 = \DFF_211.Q ;
  assign g5751 = g41;
  assign g5752 = g85;
  assign g5753 = g94;
  assign g5754 = g104;
  assign g5755 = \DFF_400.D ;
  assign g5763 = \DFF_226.D ;
  assign g5766 = g86;
  assign g5767 = g95;
  assign g5768 = g28;
  assign g5770 = \DFF_237.D ;
  assign g5777 = \DFF_21.D ;
  assign g5778 = g87;
  assign g5779 = g96;
  assign g578 = \DFF_464.Q ;
  assign g5787 = g88;
  assign g579 = \DFF_502.Q ;
  assign g5794 = g99;
  assign g58 = \DFF_91.Q ;
  assign g580 = \DFF_187.Q ;
  assign g5800 = g100;
  assign g581 = \DFF_476.Q ;
  assign g5811 = g42;
  assign g5815 = g43;
  assign g5817 = g5816;
  assign g582 = \DFF_451.Q ;
  assign g5821 = g44;
  assign g5826 = g45;
  assign g583 = \DFF_411.Q ;
  assign g5830 = g48;
  assign g5839 = g46;
  assign g584 = \DFF_464.Q ;
  assign g5843 = g47;
  assign g5844 = \DFF_112.D ;
  assign g5849 = \DFF_227.D ;
  assign g585 = \DFF_502.Q ;
  assign g5858 = \DFF_531.D ;
  assign g586 = \DFF_187.Q ;
  assign g5862 = g29;
  assign g5864 = g6920;
  assign g5865 = g6926;
  assign g587 = \DFF_476.Q ;
  assign g5874 = g6932;
  assign g5879 = g6942;
  assign g588 = \DFF_451.Q ;
  assign g5884 = g6949;
  assign g5887 = \DFF_179.D ;
  assign g5889 = g6955;
  assign g589 = \DFF_411.Q ;
  assign g590 = \DFF_54.Q ;
  assign g5904 = g109;
  assign g591 = \DFF_358.Q ;
  assign g5910 = \DFF_292.D ;
  assign g5914 = \DFF_27.D ;
  assign g5918 = \DFF_380.D ;
  assign g5919 = g109;
  assign g5936 = \DFF_438.D ;
  assign g5937 = \DFF_318.D ;
  assign g5941 = \DFF_262.D ;
  assign g5943 = \DFF_232.D ;
  assign g5947 = g83;
  assign g5948 = \DFF_525.D ;
  assign g5980 = \DFF_372.D ;
  assign g5982 = \DFF_240.D ;
  assign g5987 = g41;
  assign g599 = \DFF_310.Q ;
  assign g5992 = \DFF_7.D ;
  assign g5994 = \DFF_383.D ;
  assign g5996 = \DFF_397.D ;
  assign g6000 = \DFF_500.D ;
  assign g6002 = \DFF_356.D ;
  assign g6015 = \DFF_446.D ;
  assign g6026 = \DFF_193.D ;
  assign g6030 = \DFF_31.D ;
  assign g6035 = \DFF_443.D ;
  assign g6036 = \DFF_417.D ;
  assign g6038 = \DFF_244.D ;
  assign g6040 = \DFF_278.D ;
  assign g6042 = \DFF_222.D ;
  assign g6045 = \DFF_246.D ;
  assign g6049 = \DFF_270.D ;
  assign g605 = \DFF_362.Q ;
  assign g6051 = \DFF_323.D ;
  assign g6054 = \DFF_376.D ;
  assign g6059 = \DFF_173.D ;
  assign g6068 = \DFF_402.D ;
  assign g6071 = \DFF_94.D ;
  assign g6080 = \DFF_290.D ;
  assign g6088 = \DFF_16.D ;
  assign g6093 = \DFF_56.D ;
  assign g6096 = \DFF_82.D ;
  assign g6099 = \DFF_170.D ;
  assign g61 = \DFF_287.Q ;
  assign g6100 = \DFF_214.D ;
  assign g6103 = \DFF_457.D ;
  assign g6104 = g6842;
  assign g6106 = \DFF_122.D ;
  assign g6107 = \DFF_399.D ;
  assign g6108 = \DFF_366.D ;
  assign g611 = \DFF_135.Q ;
  assign g6110 = \DFF_145.D ;
  assign g6111 = \DFF_174.D ;
  assign g6112 = \DFF_353.D ;
  assign g6114 = \DFF_113.D ;
  assign g6115 = \DFF_468.D ;
  assign g6116 = \DFF_416.D ;
  assign g6117 = \DFF_241.D ;
  assign g6118 = \DFF_517.D ;
  assign g6120 = g83;
  assign g6123 = \DFF_253.D ;
  assign g6126 = \DFF_127.D ;
  assign g6127 = \DFF_158.D ;
  assign g6132 = \DFF_347.Q ;
  assign g6155 = \DFF_276.D ;
  assign g6163 = \DFF_452.D ;
  assign g617 = \DFF_261.Q ;
  assign g6179 = \DFF_473.D ;
  assign g6180 = \DFF_165.D ;
  assign g6193 = \DFF_494.D ;
  assign g6198 = \DFF_97.D ;
  assign g6205 = \DFF_315.D ;
  assign g6215 = \DFF_201.D ;
  assign g6216 = \DFF_24.D ;
  assign g622 = \DFF_43.Q ;
  assign g6224 = \DFF_118.D ;
  assign g6234 = \DFF_169.D ;
  assign g6237 = \DFF_407.D ;
  assign g6241 = g101;
  assign g6242 = \DFF_149.D ;
  assign g6243 = \DFF_429.D ;
  assign g6244 = \DFF_90.D ;
  assign g6248 = g102;
  assign g6249 = g101;
  assign g6251 = \DFF_389.D ;
  assign g6253 = g29;
  assign g6254 = g30;
  assign g6255 = g31;
  assign g6256 = g41;
  assign g6257 = g42;
  assign g6258 = g43;
  assign g6259 = g44;
  assign g6260 = g45;
  assign g6261 = g46;
  assign g6262 = g47;
  assign g6263 = g48;
  assign g6264 = g82;
  assign g6265 = g83;
  assign g6266 = g84;
  assign g6267 = g85;
  assign g6268 = g86;
  assign g6269 = g87;
  assign g627 = \DFF_191.Q ;
  assign g6270 = g88;
  assign g6271 = g89;
  assign g6272 = g90;
  assign g6273 = g91;
  assign g6274 = g92;
  assign g6275 = g93;
  assign g6276 = g94;
  assign g6277 = g95;
  assign g6278 = g96;
  assign g6279 = g99;
  assign g6280 = g100;
  assign g6281 = g101;
  assign g6282 = g102;
  assign g6283 = g103;
  assign g6284 = g104;
  assign g6285 = g28;
  assign g6286 = g101;
  assign g6287 = g102;
  assign g6288 = g103;
  assign g6289 = g104;
  assign g6290 = g28;
  assign g6291 = g29;
  assign g6292 = g101;
  assign g6293 = g102;
  assign g6294 = g103;
  assign g6295 = g104;
  assign g6296 = g28;
  assign g6297 = g29;
  assign g6298 = g83;
  assign g6299 = \DFF_214.D ;
  assign g630 = \DFF_336.Q ;
  assign g6300 = \DFF_438.D ;
  assign g6301 = \DFF_232.D ;
  assign g6302 = \DFF_525.D ;
  assign g6303 = \DFF_240.D ;
  assign g6304 = \DFF_7.D ;
  assign g6305 = \DFF_383.D ;
  assign g6306 = \DFF_457.D ;
  assign g6307 = \DFF_399.D ;
  assign g6308 = \DFF_366.D ;
  assign g6309 = \DFF_145.D ;
  assign g631 = \DFF_136.Q ;
  assign g6310 = \DFF_353.D ;
  assign g6311 = \DFF_468.D ;
  assign g6312 = \DFF_416.D ;
  assign g6313 = \DFF_517.D ;
  assign g632 = \DFF_117.Q ;
  assign g6330 = \DFF_241.D ;
  assign g6331 = \DFF_484.D ;
  assign g6332 = \DFF_424.D ;
  assign g6333 = \DFF_66.D ;
  assign g6334 = \DFF_284.D ;
  assign g6336 = \DFF_174.D ;
  assign g6337 = \DFF_113.D ;
  assign g6338 = g83;
  assign g6339 = \DFF_318.D ;
  assign g6340 = \DFF_380.D ;
  assign g6344 = \DFF_127.D ;
  assign g635 = \DFF_157.Q ;
  assign g636 = \DFF_360.Q ;
  assign g6365 = g42;
  assign g6382 = g43;
  assign g6386 = \DFF_452.D ;
  assign g6388 = \DFF_407.D ;
  assign g639 = \DFF_72.Q ;
  assign g6392 = \DFF_71.D ;
  assign g6396 = \DFF_149.D ;
  assign g6397 = \DFF_429.D ;
  assign g6398 = \DFF_473.D ;
  assign g6399 = \DFF_165.D ;
  assign g64 = \DFF_513.Q ;
  assign g6406 = \DFF_389.D ;
  assign g6412 = \DFF_494.D ;
  assign g6419 = \DFF_97.D ;
  assign g6426 = \DFF_315.D ;
  assign g643 = \DFF_518.Q ;
  assign g6433 = \DFF_201.D ;
  assign g6434 = \DFF_24.D ;
  assign g6439 = \DFF_296.D ;
  assign g6442 = \DFF_118.D ;
  assign g6445 = \DFF_169.D ;
  assign g6450 = \DFF_90.D ;
  assign g6453 = \DFF_233.Q ;
  assign g6454 = g48;
  assign g646 = \DFF_64.Q ;
  assign g6468 = \DFF_520.D ;
  assign g6469 = \DFF_140.D ;
  assign g6470 = \DFF_371.D ;
  assign g6471 = \DFF_141.D ;
  assign g6478 = \DFF_17.D ;
  assign g6479 = \DFF_425.D ;
  assign g6480 = \DFF_392.D ;
  assign g6481 = \DFF_456.D ;
  assign g6482 = g44;
  assign g650 = \DFF_403.Q ;
  assign g6500 = \DFF_20.D ;
  assign g6501 = \DFF_218.D ;
  assign g6502 = \DFF_268.D ;
  assign g6503 = g45;
  assign g6506 = \DFF_254.D ;
  assign g6507 = \DFF_81.D ;
  assign g6508 = \DFF_523.D ;
  assign g6509 = g46;
  assign g6513 = \DFF_391.D ;
  assign g6514 = \DFF_466.D ;
  assign g6515 = \DFF_477.D ;
  assign g6516 = \DFF_332.D ;
  assign g6517 = g47;
  assign g6521 = \DFF_400.D ;
  assign g6522 = \DFF_505.D ;
  assign g6523 = \DFF_453.D ;
  assign g6524 = \DFF_138.D ;
  assign g6525 = \DFF_59.D ;
  assign g6526 = \DFF_49.D ;
  assign g6527 = \DFF_237.D ;
  assign g6528 = \DFF_164.D ;
  assign g6529 = \DFF_463.D ;
  assign g6531 = \DFF_363.D ;
  assign g6533 = \DFF_42.D ;
  assign g6534 = \DFF_514.D ;
  assign g6536 = \DFF_112.D ;
  assign g6537 = \DFF_426.D ;
  assign g6538 = \DFF_10.D ;
  assign g6539 = \DFF_227.D ;
  assign g654 = \DFF_196.Q ;
  assign g6541 = \DFF_326.D ;
  assign g6542 = \DFF_256.D ;
  assign g6543 = g872;
  assign g6545 = \DFF_39.D ;
  assign g6546 = \DFF_130.D ;
  assign g6547 = g873;
  assign g6551 = \DFF_258.D ;
  assign g6553 = \DFF_270.D ;
  assign g6558 = \DFF_276.D ;
  assign g6571 = \DFF_531.D ;
  assign g658 = \DFF_395.Q ;
  assign g6584 = \DFF_292.D ;
  assign g6588 = \DFF_27.D ;
  assign g6594 = \DFF_179.D ;
  assign g6596 = g109;
  assign g6620 = \DFF_372.D ;
  assign g6621 = \DFF_63.D ;
  assign g6627 = \DFF_91.D ;
  assign g6629 = g6920;
  assign g6634 = \DFF_226.D ;
  assign g6635 = g6926;
  assign g6638 = \DFF_513.D ;
  assign g664 = \DFF_180.Q ;
  assign g6641 = g6932;
  assign g6644 = \DFF_397.D ;
  assign g6648 = \DFF_226.D ;
  assign g6649 = g6942;
  assign g6652 = \DFF_500.D ;
  assign g6653 = \DFF_224.D ;
  assign g6656 = \DFF_29.D ;
  assign g6657 = g6949;
  assign g6660 = \DFF_356.D ;
  assign g6667 = g6955;
  assign g6670 = \DFF_446.D ;
  assign g6672 = \DFF_336.D ;
  assign g6674 = g48;
  assign g6679 = \DFF_528.D ;
  assign g668 = \DFF_381.Q ;
  assign g6680 = \DFF_193.D ;
  assign g6685 = \DFF_31.D ;
  assign g6686 = \DFF_443.D ;
  assign g6688 = \DFF_417.D ;
  assign g6692 = \DFF_244.D ;
  assign g6694 = \DFF_278.D ;
  assign g6695 = \DFF_222.D ;
  assign g6698 = \DFF_246.D ;
  assign g67 = \DFF_479.Q ;
  assign g6703 = \DFF_21.D ;
  assign g6705 = \DFF_323.D ;
  assign g6706 = \DFF_376.D ;
  assign g6708 = \DFF_173.D ;
  assign g6710 = \DFF_402.D ;
  assign g6715 = \DFF_94.D ;
  assign g6717 = \DFF_290.D ;
  assign g6719 = \DFF_16.D ;
  assign g6723 = \DFF_56.D ;
  assign g6728 = \DFF_30.D ;
  assign g6729 = \DFF_82.D ;
  assign g673 = \DFF_488.Q ;
  assign g6733 = \DFF_393.D ;
  assign g6734 = \DFF_170.D ;
  assign g6735 = g6842;
  assign g6747 = \DFF_289.D ;
  assign g6751 = \DFF_158.D ;
  assign g6755 = \DFF_385.D ;
  assign g6757 = \DFF_220.D ;
  assign g6759 = \DFF_307.D ;
  assign g677 = \DFF_450.Q ;
  assign g6786 = \DFF_364.D ;
  assign g6793 = \DFF_253.D ;
  assign g6795 = \DFF_18.D ;
  assign g6796 = g27;
  assign g6797 = \DFF_112.D ;
  assign g6798 = \DFF_407.D ;
  assign g6799 = \DFF_149.D ;
  assign g6800 = \DFF_227.D ;
  assign g6801 = \DFF_429.D ;
  assign g6802 = \DFF_389.D ;
  assign g6803 = \DFF_376.D ;
  assign g6804 = \DFF_292.D ;
  assign g6805 = \DFF_27.D ;
  assign g6806 = \DFF_173.D ;
  assign g6807 = \DFF_402.D ;
  assign g6808 = \DFF_94.D ;
  assign g6809 = \DFF_290.D ;
  assign g6810 = \DFF_16.D ;
  assign g6811 = \DFF_56.D ;
  assign g6812 = \DFF_82.D ;
  assign g6813 = \DFF_170.D ;
  assign g6814 = \DFF_158.D ;
  assign g6815 = \DFF_31.D ;
  assign g6816 = \DFF_417.D ;
  assign g6817 = \DFF_278.D ;
  assign g6818 = \DFF_226.D ;
  assign g6819 = \DFF_88.D ;
  assign g682 = \DFF_60.Q ;
  assign g6820 = \DFF_303.D ;
  assign g6821 = \DFF_142.D ;
  assign g6822 = \DFF_163.D ;
  assign g6823 = \DFF_132.D ;
  assign g6824 = \DFF_125.D ;
  assign g6825 = \DFF_484.D ;
  assign g6826 = \DFF_67.D ;
  assign g6827 = \DFF_327.D ;
  assign g6828 = \DFF_331.D ;
  assign g6829 = \DFF_487.D ;
  assign g6830 = \DFF_5.D ;
  assign g6831 = \DFF_189.D ;
  assign g6832 = \DFF_105.D ;
  assign g6833 = \DFF_396.D ;
  assign g6834 = \DFF_185.D ;
  assign g6835 = \DFF_424.D ;
  assign g6836 = \DFF_66.D ;
  assign g6837 = \DFF_284.D ;
  assign g6838 = \DFF_153.D ;
  assign g6839 = \DFF_76.D ;
  assign g6840 = \DFF_182.D ;
  assign g6841 = \DFF_33.D ;
  assign g6843 = \DFF_372.D ;
  assign g6844 = \DFF_276.D ;
  assign g6845 = \DFF_323.D ;
  assign g6846 = \DFF_21.D ;
  assign g6852 = \DFF_30.D ;
  assign g6854 = \DFF_393.D ;
  assign g6857 = \DFF_385.D ;
  assign g686 = \DFF_316.Q ;
  assign g6860 = g41;
  assign g6869 = \DFF_289.D ;
  assign g6877 = \DFF_253.D ;
  assign g6881 = \DFF_127.D ;
  assign g6888 = \DFF_220.D ;
  assign g6893 = \DFF_307.D ;
  assign g6894 = \DFF_413.D ;
  assign g6895 = \DFF_515.D ;
  assign g6896 = \DFF_364.D ;
  assign g6897 = \DFF_386.D ;
  assign g6898 = \DFF_497.D ;
  assign g6900 = \DFF_485.D ;
  assign g6901 = \DFF_259.D ;
  assign g6902 = \DFF_414.D ;
  assign g6903 = \DFF_452.D ;
  assign g6904 = \DFF_18.D ;
  assign g6905 = \DFF_380.D ;
  assign g6906 = \DFF_176.D ;
  assign g6907 = \DFF_251.D ;
  assign g6908 = \DFF_428.D ;
  assign g6909 = \DFF_111.D ;
  assign g691 = \DFF_521.Q ;
  assign g6910 = \DFF_345.D ;
  assign g6911 = \DFF_197.D ;
  assign g6912 = \DFF_167.D ;
  assign g6913 = \DFF_473.D ;
  assign g6914 = \DFF_165.D ;
  assign g6915 = \DFF_390.D ;
  assign g6916 = \DFF_279.D ;
  assign g6918 = \DFF_108.D ;
  assign g6919 = g5816;
  assign g6921 = g6920;
  assign g6922 = \DFF_46.D ;
  assign g6923 = \DFF_511.D ;
  assign g6924 = \DFF_87.D ;
  assign g6925 = \DFF_494.D ;
  assign g6927 = g6926;
  assign g6928 = \DFF_133.D ;
  assign g6929 = \DFF_229.D ;
  assign g6930 = \DFF_115.D ;
  assign g6931 = \DFF_97.D ;
  assign g6933 = g6932;
  assign g6934 = \DFF_123.D ;
  assign g6938 = \DFF_315.D ;
  assign g6939 = \DFF_29.D ;
  assign g6943 = g6942;
  assign g6947 = \DFF_201.D ;
  assign g6948 = \DFF_24.D ;
  assign g695 = \DFF_11.Q ;
  assign g6950 = g6949;
  assign g6954 = \DFF_118.D ;
  assign g6956 = g6955;
  assign g6960 = \DFF_169.D ;
  assign g6970 = \DFF_90.D ;
  assign g6983 = \DFF_75.D ;
  assign g6993 = \DFF_528.D ;
  assign g7 = \DFF_445.Q ;
  assign g70 = \DFF_224.Q ;
  assign g700 = \DFF_281.Q ;
  assign g7007 = \DFF_296.D ;
  assign g7008 = \DFF_520.D ;
  assign g7009 = \DFF_140.D ;
  assign g7010 = \DFF_371.D ;
  assign g7020 = \DFF_17.D ;
  assign g7021 = \DFF_425.D ;
  assign g7023 = \DFF_392.D ;
  assign g7024 = \DFF_456.D ;
  assign g7026 = \DFF_20.D ;
  assign g7027 = \DFF_218.D ;
  assign g7029 = \DFF_254.D ;
  assign g7030 = \DFF_81.D ;
  assign g7032 = \DFF_4.D ;
  assign g7033 = \DFF_391.D ;
  assign g7034 = \DFF_466.D ;
  assign g7035 = \DFF_477.D ;
  assign g7037 = \DFF_400.D ;
  assign g7038 = \DFF_505.D ;
  assign g7039 = \DFF_453.D ;
  assign g704 = \DFF_57.Q ;
  assign g7040 = \DFF_138.D ;
  assign g7042 = \DFF_237.D ;
  assign g7043 = \DFF_164.D ;
  assign g7044 = \DFF_463.D ;
  assign g7047 = \DFF_42.D ;
  assign g7048 = \DFF_514.D ;
  assign g7049 = \DFF_141.D ;
  assign g7051 = \DFF_426.D ;
  assign g7052 = \DFF_10.D ;
  assign g7053 = g872;
  assign g7056 = \DFF_326.D ;
  assign g7057 = \DFF_256.D ;
  assign g7058 = g873;
  assign g7064 = \DFF_39.D ;
  assign g7065 = \DFF_130.D ;
  assign g7066 = \DFF_268.D ;
  assign g7069 = \DFF_258.D ;
  assign g7070 = \DFF_523.D ;
  assign g7072 = \DFF_332.D ;
  assign g7073 = \DFF_59.D ;
  assign g7076 = \DFF_49.D ;
  assign g7078 = \DFF_363.D ;
  assign g7082 = \DFF_397.D ;
  assign g7089 = \DFF_500.D ;
  assign g709 = \DFF_15.Q ;
  assign g7093 = \DFF_356.D ;
  assign g7097 = \DFF_531.D ;
  assign g7098 = \DFF_446.D ;
  assign g7103 = \DFF_193.D ;
  assign g7106 = \DFF_35.D ;
  assign g7107 = \DFF_443.D ;
  assign g7110 = \DFF_244.D ;
  assign g7113 = \DFF_222.D ;
  assign g7116 = \DFF_246.D ;
  assign g7119 = \DFF_270.D ;
  assign g7122 = \DFF_179.D ;
  assign g7126 = \DFF_71.D ;
  assign g713 = \DFF_6.Q ;
  assign g7133 = \DFF_103.D ;
  assign g7134 = \DFF_64.D ;
  assign g7137 = \DFF_403.D ;
  assign g7143 = \DFF_496.D ;
  assign g7144 = \DFF_336.D ;
  assign g7147 = \DFF_63.D ;
  assign g718 = \DFF_48.Q ;
  assign g7183 = \DFF_213.D ;
  assign g7187 = \DFF_91.D ;
  assign g7189 = \DFF_287.D ;
  assign g7191 = \DFF_247.D ;
  assign g7192 = g48;
  assign g7195 = \DFF_513.D ;
  assign g7202 = \DFF_184.D ;
  assign g7203 = \DFF_274.D ;
  assign g7204 = \DFF_479.D ;
  assign g7211 = \DFF_422.D ;
  assign g7212 = \DFF_224.D ;
  assign g7218 = \DFF_527.D ;
  assign g7219 = \DFF_533.D ;
  assign g722 = \DFF_286.Q ;
  assign g7225 = \DFF_236.D ;
  assign g7231 = \DFF_439.D ;
  assign g7236 = \DFF_110.D ;
  assign g7240 = \DFF_305.D ;
  assign g7242 = \DFF_348.D ;
  assign g7244 = \DFF_192.D ;
  assign g7245 = \DFF_298.D ;
  assign g7257 = \DFF_234.D ;
  assign g7258 = \DFF_160.D ;
  assign g727 = \DFF_427.Q ;
  assign g7284 = g27;
  assign g7285 = \DFF_71.D ;
  assign g7287 = \DFF_336.D ;
  assign g7288 = \DFF_253.D ;
  assign g7289 = \DFF_127.D ;
  assign g7290 = \DFF_32.D ;
  assign g7291 = \DFF_498.D ;
  assign g7292 = \DFF_61.D ;
  assign g7293 = \DFF_250.D ;
  assign g7294 = \DFF_486.D ;
  assign g7295 = \DFF_401.D ;
  assign g7296 = \DFF_510.D ;
  assign g7297 = \DFF_202.D ;
  assign g7298 = \DFF_334.D ;
  assign g7299 = \DFF_231.D ;
  assign g73 = \DFF_533.Q ;
  assign g7300 = \DFF_355.D ;
  assign g7301 = \DFF_442.D ;
  assign g7302 = \DFF_58.D ;
  assign g7303 = \DFF_322.D ;
  assign g7304 = \DFF_400.D ;
  assign g7305 = \DFF_88.D ;
  assign g7306 = \DFF_303.D ;
  assign g7307 = \DFF_142.D ;
  assign g7308 = \DFF_163.D ;
  assign g7309 = \DFF_132.D ;
  assign g731 = \DFF_359.Q ;
  assign g7310 = \DFF_125.D ;
  assign g7311 = \DFF_67.D ;
  assign g7312 = \DFF_327.D ;
  assign g7313 = \DFF_331.D ;
  assign g7314 = \DFF_487.D ;
  assign g7315 = \DFF_5.D ;
  assign g7316 = \DFF_189.D ;
  assign g7317 = \DFF_105.D ;
  assign g7318 = \DFF_396.D ;
  assign g7319 = \DFF_185.D ;
  assign g7320 = \DFF_452.D ;
  assign g7321 = \DFF_473.D ;
  assign g7322 = \DFF_153.D ;
  assign g7323 = \DFF_76.D ;
  assign g7324 = \DFF_182.D ;
  assign g7325 = \DFF_33.D ;
  assign g7326 = \DFF_237.D ;
  assign g7327 = \DFF_165.D ;
  assign g7328 = \DFF_97.D ;
  assign g7329 = \DFF_201.D ;
  assign g7330 = \DFF_24.D ;
  assign g7331 = \DFF_169.D ;
  assign g7332 = \DFF_90.D ;
  assign g7333 = \DFF_494.D ;
  assign g7334 = \DFF_315.D ;
  assign g7335 = \DFF_118.D ;
  assign g7336 = \DFF_179.D ;
  assign g7337 = \DFF_531.D ;
  assign g7338 = \DFF_391.D ;
  assign g7339 = \DFF_505.D ;
  assign g7340 = \DFF_164.D ;
  assign g7341 = \DFF_42.D ;
  assign g7342 = \DFF_426.D ;
  assign g7343 = \DFF_326.D ;
  assign g7344 = \DFF_39.D ;
  assign g7345 = \DFF_258.D ;
  assign g7346 = \DFF_453.D ;
  assign g7347 = \DFF_463.D ;
  assign g7348 = \DFF_514.D ;
  assign g7349 = \DFF_10.D ;
  assign g7350 = \DFF_256.D ;
  assign g7351 = \DFF_130.D ;
  assign g7352 = \DFF_520.D ;
  assign g7353 = \DFF_140.D ;
  assign g7354 = \DFF_17.D ;
  assign g7355 = \DFF_392.D ;
  assign g7356 = \DFF_20.D ;
  assign g7357 = \DFF_254.D ;
  assign g7358 = \DFF_466.D ;
  assign g7359 = \DFF_138.D ;
  assign g736 = \DFF_86.Q ;
  assign g7360 = \DFF_371.D ;
  assign g7361 = \DFF_425.D ;
  assign g7362 = \DFF_456.D ;
  assign g7363 = \DFF_218.D ;
  assign g7364 = \DFF_81.D ;
  assign g7365 = \DFF_477.D ;
  assign g7366 = \DFF_385.D ;
  assign g7369 = g42;
  assign g7374 = \DFF_4.D ;
  assign g7376 = \DFF_247.D ;
  assign g7377 = \DFF_192.D ;
  assign g7380 = g43;
  assign g7387 = \DFF_184.D ;
  assign g7388 = \DFF_234.D ;
  assign g7390 = g44;
  assign g7395 = g45;
  assign g7415 = \DFF_30.D ;
  assign g7421 = \DFF_393.D ;
  assign g7441 = \DFF_518.D ;
  assign g7445 = \DFF_289.D ;
  assign g7446 = g82;
  assign g745 = \DFF_89.Q ;
  assign g7450 = g82;
  assign g7454 = g82;
  assign g746 = \DFF_304.Q ;
  assign g7460 = g82;
  assign g7464 = \DFF_220.D ;
  assign g7467 = g82;
  assign g7473 = g82;
  assign g7477 = \DFF_413.D ;
  assign g7497 = g82;
  assign g7501 = \DFF_307.D ;
  assign g7502 = \DFF_515.D ;
  assign g7505 = g82;
  assign g7509 = \DFF_497.D ;
  assign g7512 = g82;
  assign g7516 = g82;
  assign g7520 = \DFF_364.D ;
  assign g7521 = \DFF_386.D ;
  assign g7522 = \DFF_414.D ;
  assign g7525 = \DFF_18.D ;
  assign g7527 = g82;
  assign g7530 = \DFF_485.D ;
  assign g7531 = \DFF_259.D ;
  assign g7532 = \DFF_428.D ;
  assign g7534 = \DFF_111.D ;
  assign g7537 = \DFF_380.D ;
  assign g7538 = \DFF_176.D ;
  assign g7539 = \DFF_251.D ;
  assign g754 = \DFF_431.Q ;
  assign g7540 = \DFF_167.D ;
  assign g7541 = \DFF_324.D ;
  assign g7543 = g872;
  assign g7544 = \DFF_345.D ;
  assign g7545 = \DFF_197.D ;
  assign g7546 = \DFF_108.D ;
  assign g755 = \DFF_462.Q ;
  assign g7550 = g42;
  assign g7555 = g5816;
  assign g7556 = g873;
  assign g7559 = \DFF_390.D ;
  assign g756 = \DFF_156.Q ;
  assign g7560 = \DFF_279.D ;
  assign g7561 = \DFF_87.D ;
  assign g7562 = g43;
  assign g7568 = \DFF_270.D ;
  assign g7569 = \DFF_46.D ;
  assign g757 = \DFF_37.Q ;
  assign g7570 = \DFF_511.D ;
  assign g7571 = \DFF_115.D ;
  assign g7574 = g44;
  assign g7579 = \DFF_133.D ;
  assign g758 = \DFF_112.Q ;
  assign g7580 = \DFF_229.D ;
  assign g7581 = \DFF_418.D ;
  assign g7585 = \DFF_123.D ;
  assign g7586 = \DFF_119.D ;
  assign g7589 = \DFF_160.D ;
  assign g7590 = \DFF_28.D ;
  assign g7594 = \DFF_35.D ;
  assign g76 = \DFF_49.Q ;
  assign g7608 = \DFF_29.D ;
  assign g7611 = \DFF_296.D ;
  assign g7618 = \DFF_75.D ;
  assign g7619 = \DFF_528.D ;
  assign g762 = \DFF_407.Q ;
  assign g7626 = \DFF_72.D ;
  assign g7627 = \DFF_141.D ;
  assign g7628 = \DFF_268.D ;
  assign g7629 = \DFF_523.D ;
  assign g7630 = \DFF_332.D ;
  assign g7631 = \DFF_397.D ;
  assign g7632 = \DFF_361.D ;
  assign g7633 = \DFF_59.D ;
  assign g7634 = \DFF_500.D ;
  assign g7635 = \DFF_356.D ;
  assign g7636 = \DFF_446.D ;
  assign g7637 = \DFF_49.D ;
  assign g7648 = \DFF_274.D ;
  assign g7649 = \DFF_193.D ;
  assign g7650 = \DFF_363.D ;
  assign g7656 = \DFF_422.D ;
  assign g7657 = \DFF_443.D ;
  assign g7658 = \DFF_527.D ;
  assign g7659 = \DFF_244.D ;
  assign g766 = \DFF_149.Q ;
  assign g7660 = \DFF_196.D ;
  assign g7662 = \DFF_236.D ;
  assign g7663 = \DFF_222.D ;
  assign g7669 = \DFF_439.D ;
  assign g7672 = \DFF_246.D ;
  assign g7673 = \DFF_110.D ;
  assign g7675 = \DFF_305.D ;
  assign g7676 = \DFF_348.D ;
  assign g7677 = g82;
  assign g7678 = \DFF_298.D ;
  assign g7680 = g82;
  assign g7681 = g82;
  assign g7682 = g82;
  assign g7683 = g82;
  assign g7684 = g82;
  assign g7685 = g82;
  assign g7686 = g82;
  assign g7688 = g82;
  assign g7692 = g82;
  assign g7696 = g82;
  assign g770 = \DFF_253.Q ;
  assign g7705 = \DFF_301.D ;
  assign g7706 = \DFF_103.D ;
  assign g7709 = \DFF_387.D ;
  assign g7723 = \DFF_496.D ;
  assign g7724 = \DFF_63.D ;
  assign g7725 = \DFF_213.D ;
  assign g7726 = \DFF_91.D ;
  assign g7727 = \DFF_64.D ;
  assign g7728 = \DFF_287.D ;
  assign g7729 = \DFF_403.D ;
  assign g7731 = \DFF_513.D ;
  assign g7733 = \DFF_479.D ;
  assign g7735 = \DFF_224.D ;
  assign g7737 = \DFF_533.D ;
  assign g774 = \DFF_30.Q ;
  assign g7744 = g27;
  assign g7745 = \DFF_380.D ;
  assign g7746 = \DFF_296.D ;
  assign g7747 = \DFF_220.D ;
  assign g7748 = \DFF_307.D ;
  assign g7749 = \DFF_364.D ;
  assign g7750 = \DFF_397.D ;
  assign g7751 = \DFF_270.D ;
  assign g7752 = \DFF_500.D ;
  assign g7753 = \DFF_356.D ;
  assign g7754 = \DFF_446.D ;
  assign g7755 = \DFF_193.D ;
  assign g7756 = \DFF_443.D ;
  assign g7757 = \DFF_244.D ;
  assign g7758 = \DFF_222.D ;
  assign g7759 = \DFF_246.D ;
  assign g7760 = \DFF_386.D ;
  assign g7761 = \DFF_485.D ;
  assign g7762 = \DFF_176.D ;
  assign g7763 = \DFF_345.D ;
  assign g7764 = \DFF_390.D ;
  assign g7765 = \DFF_46.D ;
  assign g7766 = \DFF_133.D ;
  assign g7767 = \DFF_123.D ;
  assign g7768 = \DFF_259.D ;
  assign g7769 = \DFF_251.D ;
  assign g7770 = \DFF_197.D ;
  assign g7771 = \DFF_279.D ;
  assign g7772 = \DFF_511.D ;
  assign g7773 = \DFF_229.D ;
  assign g7774 = \DFF_496.D ;
  assign g7775 = \DFF_49.D ;
  assign g7776 = \DFF_363.D ;
  assign g7777 = \DFF_63.D ;
  assign g7778 = \DFF_213.D ;
  assign g7779 = \DFF_91.D ;
  assign g778 = \DFF_247.Q ;
  assign g7780 = \DFF_287.D ;
  assign g7781 = \DFF_513.D ;
  assign g7782 = \DFF_479.D ;
  assign g7783 = \DFF_224.D ;
  assign g7784 = \DFF_533.D ;
  assign g7785 = \DFF_30.D ;
  assign g7786 = \DFF_393.D ;
  assign g7787 = \DFF_274.D ;
  assign g7788 = \DFF_160.D ;
  assign g7789 = \DFF_35.D ;
  assign g7790 = \DFF_422.D ;
  assign g7791 = \DFF_527.D ;
  assign g7792 = \DFF_236.D ;
  assign g7793 = \DFF_439.D ;
  assign g7794 = \DFF_110.D ;
  assign g7795 = \DFF_305.D ;
  assign g7796 = \DFF_348.D ;
  assign g7797 = \DFF_298.D ;
  assign g7798 = \DFF_413.D ;
  assign g7799 = \DFF_192.D ;
  assign g7800 = \DFF_234.D ;
  assign g7801 = \DFF_515.D ;
  assign g7802 = \DFF_497.D ;
  assign g7803 = \DFF_414.D ;
  assign g7804 = \DFF_428.D ;
  assign g7805 = \DFF_167.D ;
  assign g7806 = \DFF_108.D ;
  assign g7807 = \DFF_87.D ;
  assign g7808 = \DFF_115.D ;
  assign g7809 = \DFF_289.D ;
  assign g7810 = \DFF_103.D ;
  assign g7811 = \DFF_268.D ;
  assign g7812 = \DFF_523.D ;
  assign g7813 = \DFF_332.D ;
  assign g7814 = \DFF_59.D ;
  assign g7815 = \DFF_141.D ;
  assign g7816 = \DFF_18.D ;
  assign g7817 = \DFF_111.D ;
  assign g782 = \DFF_301.Q ;
  assign g7843 = \DFF_147.D ;
  assign g7844 = \DFF_301.D ;
  assign g7845 = \DFF_64.D ;
  assign g7848 = \DFF_387.D ;
  assign g7849 = \DFF_403.D ;
  assign g786 = \DFF_38.Q ;
  assign g7896 = \DFF_247.D ;
  assign g7899 = \DFF_184.D ;
  assign g79 = \DFF_363.Q ;
  assign g790 = \DFF_434.Q ;
  assign g7904 = g5816;
  assign g7906 = \DFF_4.D ;
  assign g7921 = g6920;
  assign g7922 = \DFF_518.D ;
  assign g7924 = g6926;
  assign g7925 = g6932;
  assign g7927 = g6942;
  assign g7928 = g6949;
  assign g7929 = g6955;
  assign g7930 = \DFF_104.D ;
  assign g794 = \DFF_227.Q ;
  assign g7959 = \DFF_72.D ;
  assign g7966 = \DFF_324.D ;
  assign g7975 = \DFF_418.D ;
  assign g7976 = \DFF_119.D ;
  assign g7977 = \DFF_29.D ;
  assign g7979 = \DFF_28.D ;
  assign g798 = \DFF_429.Q ;
  assign g7981 = \DFF_269.D ;
  assign g7982 = \DFF_75.D ;
  assign g7983 = \DFF_528.D ;
  assign g7984 = g872;
  assign g7985 = g873;
  assign g7989 = g82;
  assign g7991 = g82;
  assign g7993 = g82;
  assign g7995 = g82;
  assign g7998 = g82;
  assign g7999 = g82;
  assign g8 = \DFF_267.Q ;
  assign g8001 = g82;
  assign g8002 = g82;
  assign g8003 = \DFF_196.D ;
  assign g8004 = g82;
  assign g8007 = g82;
  assign g8008 = g82;
  assign g8009 = \DFF_361.D ;
  assign g8019 = \DFF_38.D ;
  assign g802 = \DFF_389.Q ;
  assign g8024 = \DFF_99.D ;
  assign g8039 = \DFF_172.D ;
  assign g8040 = \DFF_273.D ;
  assign g8041 = \DFF_34.D ;
  assign g8042 = \DFF_306.D ;
  assign g8043 = \DFF_277.D ;
  assign g8044 = \DFF_508.D ;
  assign g8045 = \DFF_139.D ;
  assign g8046 = \DFF_95.D ;
  assign g8047 = \DFF_314.D ;
  assign g8048 = \DFF_337.D ;
  assign g8049 = \DFF_382.D ;
  assign g8050 = \DFF_102.D ;
  assign g8051 = \DFF_98.D ;
  assign g8052 = \DFF_437.D ;
  assign g8053 = \DFF_474.D ;
  assign g8054 = \DFF_490.D ;
  assign g8055 = \DFF_519.D ;
  assign g8059 = \DFF_444.D ;
  assign g806 = \DFF_127.Q ;
  assign g8060 = \DFF_190.D ;
  assign g8061 = g872;
  assign g8062 = g873;
  assign g8063 = \DFF_72.D ;
  assign g8064 = \DFF_518.D ;
  assign g8065 = \DFF_64.D ;
  assign g8066 = \DFF_403.D ;
  assign g8067 = \DFF_196.D ;
  assign g8076 = \DFF_247.D ;
  assign g8077 = \DFF_184.D ;
  assign g8078 = \DFF_528.D ;
  assign g8079 = \DFF_29.D ;
  assign g8080 = \DFF_75.D ;
  assign g8093 = \DFF_38.D ;
  assign g8096 = \DFF_99.D ;
  assign g810 = \DFF_393.Q ;
  assign g8116 = \DFF_172.D ;
  assign g8121 = \DFF_273.D ;
  assign g8122 = \DFF_34.D ;
  assign g8125 = \DFF_306.D ;
  assign g8126 = \DFF_277.D ;
  assign g8128 = \DFF_508.D ;
  assign g8132 = \DFF_301.D ;
  assign g8133 = \DFF_139.D ;
  assign g8134 = \DFF_95.D ;
  assign g8137 = \DFF_314.D ;
  assign g8138 = \DFF_337.D ;
  assign g814 = \DFF_184.Q ;
  assign g8140 = \DFF_387.D ;
  assign g8141 = \DFF_382.D ;
  assign g8142 = \DFF_102.D ;
  assign g8144 = \DFF_98.D ;
  assign g8145 = \DFF_437.D ;
  assign g8147 = \DFF_243.D ;
  assign g8149 = \DFF_474.D ;
  assign g8150 = \DFF_490.D ;
  assign g8152 = \DFF_519.D ;
  assign g8155 = \DFF_444.D ;
  assign g8156 = \DFF_190.D ;
  assign g8160 = \DFF_147.D ;
  assign g8164 = g41;
  assign g8171 = \DFF_4.D ;
  assign g8173 = \DFF_346.D ;
  assign g8178 = g6920;
  assign g8179 = g6926;
  assign g818 = \DFF_387.Q ;
  assign g8181 = g6932;
  assign g8182 = g6942;
  assign g8183 = g6949;
  assign g8184 = g6955;
  assign g8186 = \DFF_269.D ;
  assign g8187 = g8352;
  assign g8191 = \DFF_104.D ;
  assign g8192 = g5816;
  assign g8193 = \DFF_74.D ;
  assign g8194 = \DFF_435.D ;
  assign g8195 = \DFF_324.D ;
  assign g8196 = \DFF_418.D ;
  assign g8197 = \DFF_119.D ;
  assign g8198 = \DFF_28.D ;
  assign g8200 = g8347;
  assign g8203 = g8313;
  assign g8206 = g8316;
  assign g8210 = g8318;
  assign g8214 = g8323;
  assign g822 = \DFF_99.Q ;
  assign g8221 = g8328;
  assign g8226 = g8331;
  assign g8230 = g8335;
  assign g8233 = g41;
  assign g8236 = g8340;
  assign g8241 = g8349;
  assign g8244 = \DFF_434.D ;
  assign g8245 = \DFF_347.D ;
  assign g8250 = \DFF_83.D ;
  assign g8251 = \DFF_361.D ;
  assign g8254 = \DFF_340.D ;
  assign g826 = \DFF_347.Q ;
  assign g8260 = \DFF_13.D ;
  assign g8271 = g5816;
  assign g8272 = \DFF_4.D ;
  assign g8273 = \DFF_301.D ;
  assign g8274 = \DFF_387.D ;
  assign g8275 = \DFF_269.D ;
  assign g8276 = \DFF_361.D ;
  assign g8277 = \DFF_418.D ;
  assign g8278 = \DFF_119.D ;
  assign g8279 = \DFF_28.D ;
  assign g8280 = \DFF_324.D ;
  assign g8281 = \DFF_349.D ;
  assign g8282 = \DFF_85.D ;
  assign g8283 = \DFF_493.D ;
  assign g8284 = \DFF_209.D ;
  assign g8285 = \DFF_339.D ;
  assign g8286 = \DFF_373.D ;
  assign g8287 = \DFF_313.D ;
  assign g8288 = \DFF_155.D ;
  assign g829 = \DFF_55.Q ;
  assign g8292 = \DFF_434.D ;
  assign g8294 = \DFF_347.D ;
  assign g8304 = \DFF_83.D ;
  assign g8306 = \DFF_340.D ;
  assign g8310 = \DFF_13.D ;
  assign g8311 = \DFF_38.D ;
  assign g8312 = \DFF_99.D ;
  assign g8314 = g8313;
  assign g8315 = \DFF_172.D ;
  assign g8317 = g8316;
  assign g8319 = g8318;
  assign g8320 = \DFF_273.D ;
  assign g8321 = \DFF_34.D ;
  assign g8324 = g8323;
  assign g8325 = \DFF_306.D ;
  assign g8326 = \DFF_277.D ;
  assign g8329 = g8328;
  assign g833 = \DFF_338.Q ;
  assign g8330 = \DFF_508.D ;
  assign g8332 = g8331;
  assign g8333 = \DFF_139.D ;
  assign g8334 = \DFF_95.D ;
  assign g8336 = g8335;
  assign g8337 = g6920;
  assign g8338 = \DFF_314.D ;
  assign g8339 = \DFF_337.D ;
  assign g8341 = g8340;
  assign g8342 = g6926;
  assign g8343 = \DFF_382.D ;
  assign g8344 = \DFF_102.D ;
  assign g8345 = \DFF_98.D ;
  assign g8346 = \DFF_437.D ;
  assign g8348 = g8347;
  assign g8350 = g8349;
  assign g8351 = g6932;
  assign g8353 = g8352;
  assign g8354 = g6942;
  assign g8355 = \DFF_474.D ;
  assign g8356 = \DFF_490.D ;
  assign g8357 = \DFF_519.D ;
  assign g8358 = g6949;
  assign g8359 = g6955;
  assign g8360 = \DFF_444.D ;
  assign g8361 = \DFF_190.D ;
  assign g8362 = \DFF_147.D ;
  assign g8363 = \DFF_243.D ;
  assign g837 = \DFF_309.Q ;
  assign g8375 = \DFF_346.D ;
  assign g8376 = \DFF_104.D ;
  assign g8378 = \DFF_74.D ;
  assign g8379 = \DFF_435.D ;
  assign g8381 = g41;
  assign g8384 = \DFF_223.D ;
  assign g841 = \DFF_412.Q ;
  assign g8418 = \DFF_382.D ;
  assign g8419 = \DFF_474.D ;
  assign g8420 = \DFF_444.D ;
  assign g8421 = \DFF_508.D ;
  assign g8422 = \DFF_314.D ;
  assign g8423 = \DFF_102.D ;
  assign g8424 = \DFF_490.D ;
  assign g8425 = \DFF_190.D ;
  assign g8426 = \DFF_147.D ;
  assign g8427 = \DFF_337.D ;
  assign g8428 = \DFF_488.D ;
  assign g8429 = \DFF_60.D ;
  assign g8430 = \DFF_521.D ;
  assign g8431 = \DFF_281.D ;
  assign g8432 = \DFF_15.D ;
  assign g8433 = \DFF_48.D ;
  assign g8434 = \DFF_427.D ;
  assign g8435 = \DFF_86.D ;
  assign g8436 = \DFF_38.D ;
  assign g8437 = \DFF_99.D ;
  assign g8438 = \DFF_306.D ;
  assign g8439 = \DFF_139.D ;
  assign g8440 = \DFF_98.D ;
  assign g8441 = \DFF_172.D ;
  assign g8442 = \DFF_273.D ;
  assign g8443 = \DFF_277.D ;
  assign g8444 = \DFF_95.D ;
  assign g8445 = \DFF_437.D ;
  assign g8446 = \DFF_519.D ;
  assign g8447 = \DFF_34.D ;
  assign g8448 = \DFF_74.D ;
  assign g8449 = \DFF_435.D ;
  assign g845 = \DFF_433.Q ;
  assign g8450 = \DFF_104.D ;
  assign g8472 = \DFF_434.D ;
  assign g8473 = \DFF_347.D ;
  assign g8476 = \DFF_83.D ;
  assign g8478 = \DFF_340.D ;
  assign g8480 = \DFF_13.D ;
  assign g849 = \DFF_343.Q ;
  assign g8500 = \DFF_243.D ;
  assign g8505 = \DFF_261.D ;
  assign g8513 = g6920;
  assign g8514 = g6926;
  assign g8515 = g6932;
  assign g8516 = g6942;
  assign g8517 = g6949;
  assign g8518 = g6955;
  assign g8519 = \DFF_346.D ;
  assign g853 = \DFF_405.Q ;
  assign g8559 = \DFF_532.D ;
  assign g8560 = \DFF_223.D ;
  assign g8561 = g6920;
  assign g8562 = g6926;
  assign g8563 = g6932;
  assign g8564 = g6942;
  assign g8565 = g6949;
  assign g8566 = g6955;
  assign g8567 = \DFF_434.D ;
  assign g8568 = \DFF_347.D ;
  assign g8569 = \DFF_243.D ;
  assign g857 = \DFF_367.Q ;
  assign g8570 = \DFF_83.D ;
  assign g8571 = \DFF_340.D ;
  assign g8572 = \DFF_13.D ;
  assign g8573 = \DFF_346.D ;
  assign g8575 = \DFF_532.D ;
  assign g8588 = \DFF_223.D ;
  assign g8600 = g8313;
  assign g8601 = g8316;
  assign g8604 = g8318;
  assign g8606 = g8323;
  assign g8608 = g8328;
  assign g861 = \DFF_248.Q ;
  assign g8610 = g8331;
  assign g8613 = g8335;
  assign g8622 = g8340;
  assign g8624 = g8347;
  assign g8625 = g8349;
  assign g8626 = g8352;
  assign g8631 = \DFF_360.D ;
  assign g8649 = \DFF_180.D ;
  assign g865 = \DFF_269.Q ;
  assign g8650 = \DFF_261.D ;
  assign g868 = \DFF_441.Q ;
  assign g869 = \DFF_188.Q ;
  assign g8694 = \DFF_223.D ;
  assign g8695 = \DFF_532.D ;
  assign g8714 = \DFF_360.D ;
  assign g874 = \DFF_357.Q ;
  assign g8747 = \DFF_180.D ;
  assign g875 = \DFF_398.Q ;
  assign g8758 = \DFF_261.D ;
  assign g876 = \DFF_93.Q ;
  assign g8765 = \DFF_415.D ;
  assign g8766 = \DFF_36.D ;
  assign g8767 = \DFF_128.D ;
  assign g8768 = \DFF_503.D ;
  assign g8769 = \DFF_109.D ;
  assign g8770 = \DFF_482.D ;
  assign g8771 = \DFF_516.D ;
  assign g8772 = \DFF_47.D ;
  assign g8773 = \DFF_374.D ;
  assign g8774 = \DFF_249.D ;
  assign g8775 = \DFF_235.D ;
  assign g8776 = \DFF_495.D ;
  assign g8777 = \DFF_199.D ;
  assign g8779 = \DFF_404.D ;
  assign g878 = \DFF_53.Q ;
  assign g8780 = \DFF_261.D ;
  assign g8781 = \DFF_360.D ;
  assign g8782 = \DFF_180.D ;
  assign g8784 = \DFF_482.D ;
  assign g8785 = \DFF_516.D ;
  assign g8788 = \DFF_374.D ;
  assign g8790 = \DFF_249.D ;
  assign g8792 = \DFF_495.D ;
  assign g8794 = \DFF_415.D ;
  assign g8795 = \DFF_199.D ;
  assign g8797 = \DFF_36.D ;
  assign g8798 = \DFF_404.D ;
  assign g8800 = \DFF_128.D ;
  assign g8802 = \DFF_503.D ;
  assign g8803 = \DFF_109.D ;
  assign g8804 = \DFF_47.D ;
  assign g8805 = \DFF_235.D ;
  assign g8806 = g8977;
  assign g8810 = g8978;
  assign g8811 = g8979;
  assign g8812 = g8980;
  assign g8813 = g8981;
  assign g8814 = g8982;
  assign g8815 = g8983;
  assign g8816 = g8984;
  assign g8817 = g8976;
  assign g8818 = g8985;
  assign g8819 = g8986;
  assign g882 = \DFF_121.Q ;
  assign g8820 = \DFF_43.D ;
  assign g883 = \DFF_291.Q ;
  assign g8868 = \DFF_482.D ;
  assign g8869 = \DFF_516.D ;
  assign g8870 = \DFF_374.D ;
  assign g8871 = \DFF_249.D ;
  assign g8872 = \DFF_495.D ;
  assign g8873 = \DFF_199.D ;
  assign g8874 = \DFF_404.D ;
  assign g8883 = \DFF_450.D ;
  assign g8884 = \DFF_415.D ;
  assign g8885 = \DFF_316.D ;
  assign g8886 = \DFF_36.D ;
  assign g8887 = \DFF_11.D ;
  assign g8888 = \DFF_128.D ;
  assign g8889 = \DFF_57.D ;
  assign g8890 = \DFF_503.D ;
  assign g8891 = \DFF_109.D ;
  assign g8920 = \DFF_6.D ;
  assign g8921 = \DFF_449.D ;
  assign g8922 = \DFF_381.D ;
  assign g8923 = \DFF_286.D ;
  assign g8924 = \DFF_47.D ;
  assign g8926 = \DFF_359.D ;
  assign g8928 = \DFF_235.D ;
  assign g8937 = \DFF_354.D ;
  assign g8938 = \DFF_333.D ;
  assign g8939 = \DFF_461.D ;
  assign g8940 = \DFF_300.D ;
  assign g8941 = \DFF_44.D ;
  assign g8943 = \DFF_1.D ;
  assign g8944 = \DFF_212.D ;
  assign g8945 = \DFF_271.D ;
  assign g8946 = g8977;
  assign g8948 = g8978;
  assign g8950 = g8979;
  assign g8951 = g8980;
  assign g8952 = g8981;
  assign g8953 = g8982;
  assign g8954 = g8983;
  assign g8956 = g8984;
  assign g8958 = g8976;
  assign g8959 = g8985;
  assign g8961 = g8986;
  assign g8969 = \DFF_43.D ;
  assign g8973 = \DFF_395.D ;
  assign g8987 = \DFF_36.D ;
  assign g8988 = \DFF_503.D ;
  assign g8989 = \DFF_47.D ;
  assign g8990 = \DFF_235.D ;
  assign g8991 = \DFF_415.D ;
  assign g8992 = \DFF_128.D ;
  assign g8993 = \DFF_109.D ;
  assign g9 = \DFF_179.Q ;
  assign g9009 = \DFF_354.D ;
  assign g9024 = \DFF_333.D ;
  assign g9025 = \DFF_461.D ;
  assign g9026 = \DFF_300.D ;
  assign g9027 = \DFF_44.D ;
  assign g9028 = \DFF_212.D ;
  assign g9029 = \DFF_271.D ;
  assign g9088 = g9451;
  assign g9106 = \DFF_43.D ;
  assign g9108 = \DFF_395.D ;
  assign g9109 = \DFF_381.D ;
  assign g9110 = \DFF_358.D ;
  assign g9124 = \DFF_310.D ;
  assign g9150 = \DFF_362.D ;
  assign g9262 = \DFF_449.D ;
  assign g9264 = \DFF_1.D ;
  assign g9266 = \DFF_297.D ;
  assign g9269 = \DFF_302.D ;
  assign g9270 = \DFF_450.D ;
  assign g9272 = \DFF_369.D ;
  assign g9273 = \DFF_316.D ;
  assign g928 = \DFF_243.Q ;
  assign g9290 = \DFF_11.D ;
  assign g9308 = \DFF_57.D ;
  assign g9310 = \DFF_6.D ;
  assign g9311 = \DFF_286.D ;
  assign g9312 = \DFF_359.D ;
  assign g932 = \DFF_83.Q ;
  assign g9338 = \DFF_43.D ;
  assign g9339 = \DFF_395.D ;
  assign g9340 = \DFF_381.D ;
  assign g9341 = \DFF_450.D ;
  assign g9342 = \DFF_316.D ;
  assign g9343 = \DFF_11.D ;
  assign g9344 = \DFF_57.D ;
  assign g9345 = \DFF_6.D ;
  assign g9346 = \DFF_286.D ;
  assign g9347 = \DFF_359.D ;
  assign g9348 = \DFF_449.D ;
  assign g9349 = \DFF_1.D ;
  assign g9350 = \DFF_354.D ;
  assign g9351 = \DFF_333.D ;
  assign g9352 = \DFF_461.D ;
  assign g9353 = \DFF_300.D ;
  assign g9354 = \DFF_44.D ;
  assign g9355 = \DFF_212.D ;
  assign g9356 = \DFF_271.D ;
  assign g936 = \DFF_340.Q ;
  assign g9360 = \DFF_369.D ;
  assign g940 = \DFF_13.Q ;
  assign g944 = \DFF_312.Q ;
  assign g9452 = g9451;
  assign g947 = \DFF_454.Q ;
  assign g950 = \DFF_365.Q ;
  assign g9507 = \DFF_357.D ;
  assign g9508 = \DFF_398.D ;
  assign g9525 = \DFF_137.D ;
  assign g9526 = \DFF_526.D ;
  assign g953 = \DFF_317.Q ;
  assign g9532 = \DFF_358.D ;
  assign g9533 = \DFF_310.D ;
  assign g9535 = \DFF_362.D ;
  assign g9555 = \DFF_455.D ;
  assign g956 = \DFF_408.Q ;
  assign g959 = \DFF_106.Q ;
  assign g962 = \DFF_148.Q ;
  assign g965 = \DFF_181.Q ;
  assign g9661 = \DFF_297.D ;
  assign g9666 = \DFF_302.D ;
  assign g9670 = \DFF_297.D ;
  assign g9671 = \DFF_302.D ;
  assign g9672 = \DFF_369.D ;
  assign g968 = \DFF_351.Q ;
  assign g97 = g872;
  assign g971 = \DFF_294.Q ;
  assign g9721 = \DFF_135.D ;
  assign g9732 = \DFF_137.D ;
  assign g9733 = \DFF_526.D ;
  assign g976 = \DFF_14.Q ;
  assign g9762 = \DFF_357.D ;
  assign g9763 = \DFF_398.D ;
  assign g9765 = \DFF_358.D ;
  assign g9767 = \DFF_310.D ;
  assign g9769 = \DFF_362.D ;
  assign g98 = g873;
  assign g981 = \DFF_52.Q ;
  assign g9813 = \DFF_455.D ;
  assign g9818 = \DFF_358.D ;
  assign g9819 = \DFF_310.D ;
  assign g9820 = \DFF_362.D ;
  assign g9821 = \DFF_357.D ;
  assign g9822 = \DFF_398.D ;
  assign g9823 = \DFF_137.D ;
  assign g9824 = \DFF_526.D ;
  assign g9825 = \DFF_297.D ;
  assign g9826 = \DFF_302.D ;
  assign g9827 = \DFF_369.D ;
  assign g9832 = \DFF_455.D ;
  assign g9845 = g9451;
  assign g986 = \DFF_293.Q ;
  assign g9875 = \DFF_135.D ;
  assign g9895 = \DFF_455.D ;
  assign g991 = \DFF_497.Q ;
  assign g9919 = \DFF_135.D ;
  assign g9930 = \DFF_135.D ;
  assign g9931 = g9961;
  assign g995 = \DFF_515.Q ;
  assign g9958 = g9961;
  assign g999 = \DFF_428.Q ;
endmodule
