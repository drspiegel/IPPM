
module s832(GND, VDD, CK, G0, G1, G10, G11, G12, G13, G14, G15, G16, G18, G2, G288, G290, G292, G296, G298, G3, G300, G302, G310, G312, G315, G322, G325, G327, G4, G43, G45, G47, G49, G5, G53, G55, G6, G7, G8, G9);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  input CK;
  wire \DFF_0.CK ;
  wire \DFF_0.D ;
  wire \DFF_0.Q ;
  wire \DFF_1.CK ;
  wire \DFF_1.D ;
  wire \DFF_1.Q ;
  wire \DFF_2.CK ;
  wire \DFF_2.D ;
  wire \DFF_2.Q ;
  wire \DFF_3.CK ;
  wire \DFF_3.D ;
  wire \DFF_3.Q ;
  wire \DFF_4.CK ;
  wire \DFF_4.D ;
  wire \DFF_4.Q ;
  input G0;
  input G1;
  input G10;
  wire G102;
  input G11;
  input G12;
  input G13;
  input G14;
  input G15;
  input G16;
  input G18;
  input G2;
  output G288;
  output G290;
  output G292;
  output G296;
  output G298;
  input G3;
  output G300;
  output G302;
  output G310;
  output G312;
  output G315;
  output G322;
  output G325;
  output G327;
  wire G38;
  wire G39;
  input G4;
  wire G40;
  wire G41;
  wire G42;
  output G43;
  output G45;
  output G47;
  output G49;
  input G5;
  output G53;
  output G55;
  input G6;
  input G7;
  input G8;
  input G9;
  wire G90;
  wire G93;
  wire G96;
  wire G99;
  input GND;
  input VDD;
  al_inv _133_ (
    .a(G4),
    .y(_095_)
  );
  al_inv _134_ (
    .a(G16),
    .y(_096_)
  );
  al_nand3ftt _135_ (
    .a(\DFF_0.Q ),
    .b(\DFF_3.Q ),
    .c(\DFF_4.Q ),
    .y(_097_)
  );
  al_nand3 _136_ (
    .a(\DFF_3.Q ),
    .b(\DFF_2.Q ),
    .c(\DFF_4.Q ),
    .y(_098_)
  );
  al_aoi21 _137_ (
    .a(_097_),
    .b(_098_),
    .c(\DFF_1.Q ),
    .y(_099_)
  );
  al_or2 _138_ (
    .a(\DFF_0.Q ),
    .b(\DFF_1.Q ),
    .y(_100_)
  );
  al_ao21ftt _139_ (
    .a(_100_),
    .b(\DFF_2.Q ),
    .c(_099_),
    .y(_101_)
  );
  al_ao21ftf _140_ (
    .a(_096_),
    .b(_095_),
    .c(_101_),
    .y(_102_)
  );
  al_and3fft _141_ (
    .a(\DFF_3.Q ),
    .b(\DFF_4.Q ),
    .c(\DFF_0.Q ),
    .y(_103_)
  );
  al_nand2 _142_ (
    .a(G4),
    .b(\DFF_1.Q ),
    .y(_104_)
  );
  al_oai21ftf _143_ (
    .a(\DFF_2.Q ),
    .b(_103_),
    .c(_104_),
    .y(_105_)
  );
  al_aoi21 _144_ (
    .a(\DFF_3.Q ),
    .b(\DFF_4.Q ),
    .c(G16),
    .y(_106_)
  );
  al_nand3ftt _145_ (
    .a(\DFF_2.Q ),
    .b(\DFF_1.Q ),
    .c(_106_),
    .y(_107_)
  );
  al_or3 _146_ (
    .a(\DFF_2.Q ),
    .b(\DFF_1.Q ),
    .c(\DFF_4.Q ),
    .y(_108_)
  );
  al_nor2 _147_ (
    .a(\DFF_0.Q ),
    .b(\DFF_3.Q ),
    .y(_109_)
  );
  al_and3ftt _148_ (
    .a(G1),
    .b(G16),
    .c(_109_),
    .y(_110_)
  );
  al_aoi21ftf _149_ (
    .a(_108_),
    .b(_110_),
    .c(_107_),
    .y(_111_)
  );
  al_nand3 _150_ (
    .a(_105_),
    .b(_111_),
    .c(_102_),
    .y(G302)
  );
  al_nand2 _151_ (
    .a(\DFF_3.Q ),
    .b(\DFF_4.Q ),
    .y(_112_)
  );
  al_and3ftt _152_ (
    .a(\DFF_0.Q ),
    .b(\DFF_2.Q ),
    .c(\DFF_1.Q ),
    .y(_113_)
  );
  al_or3 _153_ (
    .a(\DFF_0.Q ),
    .b(\DFF_3.Q ),
    .c(_108_),
    .y(_114_)
  );
  al_ao21ftf _154_ (
    .a(_112_),
    .b(_113_),
    .c(_114_),
    .y(G315)
  );
  al_and3fft _155_ (
    .a(\DFF_0.Q ),
    .b(_108_),
    .c(\DFF_3.Q ),
    .y(G53)
  );
  al_and2 _156_ (
    .a(G15),
    .b(G53),
    .y(G43)
  );
  al_nand3ftt _157_ (
    .a(\DFF_4.Q ),
    .b(\DFF_3.Q ),
    .c(\DFF_2.Q ),
    .y(_115_)
  );
  al_nor3fft _158_ (
    .a(G15),
    .b(G16),
    .c(_100_),
    .y(_116_)
  );
  al_ao21 _159_ (
    .a(G12),
    .b(G10),
    .c(G11),
    .y(_117_)
  );
  al_nand3ftt _160_ (
    .a(_115_),
    .b(_117_),
    .c(_116_),
    .y(_118_)
  );
  al_nor2 _161_ (
    .a(G12),
    .b(G10),
    .y(_119_)
  );
  al_and3fft _162_ (
    .a(_119_),
    .b(_118_),
    .c(_095_),
    .y(G45)
  );
  al_and3fft _163_ (
    .a(\DFF_3.Q ),
    .b(\DFF_4.Q ),
    .c(_113_),
    .y(G288)
  );
  al_and2ft _164_ (
    .a(G5),
    .b(G288),
    .y(G47)
  );
  al_nand2 _165_ (
    .a(\DFF_2.Q ),
    .b(\DFF_1.Q ),
    .y(_120_)
  );
  al_and3fft _166_ (
    .a(\DFF_3.Q ),
    .b(\DFF_4.Q ),
    .c(G5),
    .y(_121_)
  );
  al_and3fft _167_ (
    .a(\DFF_0.Q ),
    .b(_120_),
    .c(_121_),
    .y(G55)
  );
  al_inv _168_ (
    .a(\DFF_4.Q ),
    .y(_122_)
  );
  al_or2 _169_ (
    .a(\DFF_3.Q ),
    .b(\DFF_2.Q ),
    .y(_123_)
  );
  al_nand2 _170_ (
    .a(G15),
    .b(\DFF_1.Q ),
    .y(_124_)
  );
  al_and3fft _171_ (
    .a(_123_),
    .b(_124_),
    .c(_122_),
    .y(G290)
  );
  al_nor2 _172_ (
    .a(G4),
    .b(\DFF_2.Q ),
    .y(_125_)
  );
  al_and2 _173_ (
    .a(G8),
    .b(G9),
    .y(_126_)
  );
  al_nand3 _174_ (
    .a(G7),
    .b(G6),
    .c(_126_),
    .y(_127_)
  );
  al_or3fft _175_ (
    .a(G15),
    .b(\DFF_0.Q ),
    .c(_127_),
    .y(_128_)
  );
  al_ao21 _176_ (
    .a(G16),
    .b(_128_),
    .c(_112_),
    .y(_129_)
  );
  al_nor3fft _177_ (
    .a(\DFF_1.Q ),
    .b(_125_),
    .c(_129_),
    .y(G292)
  );
  al_and3ftt _178_ (
    .a(\DFF_4.Q ),
    .b(\DFF_3.Q ),
    .c(_113_),
    .y(G296)
  );
  al_and3 _179_ (
    .a(G15),
    .b(\DFF_3.Q ),
    .c(G14),
    .y(_130_)
  );
  al_and3fft _180_ (
    .a(\DFF_0.Q ),
    .b(_108_),
    .c(_130_),
    .y(G298)
  );
  al_nor2 _181_ (
    .a(G16),
    .b(G1),
    .y(_131_)
  );
  al_nor3fft _182_ (
    .a(G3),
    .b(_131_),
    .c(_114_),
    .y(G300)
  );
  al_and3ftt _183_ (
    .a(\DFF_3.Q ),
    .b(\DFF_4.Q ),
    .c(_113_),
    .y(G310)
  );
  al_nor3ftt _184_ (
    .a(G16),
    .b(_097_),
    .c(_120_),
    .y(G312)
  );
  al_nand3 _185_ (
    .a(\DFF_2.Q ),
    .b(\DFF_1.Q ),
    .c(\DFF_4.Q ),
    .y(_132_)
  );
  al_nand3fft _186_ (
    .a(\DFF_0.Q ),
    .b(\DFF_3.Q ),
    .c(G1),
    .y(_000_)
  );
  al_aoi21 _187_ (
    .a(_108_),
    .b(_132_),
    .c(_000_),
    .y(G322)
  );
  al_nor3ftt _188_ (
    .a(\DFF_4.Q ),
    .b(_123_),
    .c(_124_),
    .y(G327)
  );
  al_nand2ft _189_ (
    .a(\DFF_1.Q ),
    .b(\DFF_0.Q ),
    .y(_001_)
  );
  al_nor2 _190_ (
    .a(\DFF_2.Q ),
    .b(\DFF_1.Q ),
    .y(_002_)
  );
  al_oai21ftf _191_ (
    .a(_120_),
    .b(_002_),
    .c(_103_),
    .y(_003_)
  );
  al_ao21 _192_ (
    .a(_001_),
    .b(_003_),
    .c(_099_),
    .y(G49)
  );
  al_ao21 _193_ (
    .a(\DFF_3.Q ),
    .b(\DFF_2.Q ),
    .c(\DFF_1.Q ),
    .y(_004_)
  );
  al_and3 _194_ (
    .a(\DFF_0.Q ),
    .b(G16),
    .c(_115_),
    .y(_005_)
  );
  al_nand3 _195_ (
    .a(_132_),
    .b(_004_),
    .c(_005_),
    .y(_006_)
  );
  al_ao21 _196_ (
    .a(_006_),
    .b(_118_),
    .c(G4),
    .y(_007_)
  );
  al_and2ft _197_ (
    .a(G0),
    .b(\DFF_0.Q ),
    .y(_008_)
  );
  al_aoi21ftt _198_ (
    .a(\DFF_3.Q ),
    .b(\DFF_0.Q ),
    .c(_132_),
    .y(_009_)
  );
  al_ao21ftf _199_ (
    .a(_008_),
    .b(_000_),
    .c(_009_),
    .y(_010_)
  );
  al_nand2ft _200_ (
    .a(\DFF_4.Q ),
    .b(\DFF_0.Q ),
    .y(_011_)
  );
  al_aoi21ttf _201_ (
    .a(\DFF_0.Q ),
    .b(G16),
    .c(\DFF_4.Q ),
    .y(_012_)
  );
  al_oai21ttf _202_ (
    .a(_011_),
    .b(_008_),
    .c(_012_),
    .y(_013_)
  );
  al_or3 _203_ (
    .a(\DFF_0.Q ),
    .b(G16),
    .c(G1),
    .y(_014_)
  );
  al_and3ftt _204_ (
    .a(\DFF_3.Q ),
    .b(_014_),
    .c(_002_),
    .y(_015_)
  );
  al_aoi21ftf _205_ (
    .a(_013_),
    .b(_015_),
    .c(_010_),
    .y(_016_)
  );
  al_aoi21 _206_ (
    .a(_016_),
    .b(_007_),
    .c(G18),
    .y(\DFF_0.D )
  );
  al_nand2ft _207_ (
    .a(G4),
    .b(_103_),
    .y(_017_)
  );
  al_ao21ftf _208_ (
    .a(_112_),
    .b(_008_),
    .c(_017_),
    .y(_018_)
  );
  al_or3 _209_ (
    .a(\DFF_3.Q ),
    .b(G1),
    .c(G3),
    .y(_019_)
  );
  al_nand2 _210_ (
    .a(\DFF_4.Q ),
    .b(_019_),
    .y(_020_)
  );
  al_nand3ftt _211_ (
    .a(_121_),
    .b(_113_),
    .c(_020_),
    .y(_021_)
  );
  al_aoi21ftf _212_ (
    .a(_120_),
    .b(_018_),
    .c(_021_),
    .y(_022_)
  );
  al_and3fft _213_ (
    .a(G4),
    .b(\DFF_1.Q ),
    .c(G16),
    .y(_023_)
  );
  al_ao21ftf _214_ (
    .a(\DFF_4.Q ),
    .b(\DFF_0.Q ),
    .c(_023_),
    .y(_024_)
  );
  al_and3ftt _215_ (
    .a(\DFF_4.Q ),
    .b(G11),
    .c(_119_),
    .y(_025_)
  );
  al_and2 _216_ (
    .a(G15),
    .b(\DFF_2.Q ),
    .y(_026_)
  );
  al_and2ft _217_ (
    .a(\DFF_4.Q ),
    .b(G10),
    .y(_027_)
  );
  al_nand3fft _218_ (
    .a(G12),
    .b(G11),
    .c(_027_),
    .y(_028_)
  );
  al_and3 _219_ (
    .a(\DFF_3.Q ),
    .b(_026_),
    .c(_028_),
    .y(_029_)
  );
  al_nand3fft _220_ (
    .a(_024_),
    .b(_025_),
    .c(_029_),
    .y(_030_)
  );
  al_and3ftt _221_ (
    .a(G3),
    .b(G2),
    .c(_131_),
    .y(_031_)
  );
  al_nand3ftt _222_ (
    .a(_108_),
    .b(_109_),
    .c(_031_),
    .y(_032_)
  );
  al_or3fft _223_ (
    .a(\DFF_1.Q ),
    .b(_125_),
    .c(_106_),
    .y(_033_)
  );
  al_and3 _224_ (
    .a(_032_),
    .b(_033_),
    .c(_030_),
    .y(_034_)
  );
  al_aoi21 _225_ (
    .a(_022_),
    .b(_034_),
    .c(G18),
    .y(\DFF_1.D )
  );
  al_nor2 _226_ (
    .a(\DFF_2.Q ),
    .b(\DFF_4.Q ),
    .y(_035_)
  );
  al_oa21ftt _227_ (
    .a(G15),
    .b(G14),
    .c(\DFF_3.Q ),
    .y(_036_)
  );
  al_and3fft _228_ (
    .a(_100_),
    .b(_036_),
    .c(_035_),
    .y(_037_)
  );
  al_oai21 _229_ (
    .a(\DFF_3.Q ),
    .b(_031_),
    .c(_037_),
    .y(_038_)
  );
  al_aoi21ftt _230_ (
    .a(\DFF_3.Q ),
    .b(\DFF_0.Q ),
    .c(_024_),
    .y(_039_)
  );
  al_oai21ftf _231_ (
    .a(G15),
    .b(_097_),
    .c(\DFF_2.Q ),
    .y(_040_)
  );
  al_oai21ttf _232_ (
    .a(G10),
    .b(G11),
    .c(\DFF_4.Q ),
    .y(_041_)
  );
  al_nand3 _233_ (
    .a(\DFF_3.Q ),
    .b(_041_),
    .c(_026_),
    .y(_042_)
  );
  al_nand3 _234_ (
    .a(_040_),
    .b(_042_),
    .c(_039_),
    .y(_043_)
  );
  al_and3 _235_ (
    .a(_038_),
    .b(_043_),
    .c(_022_),
    .y(_044_)
  );
  al_oa21ftf _236_ (
    .a(_044_),
    .b(G292),
    .c(G18),
    .y(\DFF_2.D )
  );
  al_nand2ft _237_ (
    .a(\DFF_3.Q ),
    .b(\DFF_4.Q ),
    .y(_045_)
  );
  al_aoi21ftt _238_ (
    .a(_045_),
    .b(_026_),
    .c(_096_),
    .y(_046_)
  );
  al_ao21 _239_ (
    .a(\DFF_3.Q ),
    .b(\DFF_4.Q ),
    .c(\DFF_2.Q ),
    .y(_047_)
  );
  al_aoi21 _240_ (
    .a(G4),
    .b(_047_),
    .c(\DFF_1.Q ),
    .y(_048_)
  );
  al_aoi21ftf _241_ (
    .a(_036_),
    .b(_035_),
    .c(_048_),
    .y(_049_)
  );
  al_ao21ftf _242_ (
    .a(_035_),
    .b(_046_),
    .c(_049_),
    .y(_050_)
  );
  al_or3ftt _243_ (
    .a(\DFF_3.Q ),
    .b(G4),
    .c(\DFF_4.Q ),
    .y(_051_)
  );
  al_nand2ft _244_ (
    .a(\DFF_1.Q ),
    .b(_051_),
    .y(_052_)
  );
  al_oai21ftf _245_ (
    .a(G5),
    .b(\DFF_4.Q ),
    .c(\DFF_3.Q ),
    .y(_053_)
  );
  al_aoi21ttf _246_ (
    .a(G16),
    .b(\DFF_4.Q ),
    .c(\DFF_2.Q ),
    .y(_054_)
  );
  al_nand3 _247_ (
    .a(_053_),
    .b(_054_),
    .c(_052_),
    .y(_055_)
  );
  al_aoi21ftf _248_ (
    .a(G16),
    .b(_002_),
    .c(_132_),
    .y(_056_)
  );
  al_nor2ft _249_ (
    .a(G2),
    .b(_019_),
    .y(_057_)
  );
  al_aoi21ftf _250_ (
    .a(_056_),
    .b(_057_),
    .c(_055_),
    .y(_058_)
  );
  al_ao21 _251_ (
    .a(_058_),
    .b(_050_),
    .c(\DFF_0.Q ),
    .y(_059_)
  );
  al_nand3ftt _252_ (
    .a(G0),
    .b(\DFF_0.Q ),
    .c(\DFF_1.Q ),
    .y(_060_)
  );
  al_nand3 _253_ (
    .a(G13),
    .b(G15),
    .c(G16),
    .y(_061_)
  );
  al_nand3fft _254_ (
    .a(G4),
    .b(\DFF_1.Q ),
    .c(_061_),
    .y(_062_)
  );
  al_aoi21 _255_ (
    .a(_060_),
    .b(_062_),
    .c(_098_),
    .y(_063_)
  );
  al_aoi21ttf _256_ (
    .a(G15),
    .b(\DFF_4.Q ),
    .c(G16),
    .y(_064_)
  );
  al_oai21ftf _257_ (
    .a(G16),
    .b(G15),
    .c(\DFF_1.Q ),
    .y(_065_)
  );
  al_and3 _258_ (
    .a(_001_),
    .b(_125_),
    .c(_065_),
    .y(_066_)
  );
  al_aoi21ftf _259_ (
    .a(\DFF_3.Q ),
    .b(_064_),
    .c(_066_),
    .y(_067_)
  );
  al_aoi21 _260_ (
    .a(_067_),
    .b(_129_),
    .c(_063_),
    .y(_068_)
  );
  al_aoi21 _261_ (
    .a(_059_),
    .b(_068_),
    .c(G18),
    .y(\DFF_3.D )
  );
  al_or3 _262_ (
    .a(\DFF_3.Q ),
    .b(\DFF_2.Q ),
    .c(G1),
    .y(_069_)
  );
  al_and2ft _263_ (
    .a(G7),
    .b(G6),
    .y(_070_)
  );
  al_and3ftt _264_ (
    .a(G8),
    .b(G15),
    .c(\DFF_2.Q ),
    .y(_071_)
  );
  al_nand3 _265_ (
    .a(G9),
    .b(_071_),
    .c(_070_),
    .y(_072_)
  );
  al_mux2h _266_ (
    .a(G15),
    .b(_072_),
    .s(_122_),
    .y(_073_)
  );
  al_ao21 _267_ (
    .a(_069_),
    .b(_073_),
    .c(_100_),
    .y(_074_)
  );
  al_inv _268_ (
    .a(\DFF_2.Q ),
    .y(_075_)
  );
  al_nand2 _269_ (
    .a(\DFF_0.Q ),
    .b(\DFF_1.Q ),
    .y(_076_)
  );
  al_ao21 _270_ (
    .a(_075_),
    .b(_127_),
    .c(_076_),
    .y(_077_)
  );
  al_nand3 _271_ (
    .a(G13),
    .b(G15),
    .c(\DFF_4.Q ),
    .y(_078_)
  );
  al_oai21ftf _272_ (
    .a(G15),
    .b(\DFF_0.Q ),
    .c(\DFF_4.Q ),
    .y(_079_)
  );
  al_ao21 _273_ (
    .a(_079_),
    .b(_078_),
    .c(\DFF_1.Q ),
    .y(_080_)
  );
  al_ao21 _274_ (
    .a(G15),
    .b(\DFF_1.Q ),
    .c(\DFF_2.Q ),
    .y(_081_)
  );
  al_and3 _275_ (
    .a(\DFF_3.Q ),
    .b(_081_),
    .c(_080_),
    .y(_082_)
  );
  al_oai21 _276_ (
    .a(\DFF_2.Q ),
    .b(\DFF_4.Q ),
    .c(_081_),
    .y(_083_)
  );
  al_oa21 _277_ (
    .a(G15),
    .b(\DFF_4.Q ),
    .c(\DFF_1.Q ),
    .y(_084_)
  );
  al_aoi21ftf _278_ (
    .a(_084_),
    .b(_045_),
    .c(_083_),
    .y(_085_)
  );
  al_aoi21 _279_ (
    .a(_077_),
    .b(_082_),
    .c(_085_),
    .y(_086_)
  );
  al_ao21 _280_ (
    .a(_074_),
    .b(_086_),
    .c(_096_),
    .y(_087_)
  );
  al_nand2ft _281_ (
    .a(\DFF_1.Q ),
    .b(G4),
    .y(_088_)
  );
  al_aoi21 _282_ (
    .a(G2),
    .b(\DFF_4.Q ),
    .c(_120_),
    .y(_089_)
  );
  al_nand3ftt _283_ (
    .a(_121_),
    .b(_020_),
    .c(_089_),
    .y(_090_)
  );
  al_ao21ftf _284_ (
    .a(_088_),
    .b(_047_),
    .c(_090_),
    .y(_091_)
  );
  al_ao21 _285_ (
    .a(_060_),
    .b(_088_),
    .c(_098_),
    .y(_092_)
  );
  al_and3ftt _286_ (
    .a(G298),
    .b(_105_),
    .c(_092_),
    .y(_093_)
  );
  al_aoi21ftf _287_ (
    .a(\DFF_0.Q ),
    .b(_091_),
    .c(_093_),
    .y(_094_)
  );
  al_aoi21 _288_ (
    .a(_094_),
    .b(_087_),
    .c(G18),
    .y(\DFF_4.D )
  );
  al_dffl _289_ (
    .clk(CK),
    .d(\DFF_0.D ),
    .q(\DFF_0.Q )
  );
  al_dffl _290_ (
    .clk(CK),
    .d(\DFF_1.D ),
    .q(\DFF_1.Q )
  );
  al_dffl _291_ (
    .clk(CK),
    .d(\DFF_2.D ),
    .q(\DFF_2.Q )
  );
  al_dffl _292_ (
    .clk(CK),
    .d(\DFF_3.D ),
    .q(\DFF_3.Q )
  );
  al_dffl _293_ (
    .clk(CK),
    .d(\DFF_4.D ),
    .q(\DFF_4.Q )
  );
  assign \DFF_0.CK  = CK;
  assign \DFF_1.CK  = CK;
  assign \DFF_2.CK  = CK;
  assign \DFF_3.CK  = CK;
  assign \DFF_4.CK  = CK;
  assign G102 = \DFF_4.D ;
  assign G325 = G310;
  assign G38 = \DFF_0.Q ;
  assign G39 = \DFF_1.Q ;
  assign G40 = \DFF_2.Q ;
  assign G41 = \DFF_3.Q ;
  assign G42 = \DFF_4.Q ;
  assign G90 = \DFF_0.D ;
  assign G93 = \DFF_1.D ;
  assign G96 = \DFF_2.D ;
  assign G99 = \DFF_3.D ;
endmodule
