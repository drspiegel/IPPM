
module c6288(N1, N18, N35, N52, N69, N86, N103, N120, N137, N154, N171, N188, N205, N222, N239, N256, N273, N290, N307, N324, N341, N358, N375, N392, N409, N426, N443, N460, N477, N494, N511, N528, N545, N1581, N1901, N2223, N2548, N2877, N3211, N3552, N3895, N4241, N4591, N4946, N5308, N5672, N5971, N6123, N6150, N6160, N6170, N6180, N6190, N6200, N6210, N6220, N6230, N6240, N6250, N6260, N6270, N6280, N6287, N6288);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  input N1;
  input N103;
  input N120;
  input N137;
  input N154;
  output N1581;
  input N171;
  input N18;
  input N188;
  output N1901;
  input N205;
  input N222;
  output N2223;
  input N239;
  output N2548;
  input N256;
  input N273;
  output N2877;
  input N290;
  input N307;
  output N3211;
  input N324;
  input N341;
  input N35;
  output N3552;
  input N358;
  input N375;
  output N3895;
  input N392;
  input N409;
  output N4241;
  input N426;
  input N443;
  output N4591;
  input N460;
  input N477;
  input N494;
  output N4946;
  input N511;
  input N52;
  input N528;
  output N5308;
  output N545;
  output N5672;
  output N5971;
  output N6123;
  wire N6141;
  output N6150;
  output N6160;
  output N6170;
  output N6180;
  output N6190;
  output N6200;
  output N6210;
  output N6220;
  output N6230;
  output N6240;
  output N6250;
  output N6260;
  output N6270;
  output N6280;
  output N6287;
  output N6288;
  input N69;
  input N86;
  al_and2ft _1444_ (
    .a(_0045_),
    .b(_0046_),
    .y(_0048_)
  );
  al_nor2 _1445_ (
    .a(_0048_),
    .b(_1407_),
    .y(_0049_)
  );
  al_or2ft _1446_ (
    .a(_0047_),
    .b(_0049_),
    .y(N6170)
  );
  al_ao21 _1447_ (
    .a(_0048_),
    .b(_1407_),
    .c(_0045_),
    .y(_0050_)
  );
  al_ao21ttf _1448_ (
    .a(_1409_),
    .b(_0041_),
    .c(_0040_),
    .y(_0051_)
  );
  al_nand2 _1449_ (
    .a(N528),
    .b(N69),
    .y(_0052_)
  );
  al_ao21ttf _1450_ (
    .a(_1412_),
    .b(_0037_),
    .c(_0036_),
    .y(_0053_)
  );
  al_nand2 _1451_ (
    .a(N511),
    .b(N86),
    .y(_0055_)
  );
  al_ao21ttf _1452_ (
    .a(_1414_),
    .b(_0032_),
    .c(_0031_),
    .y(_0056_)
  );
  al_nand2 _1453_ (
    .a(N494),
    .b(N103),
    .y(_0057_)
  );
  al_ao21ttf _1454_ (
    .a(_1416_),
    .b(_0028_),
    .c(_0027_),
    .y(_0058_)
  );
  al_nand2 _1455_ (
    .a(N477),
    .b(N120),
    .y(_0059_)
  );
  al_ao21ttf _1456_ (
    .a(_1418_),
    .b(_0024_),
    .c(_0023_),
    .y(_0060_)
  );
  al_nand2 _1457_ (
    .a(N460),
    .b(N137),
    .y(_0061_)
  );
  al_ao21ttf _1458_ (
    .a(_1420_),
    .b(_0019_),
    .c(_0018_),
    .y(_0062_)
  );
  al_nand2 _1459_ (
    .a(N443),
    .b(N154),
    .y(_0063_)
  );
  al_ao21ttf _1460_ (
    .a(_1423_),
    .b(_0015_),
    .c(_0014_),
    .y(_0064_)
  );
  al_nand2 _1461_ (
    .a(N426),
    .b(N171),
    .y(_0066_)
  );
  al_ao21ttf _1462_ (
    .a(_1425_),
    .b(_0010_),
    .c(_0009_),
    .y(_0067_)
  );
  al_nand2 _1463_ (
    .a(N409),
    .b(N188),
    .y(_0068_)
  );
  al_ao21ttf _1464_ (
    .a(_1427_),
    .b(_0006_),
    .c(_0005_),
    .y(_0069_)
  );
  al_nand2 _1465_ (
    .a(N392),
    .b(N205),
    .y(_0070_)
  );
  al_ao21ttf _1466_ (
    .a(_1429_),
    .b(_0002_),
    .c(_0001_),
    .y(_0071_)
  );
  al_nand2 _1467_ (
    .a(N375),
    .b(N222),
    .y(_0072_)
  );
  al_ao21ttf _1468_ (
    .a(_1431_),
    .b(_1441_),
    .c(_1440_),
    .y(_0073_)
  );
  al_inv _1469_ (
    .a(N239),
    .y(_0074_)
  );
  al_ao21ttf _1470_ (
    .a(_1434_),
    .b(_1437_),
    .c(_1436_),
    .y(_0075_)
  );
  al_ao21ftf _1471_ (
    .a(_1344_),
    .b(N341),
    .c(_0075_),
    .y(_0077_)
  );
  al_and3fft _1472_ (
    .a(_1344_),
    .b(_0075_),
    .c(N341),
    .y(_0078_)
  );
  al_or2ft _1473_ (
    .a(_0077_),
    .b(_0078_),
    .y(_0079_)
  );
  al_ao21ftt _1474_ (
    .a(_0074_),
    .b(N358),
    .c(_0079_),
    .y(_0080_)
  );
  al_nand3 _1475_ (
    .a(N358),
    .b(N239),
    .c(_0079_),
    .y(_0081_)
  );
  al_nand3 _1476_ (
    .a(_0073_),
    .b(_0081_),
    .c(_0080_),
    .y(_0082_)
  );
  al_ao21 _1477_ (
    .a(_0081_),
    .b(_0080_),
    .c(_0073_),
    .y(_0083_)
  );
  al_nand3 _1478_ (
    .a(_0072_),
    .b(_0083_),
    .c(_0082_),
    .y(_0084_)
  );
  al_ao21 _1479_ (
    .a(_0083_),
    .b(_0082_),
    .c(_0072_),
    .y(_0085_)
  );
  al_nand3 _1480_ (
    .a(_0084_),
    .b(_0085_),
    .c(_0071_),
    .y(_0086_)
  );
  al_ao21 _1481_ (
    .a(_0084_),
    .b(_0085_),
    .c(_0071_),
    .y(_0088_)
  );
  al_nand3 _1482_ (
    .a(_0070_),
    .b(_0086_),
    .c(_0088_),
    .y(_0089_)
  );
  al_ao21 _1483_ (
    .a(_0086_),
    .b(_0088_),
    .c(_0070_),
    .y(_0090_)
  );
  al_nand3 _1484_ (
    .a(_0089_),
    .b(_0090_),
    .c(_0069_),
    .y(_0091_)
  );
  al_ao21 _1485_ (
    .a(_0089_),
    .b(_0090_),
    .c(_0069_),
    .y(_0092_)
  );
  al_and3 _1486_ (
    .a(_0068_),
    .b(_0091_),
    .c(_0092_),
    .y(_0093_)
  );
  al_ao21 _1487_ (
    .a(_0091_),
    .b(_0092_),
    .c(_0068_),
    .y(_0094_)
  );
  al_and3ftt _1488_ (
    .a(_0093_),
    .b(_0094_),
    .c(_0067_),
    .y(_0095_)
  );
  al_ao21ftt _1489_ (
    .a(_0093_),
    .b(_0094_),
    .c(_0067_),
    .y(_0096_)
  );
  al_nor3fft _1490_ (
    .a(_0066_),
    .b(_0096_),
    .c(_0095_),
    .y(_0097_)
  );
  al_oai21ftf _1491_ (
    .a(_0096_),
    .b(_0095_),
    .c(_0066_),
    .y(_0099_)
  );
  al_and3ftt _1492_ (
    .a(_0097_),
    .b(_0099_),
    .c(_0064_),
    .y(_0100_)
  );
  al_ao21ftt _1493_ (
    .a(_0097_),
    .b(_0099_),
    .c(_0064_),
    .y(_0101_)
  );
  al_nor3fft _1494_ (
    .a(_0063_),
    .b(_0101_),
    .c(_0100_),
    .y(_0102_)
  );
  al_oai21ftf _1495_ (
    .a(_0101_),
    .b(_0100_),
    .c(_0063_),
    .y(_0103_)
  );
  al_and3ftt _1496_ (
    .a(_0102_),
    .b(_0103_),
    .c(_0062_),
    .y(_0104_)
  );
  al_ao21ftt _1497_ (
    .a(_0102_),
    .b(_0103_),
    .c(_0062_),
    .y(_0105_)
  );
  al_nor3fft _1498_ (
    .a(_0061_),
    .b(_0105_),
    .c(_0104_),
    .y(_0106_)
  );
  al_oai21ftf _1499_ (
    .a(_0105_),
    .b(_0104_),
    .c(_0061_),
    .y(_0107_)
  );
  al_and3ftt _1500_ (
    .a(_0106_),
    .b(_0107_),
    .c(_0060_),
    .y(_0108_)
  );
  al_ao21ftt _1501_ (
    .a(_0106_),
    .b(_0107_),
    .c(_0060_),
    .y(_0110_)
  );
  al_nor3fft _1502_ (
    .a(_0059_),
    .b(_0110_),
    .c(_0108_),
    .y(_0111_)
  );
  al_oai21ftf _1503_ (
    .a(_0110_),
    .b(_0108_),
    .c(_0059_),
    .y(_0112_)
  );
  al_nand3ftt _1504_ (
    .a(_0111_),
    .b(_0112_),
    .c(_0058_),
    .y(_0113_)
  );
  al_ao21ftt _1505_ (
    .a(_0111_),
    .b(_0112_),
    .c(_0058_),
    .y(_0114_)
  );
  al_and3 _1506_ (
    .a(_0057_),
    .b(_0113_),
    .c(_0114_),
    .y(_0115_)
  );
  al_ao21 _1507_ (
    .a(_0113_),
    .b(_0114_),
    .c(_0057_),
    .y(_0116_)
  );
  al_nand3ftt _1508_ (
    .a(_0115_),
    .b(_0116_),
    .c(_0056_),
    .y(_0117_)
  );
  al_ao21ftt _1509_ (
    .a(_0115_),
    .b(_0116_),
    .c(_0056_),
    .y(_0118_)
  );
  al_and3 _1510_ (
    .a(_0055_),
    .b(_0117_),
    .c(_0118_),
    .y(_0119_)
  );
  al_ao21 _1511_ (
    .a(_0117_),
    .b(_0118_),
    .c(_0055_),
    .y(_0121_)
  );
  al_nand3ftt _1512_ (
    .a(_0119_),
    .b(_0121_),
    .c(_0053_),
    .y(_0122_)
  );
  al_ao21ftt _1513_ (
    .a(_0119_),
    .b(_0121_),
    .c(_0053_),
    .y(_0123_)
  );
  al_and3 _1514_ (
    .a(_0052_),
    .b(_0122_),
    .c(_0123_),
    .y(_0124_)
  );
  al_ao21 _1515_ (
    .a(_0122_),
    .b(_0123_),
    .c(_0052_),
    .y(_0125_)
  );
  al_and3ftt _1516_ (
    .a(_0124_),
    .b(_0125_),
    .c(_0051_),
    .y(_0126_)
  );
  al_ao21ftt _1517_ (
    .a(_0124_),
    .b(_0125_),
    .c(_0051_),
    .y(_0127_)
  );
  al_and2ft _1518_ (
    .a(_0126_),
    .b(_0127_),
    .y(_0128_)
  );
  al_nand2 _1519_ (
    .a(_0128_),
    .b(_0050_),
    .y(_0129_)
  );
  al_and3fft _1520_ (
    .a(_0045_),
    .b(_0128_),
    .c(_0047_),
    .y(_0130_)
  );
  al_nand2ft _1521_ (
    .a(_0130_),
    .b(_0129_),
    .y(N6180)
  );
  al_ao21 _1522_ (
    .a(_0128_),
    .b(_0050_),
    .c(_0126_),
    .y(_0132_)
  );
  al_ao21ttf _1523_ (
    .a(_0052_),
    .b(_0123_),
    .c(_0122_),
    .y(_0133_)
  );
  al_nand2 _1524_ (
    .a(N528),
    .b(N86),
    .y(_0134_)
  );
  al_ao21ttf _1525_ (
    .a(_0055_),
    .b(_0118_),
    .c(_0117_),
    .y(_0135_)
  );
  al_nand2 _1526_ (
    .a(N511),
    .b(N103),
    .y(_0136_)
  );
  al_ao21ttf _1527_ (
    .a(_0057_),
    .b(_0114_),
    .c(_0113_),
    .y(_0137_)
  );
  al_nand2 _1528_ (
    .a(N494),
    .b(N120),
    .y(_0138_)
  );
  al_ao21 _1529_ (
    .a(_0059_),
    .b(_0110_),
    .c(_0108_),
    .y(_0139_)
  );
  al_nand2 _1530_ (
    .a(N477),
    .b(N137),
    .y(_0140_)
  );
  al_ao21 _1531_ (
    .a(_0061_),
    .b(_0105_),
    .c(_0104_),
    .y(_0142_)
  );
  al_nand2 _1532_ (
    .a(N460),
    .b(N154),
    .y(_0143_)
  );
  al_ao21 _1533_ (
    .a(_0063_),
    .b(_0101_),
    .c(_0100_),
    .y(_0144_)
  );
  al_nand2 _1534_ (
    .a(N443),
    .b(N171),
    .y(_0145_)
  );
  al_ao21 _1535_ (
    .a(_0066_),
    .b(_0096_),
    .c(_0095_),
    .y(_0146_)
  );
  al_nand2 _1536_ (
    .a(N426),
    .b(N188),
    .y(_0147_)
  );
  al_ao21ttf _1537_ (
    .a(_0068_),
    .b(_0092_),
    .c(_0091_),
    .y(_0148_)
  );
  al_nand2 _1538_ (
    .a(N409),
    .b(N205),
    .y(_0149_)
  );
  al_ao21ttf _1539_ (
    .a(_0070_),
    .b(_0088_),
    .c(_0086_),
    .y(_0150_)
  );
  al_nand2 _1540_ (
    .a(N392),
    .b(N222),
    .y(_0151_)
  );
  al_ao21ttf _1541_ (
    .a(_0072_),
    .b(_0083_),
    .c(_0082_),
    .y(_0153_)
  );
  al_nand2 _1542_ (
    .a(N375),
    .b(N239),
    .y(_0154_)
  );
  al_nand2 _1543_ (
    .a(_0077_),
    .b(_0080_),
    .y(_0155_)
  );
  al_ao21ftf _1544_ (
    .a(_1344_),
    .b(N358),
    .c(_0155_),
    .y(_0156_)
  );
  al_or3fft _1545_ (
    .a(N358),
    .b(N256),
    .c(_0155_),
    .y(_0157_)
  );
  al_nand3 _1546_ (
    .a(_0154_),
    .b(_0156_),
    .c(_0157_),
    .y(_0158_)
  );
  al_ao21 _1547_ (
    .a(_0156_),
    .b(_0157_),
    .c(_0154_),
    .y(_0159_)
  );
  al_nand3 _1548_ (
    .a(_0153_),
    .b(_0158_),
    .c(_0159_),
    .y(_0160_)
  );
  al_ao21 _1549_ (
    .a(_0158_),
    .b(_0159_),
    .c(_0153_),
    .y(_0161_)
  );
  al_nand3 _1550_ (
    .a(_0151_),
    .b(_0160_),
    .c(_0161_),
    .y(_0162_)
  );
  al_ao21 _1551_ (
    .a(_0160_),
    .b(_0161_),
    .c(_0151_),
    .y(_0164_)
  );
  al_nand3 _1552_ (
    .a(_0150_),
    .b(_0162_),
    .c(_0164_),
    .y(_0165_)
  );
  al_ao21 _1553_ (
    .a(_0162_),
    .b(_0164_),
    .c(_0150_),
    .y(_0166_)
  );
  al_nand3 _1554_ (
    .a(_0149_),
    .b(_0165_),
    .c(_0166_),
    .y(_0167_)
  );
  al_ao21 _1555_ (
    .a(_0165_),
    .b(_0166_),
    .c(_0149_),
    .y(_0168_)
  );
  al_nand3 _1556_ (
    .a(_0167_),
    .b(_0148_),
    .c(_0168_),
    .y(_0169_)
  );
  al_ao21 _1557_ (
    .a(_0167_),
    .b(_0168_),
    .c(_0148_),
    .y(_0170_)
  );
  al_and3 _1558_ (
    .a(_0147_),
    .b(_0169_),
    .c(_0170_),
    .y(_0171_)
  );
  al_ao21 _1559_ (
    .a(_0169_),
    .b(_0170_),
    .c(_0147_),
    .y(_0172_)
  );
  al_and3ftt _1560_ (
    .a(_0171_),
    .b(_0146_),
    .c(_0172_),
    .y(_0173_)
  );
  al_ao21ftt _1561_ (
    .a(_0171_),
    .b(_0172_),
    .c(_0146_),
    .y(_0174_)
  );
  al_nor3fft _1562_ (
    .a(_0145_),
    .b(_0174_),
    .c(_0173_),
    .y(_0175_)
  );
  al_oai21ftf _1563_ (
    .a(_0174_),
    .b(_0173_),
    .c(_0145_),
    .y(_0176_)
  );
  al_and3ftt _1564_ (
    .a(_0175_),
    .b(_0144_),
    .c(_0176_),
    .y(_0177_)
  );
  al_ao21ftt _1565_ (
    .a(_0175_),
    .b(_0176_),
    .c(_0144_),
    .y(_0178_)
  );
  al_nor3fft _1566_ (
    .a(_0143_),
    .b(_0178_),
    .c(_0177_),
    .y(_0179_)
  );
  al_oai21ftf _1567_ (
    .a(_0178_),
    .b(_0177_),
    .c(_0143_),
    .y(_0180_)
  );
  al_and3ftt _1568_ (
    .a(_0179_),
    .b(_0142_),
    .c(_0180_),
    .y(_0181_)
  );
  al_ao21ftt _1569_ (
    .a(_0179_),
    .b(_0180_),
    .c(_0142_),
    .y(_0182_)
  );
  al_nor3fft _1570_ (
    .a(_0140_),
    .b(_0182_),
    .c(_0181_),
    .y(_0183_)
  );
  al_oai21ftf _1571_ (
    .a(_0182_),
    .b(_0181_),
    .c(_0140_),
    .y(_0185_)
  );
  al_and3ftt _1572_ (
    .a(_0183_),
    .b(_0139_),
    .c(_0185_),
    .y(_0186_)
  );
  al_ao21ftt _1573_ (
    .a(_0183_),
    .b(_0185_),
    .c(_0139_),
    .y(_0187_)
  );
  al_nor3fft _1574_ (
    .a(_0138_),
    .b(_0187_),
    .c(_0186_),
    .y(_0188_)
  );
  al_oai21ftf _1575_ (
    .a(_0187_),
    .b(_0186_),
    .c(_0138_),
    .y(_0189_)
  );
  al_and3ftt _1576_ (
    .a(_0188_),
    .b(_0137_),
    .c(_0189_),
    .y(_0190_)
  );
  al_ao21ftt _1577_ (
    .a(_0188_),
    .b(_0189_),
    .c(_0137_),
    .y(_0191_)
  );
  al_nor3fft _1578_ (
    .a(_0136_),
    .b(_0191_),
    .c(_0190_),
    .y(_0192_)
  );
  al_oai21ftf _1579_ (
    .a(_0191_),
    .b(_0190_),
    .c(_0136_),
    .y(_0193_)
  );
  al_nor3fft _1580_ (
    .a(_0135_),
    .b(_0193_),
    .c(_0192_),
    .y(_0194_)
  );
  al_ao21ftt _1581_ (
    .a(_0192_),
    .b(_0193_),
    .c(_0135_),
    .y(_0196_)
  );
  al_nor3fft _1582_ (
    .a(_0134_),
    .b(_0196_),
    .c(_0194_),
    .y(_0197_)
  );
  al_oai21ftf _1583_ (
    .a(_0196_),
    .b(_0194_),
    .c(_0134_),
    .y(_0198_)
  );
  al_nor3fft _1584_ (
    .a(_0133_),
    .b(_0198_),
    .c(_0197_),
    .y(_0199_)
  );
  al_ao21ftt _1585_ (
    .a(_0197_),
    .b(_0198_),
    .c(_0133_),
    .y(_0200_)
  );
  al_and2ft _1586_ (
    .a(_0199_),
    .b(_0200_),
    .y(_0201_)
  );
  al_nand2 _1587_ (
    .a(_0201_),
    .b(_0132_),
    .y(_0202_)
  );
  al_and3fft _1588_ (
    .a(_0126_),
    .b(_0201_),
    .c(_0129_),
    .y(_0203_)
  );
  al_nand2ft _1589_ (
    .a(_0203_),
    .b(_0202_),
    .y(N6190)
  );
  al_ao21 _1590_ (
    .a(_0201_),
    .b(_0132_),
    .c(_0199_),
    .y(_0204_)
  );
  al_ao21 _1591_ (
    .a(_0134_),
    .b(_0196_),
    .c(_0194_),
    .y(_0206_)
  );
  al_nand2 _1592_ (
    .a(N528),
    .b(N103),
    .y(_0207_)
  );
  al_ao21 _1593_ (
    .a(_0136_),
    .b(_0191_),
    .c(_0190_),
    .y(_0208_)
  );
  al_nand2 _1594_ (
    .a(N511),
    .b(N120),
    .y(_0209_)
  );
  al_ao21 _1595_ (
    .a(_0138_),
    .b(_0187_),
    .c(_0186_),
    .y(_0210_)
  );
  al_nand2 _1596_ (
    .a(N494),
    .b(N137),
    .y(_0211_)
  );
  al_ao21 _1597_ (
    .a(_0140_),
    .b(_0182_),
    .c(_0181_),
    .y(_0212_)
  );
  al_nand2 _1598_ (
    .a(N477),
    .b(N154),
    .y(_0213_)
  );
  al_ao21 _1599_ (
    .a(_0143_),
    .b(_0178_),
    .c(_0177_),
    .y(_0214_)
  );
  al_nand2 _1600_ (
    .a(N460),
    .b(N171),
    .y(_0215_)
  );
  al_ao21 _1601_ (
    .a(_0145_),
    .b(_0174_),
    .c(_0173_),
    .y(_0217_)
  );
  al_nand2 _1602_ (
    .a(N443),
    .b(N188),
    .y(_0218_)
  );
  al_ao21ttf _1603_ (
    .a(_0147_),
    .b(_0170_),
    .c(_0169_),
    .y(_0219_)
  );
  al_nand2 _1604_ (
    .a(N426),
    .b(N205),
    .y(_0220_)
  );
  al_ao21ttf _1605_ (
    .a(_0149_),
    .b(_0166_),
    .c(_0165_),
    .y(_0221_)
  );
  al_nand2 _1606_ (
    .a(N409),
    .b(N222),
    .y(_0222_)
  );
  al_ao21ttf _1607_ (
    .a(_0151_),
    .b(_0161_),
    .c(_0160_),
    .y(_0223_)
  );
  al_nand2 _1608_ (
    .a(N392),
    .b(N239),
    .y(_0224_)
  );
  al_ao21ttf _1609_ (
    .a(_0154_),
    .b(_0157_),
    .c(_0156_),
    .y(_0225_)
  );
  al_ao21ftf _1610_ (
    .a(_1344_),
    .b(N375),
    .c(_0225_),
    .y(_0226_)
  );
  al_or3fft _1611_ (
    .a(N375),
    .b(N256),
    .c(_0225_),
    .y(_0227_)
  );
  al_nand3 _1612_ (
    .a(_0224_),
    .b(_0226_),
    .c(_0227_),
    .y(_0228_)
  );
  al_aoi21 _1613_ (
    .a(_0226_),
    .b(_0227_),
    .c(_0224_),
    .y(_0229_)
  );
  al_or3fft _1614_ (
    .a(_0228_),
    .b(_0223_),
    .c(_0229_),
    .y(_0230_)
  );
  al_oai21ftf _1615_ (
    .a(_0228_),
    .b(_0229_),
    .c(_0223_),
    .y(_0231_)
  );
  al_nand3 _1616_ (
    .a(_0222_),
    .b(_0230_),
    .c(_0231_),
    .y(_0232_)
  );
  al_ao21 _1617_ (
    .a(_0230_),
    .b(_0231_),
    .c(_0222_),
    .y(_0233_)
  );
  al_nand3 _1618_ (
    .a(_0232_),
    .b(_0233_),
    .c(_0221_),
    .y(_0234_)
  );
  al_ao21 _1619_ (
    .a(_0232_),
    .b(_0233_),
    .c(_0221_),
    .y(_0235_)
  );
  al_nand3 _1620_ (
    .a(_0220_),
    .b(_0235_),
    .c(_0234_),
    .y(_0236_)
  );
  al_ao21 _1621_ (
    .a(_0235_),
    .b(_0234_),
    .c(_0220_),
    .y(_0239_)
  );
  al_nand3 _1622_ (
    .a(_0219_),
    .b(_0236_),
    .c(_0239_),
    .y(_0240_)
  );
  al_ao21 _1623_ (
    .a(_0236_),
    .b(_0239_),
    .c(_0219_),
    .y(_0241_)
  );
  al_nand3 _1624_ (
    .a(_0218_),
    .b(_0240_),
    .c(_0241_),
    .y(_0242_)
  );
  al_ao21 _1625_ (
    .a(_0240_),
    .b(_0241_),
    .c(_0218_),
    .y(_0243_)
  );
  al_and3 _1626_ (
    .a(_0242_),
    .b(_0217_),
    .c(_0243_),
    .y(_0244_)
  );
  al_ao21 _1627_ (
    .a(_0242_),
    .b(_0243_),
    .c(_0217_),
    .y(_0245_)
  );
  al_or3fft _1628_ (
    .a(_0215_),
    .b(_0245_),
    .c(_0244_),
    .y(_0246_)
  );
  al_oai21ftf _1629_ (
    .a(_0245_),
    .b(_0244_),
    .c(_0215_),
    .y(_0247_)
  );
  al_and3 _1630_ (
    .a(_0246_),
    .b(_0214_),
    .c(_0247_),
    .y(_0248_)
  );
  al_ao21 _1631_ (
    .a(_0246_),
    .b(_0247_),
    .c(_0214_),
    .y(_0250_)
  );
  al_or3fft _1632_ (
    .a(_0213_),
    .b(_0250_),
    .c(_0248_),
    .y(_0251_)
  );
  al_oai21ftf _1633_ (
    .a(_0250_),
    .b(_0248_),
    .c(_0213_),
    .y(_0252_)
  );
  al_and3 _1634_ (
    .a(_0251_),
    .b(_0212_),
    .c(_0252_),
    .y(_0253_)
  );
  al_ao21 _1635_ (
    .a(_0251_),
    .b(_0252_),
    .c(_0212_),
    .y(_0254_)
  );
  al_or3fft _1636_ (
    .a(_0211_),
    .b(_0254_),
    .c(_0253_),
    .y(_0255_)
  );
  al_oai21ftf _1637_ (
    .a(_0254_),
    .b(_0253_),
    .c(_0211_),
    .y(_0256_)
  );
  al_and3 _1638_ (
    .a(_0255_),
    .b(_0210_),
    .c(_0256_),
    .y(_0257_)
  );
  al_ao21 _1639_ (
    .a(_0255_),
    .b(_0256_),
    .c(_0210_),
    .y(_0258_)
  );
  al_or3fft _1640_ (
    .a(_0209_),
    .b(_0258_),
    .c(_0257_),
    .y(_0259_)
  );
  al_oai21ftf _1641_ (
    .a(_0258_),
    .b(_0257_),
    .c(_0209_),
    .y(_0261_)
  );
  al_nand3 _1642_ (
    .a(_0259_),
    .b(_0261_),
    .c(_0208_),
    .y(_0262_)
  );
  al_ao21 _1643_ (
    .a(_0259_),
    .b(_0261_),
    .c(_0208_),
    .y(_0263_)
  );
  al_and3 _1644_ (
    .a(_0207_),
    .b(_0262_),
    .c(_0263_),
    .y(_0264_)
  );
  al_ao21 _1645_ (
    .a(_0262_),
    .b(_0263_),
    .c(_0207_),
    .y(_0265_)
  );
  al_and3ftt _1646_ (
    .a(_0264_),
    .b(_0265_),
    .c(_0206_),
    .y(_0266_)
  );
  al_ao21ftt _1647_ (
    .a(_0264_),
    .b(_0265_),
    .c(_0206_),
    .y(_0267_)
  );
  al_and2ft _1648_ (
    .a(_0266_),
    .b(_0267_),
    .y(_0268_)
  );
  al_nand2 _1649_ (
    .a(_0268_),
    .b(_0204_),
    .y(_0269_)
  );
  al_and3fft _1650_ (
    .a(_0199_),
    .b(_0268_),
    .c(_0202_),
    .y(_0270_)
  );
  al_nand2ft _1651_ (
    .a(_0270_),
    .b(_0269_),
    .y(N6200)
  );
  al_ao21 _1652_ (
    .a(_0268_),
    .b(_0204_),
    .c(_0266_),
    .y(_0272_)
  );
  al_ao21ttf _1653_ (
    .a(_0207_),
    .b(_0263_),
    .c(_0262_),
    .y(_0273_)
  );
  al_nand2 _1654_ (
    .a(N528),
    .b(N120),
    .y(_0274_)
  );
  al_ao21 _1655_ (
    .a(_0209_),
    .b(_0258_),
    .c(_0257_),
    .y(_0275_)
  );
  al_nand2 _1656_ (
    .a(N511),
    .b(N137),
    .y(_0276_)
  );
  al_ao21 _1657_ (
    .a(_0211_),
    .b(_0254_),
    .c(_0253_),
    .y(_0277_)
  );
  al_nand2 _1658_ (
    .a(N494),
    .b(N154),
    .y(_0278_)
  );
  al_ao21 _1659_ (
    .a(_0213_),
    .b(_0250_),
    .c(_0248_),
    .y(_0279_)
  );
  al_nand2 _1660_ (
    .a(N477),
    .b(N171),
    .y(_0280_)
  );
  al_ao21 _1661_ (
    .a(_0215_),
    .b(_0245_),
    .c(_0244_),
    .y(_0282_)
  );
  al_nand2 _1662_ (
    .a(N460),
    .b(N188),
    .y(_0283_)
  );
  al_ao21ttf _1663_ (
    .a(_0218_),
    .b(_0241_),
    .c(_0240_),
    .y(_0284_)
  );
  al_nand2 _1664_ (
    .a(N443),
    .b(N205),
    .y(_0285_)
  );
  al_ao21ttf _1665_ (
    .a(_0220_),
    .b(_0235_),
    .c(_0234_),
    .y(_0286_)
  );
  al_nand2 _1666_ (
    .a(N426),
    .b(N222),
    .y(_0287_)
  );
  al_ao21ttf _1667_ (
    .a(_0222_),
    .b(_0231_),
    .c(_0230_),
    .y(_0288_)
  );
  al_nand2 _1668_ (
    .a(N409),
    .b(N239),
    .y(_0289_)
  );
  al_nand2 _1669_ (
    .a(N392),
    .b(N256),
    .y(_0290_)
  );
  al_ao21ttf _1670_ (
    .a(_0226_),
    .b(_0228_),
    .c(_0290_),
    .y(_0291_)
  );
  al_nand3ftt _1671_ (
    .a(_0290_),
    .b(_0226_),
    .c(_0228_),
    .y(_0293_)
  );
  al_nand3 _1672_ (
    .a(_0289_),
    .b(_0293_),
    .c(_0291_),
    .y(_0294_)
  );
  al_ao21 _1673_ (
    .a(_0293_),
    .b(_0291_),
    .c(_0289_),
    .y(_0295_)
  );
  al_nand3 _1674_ (
    .a(_0294_),
    .b(_0295_),
    .c(_0288_),
    .y(_0296_)
  );
  al_ao21 _1675_ (
    .a(_0294_),
    .b(_0295_),
    .c(_0288_),
    .y(_0297_)
  );
  al_nand3 _1676_ (
    .a(_0287_),
    .b(_0296_),
    .c(_0297_),
    .y(_0298_)
  );
  al_ao21 _1677_ (
    .a(_0296_),
    .b(_0297_),
    .c(_0287_),
    .y(_0299_)
  );
  al_nand3 _1678_ (
    .a(_0298_),
    .b(_0299_),
    .c(_0286_),
    .y(_0300_)
  );
  al_ao21 _1679_ (
    .a(_0298_),
    .b(_0299_),
    .c(_0286_),
    .y(_0301_)
  );
  al_nand3 _1680_ (
    .a(_0285_),
    .b(_0300_),
    .c(_0301_),
    .y(_0302_)
  );
  al_ao21 _1681_ (
    .a(_0300_),
    .b(_0301_),
    .c(_0285_),
    .y(_0304_)
  );
  al_nand3 _1682_ (
    .a(_0302_),
    .b(_0304_),
    .c(_0284_),
    .y(_0305_)
  );
  al_ao21 _1683_ (
    .a(_0302_),
    .b(_0304_),
    .c(_0284_),
    .y(_0306_)
  );
  al_and3 _1684_ (
    .a(_0283_),
    .b(_0305_),
    .c(_0306_),
    .y(_0307_)
  );
  al_ao21 _1685_ (
    .a(_0305_),
    .b(_0306_),
    .c(_0283_),
    .y(_0308_)
  );
  al_nand3ftt _1686_ (
    .a(_0307_),
    .b(_0308_),
    .c(_0282_),
    .y(_0309_)
  );
  al_ao21ftt _1687_ (
    .a(_0307_),
    .b(_0308_),
    .c(_0282_),
    .y(_0310_)
  );
  al_and3 _1688_ (
    .a(_0280_),
    .b(_0309_),
    .c(_0310_),
    .y(_0311_)
  );
  al_ao21 _1689_ (
    .a(_0309_),
    .b(_0310_),
    .c(_0280_),
    .y(_0312_)
  );
  al_nand3ftt _1690_ (
    .a(_0311_),
    .b(_0312_),
    .c(_0279_),
    .y(_0313_)
  );
  al_ao21ftt _1691_ (
    .a(_0311_),
    .b(_0312_),
    .c(_0279_),
    .y(_0315_)
  );
  al_and3 _1692_ (
    .a(_0278_),
    .b(_0313_),
    .c(_0315_),
    .y(_0316_)
  );
  al_ao21 _1693_ (
    .a(_0313_),
    .b(_0315_),
    .c(_0278_),
    .y(_0317_)
  );
  al_nand3ftt _1694_ (
    .a(_0316_),
    .b(_0317_),
    .c(_0277_),
    .y(_0318_)
  );
  al_ao21ftt _1695_ (
    .a(_0316_),
    .b(_0317_),
    .c(_0277_),
    .y(_0319_)
  );
  al_and3 _1696_ (
    .a(_0276_),
    .b(_0318_),
    .c(_0319_),
    .y(_0320_)
  );
  al_ao21 _1697_ (
    .a(_0318_),
    .b(_0319_),
    .c(_0276_),
    .y(_0321_)
  );
  al_nand3ftt _1698_ (
    .a(_0320_),
    .b(_0321_),
    .c(_0275_),
    .y(_0322_)
  );
  al_ao21ftt _1699_ (
    .a(_0320_),
    .b(_0321_),
    .c(_0275_),
    .y(_0323_)
  );
  al_and3 _1700_ (
    .a(_0274_),
    .b(_0322_),
    .c(_0323_),
    .y(_0324_)
  );
  al_ao21 _1701_ (
    .a(_0322_),
    .b(_0323_),
    .c(_0274_),
    .y(_0326_)
  );
  al_and3ftt _1702_ (
    .a(_0324_),
    .b(_0326_),
    .c(_0273_),
    .y(_0327_)
  );
  al_ao21ftt _1703_ (
    .a(_0324_),
    .b(_0326_),
    .c(_0273_),
    .y(_0328_)
  );
  al_and2ft _1704_ (
    .a(_0327_),
    .b(_0328_),
    .y(_0329_)
  );
  al_nand2 _1705_ (
    .a(_0329_),
    .b(_0272_),
    .y(_0330_)
  );
  al_and3fft _1706_ (
    .a(_0266_),
    .b(_0329_),
    .c(_0269_),
    .y(_0331_)
  );
  al_nand2ft _1707_ (
    .a(_0331_),
    .b(_0330_),
    .y(N6210)
  );
  al_ao21 _1708_ (
    .a(_0329_),
    .b(_0272_),
    .c(_0327_),
    .y(_0332_)
  );
  al_ao21ttf _1709_ (
    .a(_0274_),
    .b(_0323_),
    .c(_0322_),
    .y(_0333_)
  );
  al_nand2 _1710_ (
    .a(N528),
    .b(N137),
    .y(_0334_)
  );
  al_aoi21ttf _1711_ (
    .a(_0276_),
    .b(_0319_),
    .c(_0318_),
    .y(_0336_)
  );
  al_nand2 _1712_ (
    .a(N511),
    .b(N154),
    .y(_0337_)
  );
  al_aoi21ttf _1713_ (
    .a(_0278_),
    .b(_0315_),
    .c(_0313_),
    .y(_0338_)
  );
  al_nand2 _1714_ (
    .a(N494),
    .b(N171),
    .y(_0339_)
  );
  al_aoi21ttf _1715_ (
    .a(_0280_),
    .b(_0310_),
    .c(_0309_),
    .y(_0340_)
  );
  al_nand2 _1716_ (
    .a(N477),
    .b(N188),
    .y(_0341_)
  );
  al_ao21ttf _1717_ (
    .a(_0283_),
    .b(_0306_),
    .c(_0305_),
    .y(_0342_)
  );
  al_nand2 _1718_ (
    .a(N460),
    .b(N205),
    .y(_0343_)
  );
  al_ao21ttf _1719_ (
    .a(_0285_),
    .b(_0301_),
    .c(_0300_),
    .y(_0344_)
  );
  al_nand2 _1720_ (
    .a(N443),
    .b(N222),
    .y(_0345_)
  );
  al_ao21ttf _1721_ (
    .a(_0287_),
    .b(_0297_),
    .c(_0296_),
    .y(_0347_)
  );
  al_nand2 _1722_ (
    .a(N426),
    .b(N239),
    .y(_0348_)
  );
  al_nand2 _1723_ (
    .a(N409),
    .b(N256),
    .y(_0349_)
  );
  al_ao21ttf _1724_ (
    .a(_0291_),
    .b(_0294_),
    .c(_0349_),
    .y(_0350_)
  );
  al_nand3ftt _1725_ (
    .a(_0349_),
    .b(_0291_),
    .c(_0294_),
    .y(_0351_)
  );
  al_and3 _1726_ (
    .a(_0348_),
    .b(_0351_),
    .c(_0350_),
    .y(_0352_)
  );
  al_ao21 _1727_ (
    .a(_0351_),
    .b(_0350_),
    .c(_0348_),
    .y(_0353_)
  );
  al_nand3ftt _1728_ (
    .a(_0352_),
    .b(_0353_),
    .c(_0347_),
    .y(_0354_)
  );
  al_ao21ftt _1729_ (
    .a(_0352_),
    .b(_0353_),
    .c(_0347_),
    .y(_0355_)
  );
  al_nand3 _1730_ (
    .a(_0345_),
    .b(_0354_),
    .c(_0355_),
    .y(_0356_)
  );
  al_ao21 _1731_ (
    .a(_0354_),
    .b(_0355_),
    .c(_0345_),
    .y(_0358_)
  );
  al_and3 _1732_ (
    .a(_0356_),
    .b(_0358_),
    .c(_0344_),
    .y(_0359_)
  );
  al_ao21 _1733_ (
    .a(_0356_),
    .b(_0358_),
    .c(_0344_),
    .y(_0360_)
  );
  al_or3fft _1734_ (
    .a(_0343_),
    .b(_0360_),
    .c(_0359_),
    .y(_0361_)
  );
  al_oai21ftf _1735_ (
    .a(_0360_),
    .b(_0359_),
    .c(_0343_),
    .y(_0362_)
  );
  al_and3 _1736_ (
    .a(_0361_),
    .b(_0362_),
    .c(_0342_),
    .y(_0363_)
  );
  al_ao21 _1737_ (
    .a(_0361_),
    .b(_0362_),
    .c(_0342_),
    .y(_0364_)
  );
  al_nor3fft _1738_ (
    .a(_0341_),
    .b(_0364_),
    .c(_0363_),
    .y(_0365_)
  );
  al_oai21ftf _1739_ (
    .a(_0364_),
    .b(_0363_),
    .c(_0341_),
    .y(_0366_)
  );
  al_and3fft _1740_ (
    .a(_0365_),
    .b(_0340_),
    .c(_0366_),
    .y(_0367_)
  );
  al_ao21ftf _1741_ (
    .a(_0365_),
    .b(_0366_),
    .c(_0340_),
    .y(_0369_)
  );
  al_nor3fft _1742_ (
    .a(_0339_),
    .b(_0369_),
    .c(_0367_),
    .y(_0370_)
  );
  al_oai21ftf _1743_ (
    .a(_0369_),
    .b(_0367_),
    .c(_0339_),
    .y(_0371_)
  );
  al_and3fft _1744_ (
    .a(_0370_),
    .b(_0338_),
    .c(_0371_),
    .y(_0372_)
  );
  al_ao21ftf _1745_ (
    .a(_0370_),
    .b(_0371_),
    .c(_0338_),
    .y(_0373_)
  );
  al_nor3fft _1746_ (
    .a(_0337_),
    .b(_0373_),
    .c(_0372_),
    .y(_0374_)
  );
  al_oai21ftf _1747_ (
    .a(_0373_),
    .b(_0372_),
    .c(_0337_),
    .y(_0375_)
  );
  al_and3fft _1748_ (
    .a(_0374_),
    .b(_0336_),
    .c(_0375_),
    .y(_0376_)
  );
  al_ao21ftf _1749_ (
    .a(_0374_),
    .b(_0375_),
    .c(_0336_),
    .y(_0377_)
  );
  al_nor3fft _1750_ (
    .a(_0334_),
    .b(_0377_),
    .c(_0376_),
    .y(_0378_)
  );
  al_oai21ftf _1751_ (
    .a(_0377_),
    .b(_0376_),
    .c(_0334_),
    .y(_0380_)
  );
  al_and3ftt _1752_ (
    .a(_0378_),
    .b(_0333_),
    .c(_0380_),
    .y(_0381_)
  );
  al_ao21ftt _1753_ (
    .a(_0378_),
    .b(_0380_),
    .c(_0333_),
    .y(_0382_)
  );
  al_and2ft _1754_ (
    .a(_0381_),
    .b(_0382_),
    .y(_0383_)
  );
  al_and2 _1755_ (
    .a(_0383_),
    .b(_0332_),
    .y(_0384_)
  );
  al_and3fft _1756_ (
    .a(_0327_),
    .b(_0383_),
    .c(_0330_),
    .y(_0385_)
  );
  al_or2 _1757_ (
    .a(_0385_),
    .b(_0384_),
    .y(N6220)
  );
  al_ao21 _1758_ (
    .a(_0383_),
    .b(_0332_),
    .c(_0381_),
    .y(_0386_)
  );
  al_ao21 _1759_ (
    .a(_0334_),
    .b(_0377_),
    .c(_0376_),
    .y(_0387_)
  );
  al_nand2 _1760_ (
    .a(N528),
    .b(N154),
    .y(_0388_)
  );
  al_ao21 _1761_ (
    .a(_0337_),
    .b(_0373_),
    .c(_0372_),
    .y(_0390_)
  );
  al_nand2 _1762_ (
    .a(N511),
    .b(N171),
    .y(_0391_)
  );
  al_ao21 _1763_ (
    .a(_0339_),
    .b(_0369_),
    .c(_0367_),
    .y(_0392_)
  );
  al_nand2 _1764_ (
    .a(N494),
    .b(N188),
    .y(_0393_)
  );
  al_ao21 _1765_ (
    .a(_0341_),
    .b(_0364_),
    .c(_0363_),
    .y(_0394_)
  );
  al_nand2 _1766_ (
    .a(N477),
    .b(N205),
    .y(_0395_)
  );
  al_ao21 _1767_ (
    .a(_0343_),
    .b(_0360_),
    .c(_0359_),
    .y(_0396_)
  );
  al_nand2 _1768_ (
    .a(N460),
    .b(N222),
    .y(_0397_)
  );
  al_ao21ttf _1769_ (
    .a(_0345_),
    .b(_0355_),
    .c(_0354_),
    .y(_0398_)
  );
  al_ao21ttf _1770_ (
    .a(_0348_),
    .b(_0351_),
    .c(_0350_),
    .y(_0399_)
  );
  al_ao21ftf _1771_ (
    .a(_1344_),
    .b(N426),
    .c(_0399_),
    .y(_0401_)
  );
  al_and3fft _1772_ (
    .a(_1344_),
    .b(_0399_),
    .c(N426),
    .y(_0402_)
  );
  al_nor2ft _1773_ (
    .a(_0401_),
    .b(_0402_),
    .y(_0403_)
  );
  al_ao21ftf _1774_ (
    .a(_0074_),
    .b(N443),
    .c(_0403_),
    .y(_0404_)
  );
  al_and3fft _1775_ (
    .a(_0074_),
    .b(_0403_),
    .c(N443),
    .y(_0405_)
  );
  al_or3fft _1776_ (
    .a(_0398_),
    .b(_0404_),
    .c(_0405_),
    .y(_0406_)
  );
  al_oai21ftf _1777_ (
    .a(_0404_),
    .b(_0405_),
    .c(_0398_),
    .y(_0407_)
  );
  al_nand3 _1778_ (
    .a(_0397_),
    .b(_0406_),
    .c(_0407_),
    .y(_0408_)
  );
  al_ao21 _1779_ (
    .a(_0406_),
    .b(_0407_),
    .c(_0397_),
    .y(_0409_)
  );
  al_and3 _1780_ (
    .a(_0396_),
    .b(_0408_),
    .c(_0409_),
    .y(_0410_)
  );
  al_ao21 _1781_ (
    .a(_0408_),
    .b(_0409_),
    .c(_0396_),
    .y(_0412_)
  );
  al_or3fft _1782_ (
    .a(_0395_),
    .b(_0412_),
    .c(_0410_),
    .y(_0413_)
  );
  al_ao21ftt _1783_ (
    .a(_0410_),
    .b(_0412_),
    .c(_0395_),
    .y(_0414_)
  );
  al_and3 _1784_ (
    .a(_0394_),
    .b(_0413_),
    .c(_0414_),
    .y(_0415_)
  );
  al_ao21 _1785_ (
    .a(_0413_),
    .b(_0414_),
    .c(_0394_),
    .y(_0416_)
  );
  al_nor3fft _1786_ (
    .a(_0393_),
    .b(_0416_),
    .c(_0415_),
    .y(_0417_)
  );
  al_ao21ftt _1787_ (
    .a(_0415_),
    .b(_0416_),
    .c(_0393_),
    .y(_0418_)
  );
  al_nor3fft _1788_ (
    .a(_0392_),
    .b(_0418_),
    .c(_0417_),
    .y(_0419_)
  );
  al_ao21ftt _1789_ (
    .a(_0417_),
    .b(_0418_),
    .c(_0392_),
    .y(_0420_)
  );
  al_nor3fft _1790_ (
    .a(_0391_),
    .b(_0420_),
    .c(_0419_),
    .y(_0421_)
  );
  al_ao21ftt _1791_ (
    .a(_0419_),
    .b(_0420_),
    .c(_0391_),
    .y(_0423_)
  );
  al_nor3fft _1792_ (
    .a(_0390_),
    .b(_0423_),
    .c(_0421_),
    .y(_0424_)
  );
  al_ao21ftt _1793_ (
    .a(_0421_),
    .b(_0423_),
    .c(_0390_),
    .y(_0425_)
  );
  al_nor3fft _1794_ (
    .a(_0388_),
    .b(_0425_),
    .c(_0424_),
    .y(_0426_)
  );
  al_ao21ftt _1795_ (
    .a(_0424_),
    .b(_0425_),
    .c(_0388_),
    .y(_0427_)
  );
  al_nor3fft _1796_ (
    .a(_0387_),
    .b(_0427_),
    .c(_0426_),
    .y(_0428_)
  );
  al_ao21ftt _1797_ (
    .a(_0426_),
    .b(_0427_),
    .c(_0387_),
    .y(_0429_)
  );
  al_and2ft _1798_ (
    .a(_0428_),
    .b(_0429_),
    .y(_0430_)
  );
  al_nand2 _1799_ (
    .a(_0430_),
    .b(_0386_),
    .y(_0431_)
  );
  al_or3 _1800_ (
    .a(_0381_),
    .b(_0430_),
    .c(_0384_),
    .y(_0432_)
  );
  al_nand2 _1801_ (
    .a(_0432_),
    .b(_0431_),
    .y(N6230)
  );
  al_inv _1802_ (
    .a(_0428_),
    .y(_0434_)
  );
  al_ao21 _1803_ (
    .a(_0388_),
    .b(_0425_),
    .c(_0424_),
    .y(_0435_)
  );
  al_nand2 _1804_ (
    .a(N528),
    .b(N171),
    .y(_0436_)
  );
  al_aoi21 _1805_ (
    .a(_0391_),
    .b(_0420_),
    .c(_0419_),
    .y(_0437_)
  );
  al_nand2 _1806_ (
    .a(N511),
    .b(N188),
    .y(_0438_)
  );
  al_ao21 _1807_ (
    .a(_0393_),
    .b(_0416_),
    .c(_0415_),
    .y(_0439_)
  );
  al_nand2 _1808_ (
    .a(N494),
    .b(N205),
    .y(_0440_)
  );
  al_ao21 _1809_ (
    .a(_0395_),
    .b(_0412_),
    .c(_0410_),
    .y(_0441_)
  );
  al_nand2 _1810_ (
    .a(N477),
    .b(N222),
    .y(_0442_)
  );
  al_ao21ttf _1811_ (
    .a(_0397_),
    .b(_0407_),
    .c(_0406_),
    .y(_0444_)
  );
  al_nand2 _1812_ (
    .a(_0401_),
    .b(_0404_),
    .y(_0445_)
  );
  al_ao21ftf _1813_ (
    .a(_1344_),
    .b(N443),
    .c(_0445_),
    .y(_0446_)
  );
  al_and3fft _1814_ (
    .a(_1344_),
    .b(_0445_),
    .c(N443),
    .y(_0447_)
  );
  al_nor2ft _1815_ (
    .a(_0446_),
    .b(_0447_),
    .y(_0448_)
  );
  al_ao21ftf _1816_ (
    .a(_0074_),
    .b(N460),
    .c(_0448_),
    .y(_0449_)
  );
  al_and3fft _1817_ (
    .a(_0074_),
    .b(_0448_),
    .c(N460),
    .y(_0450_)
  );
  al_or3fft _1818_ (
    .a(_0444_),
    .b(_0449_),
    .c(_0450_),
    .y(_0451_)
  );
  al_oai21ftf _1819_ (
    .a(_0449_),
    .b(_0450_),
    .c(_0444_),
    .y(_0452_)
  );
  al_nand3 _1820_ (
    .a(_0442_),
    .b(_0451_),
    .c(_0452_),
    .y(_0453_)
  );
  al_ao21 _1821_ (
    .a(_0451_),
    .b(_0452_),
    .c(_0442_),
    .y(_0455_)
  );
  al_nand3 _1822_ (
    .a(_0441_),
    .b(_0453_),
    .c(_0455_),
    .y(_0456_)
  );
  al_ao21 _1823_ (
    .a(_0453_),
    .b(_0455_),
    .c(_0441_),
    .y(_0457_)
  );
  al_nand3 _1824_ (
    .a(_0440_),
    .b(_0456_),
    .c(_0457_),
    .y(_0458_)
  );
  al_ao21 _1825_ (
    .a(_0456_),
    .b(_0457_),
    .c(_0440_),
    .y(_0459_)
  );
  al_and3 _1826_ (
    .a(_0439_),
    .b(_0458_),
    .c(_0459_),
    .y(_0460_)
  );
  al_ao21 _1827_ (
    .a(_0458_),
    .b(_0459_),
    .c(_0439_),
    .y(_0461_)
  );
  al_nor3fft _1828_ (
    .a(_0438_),
    .b(_0461_),
    .c(_0460_),
    .y(_0462_)
  );
  al_ao21ftt _1829_ (
    .a(_0460_),
    .b(_0461_),
    .c(_0438_),
    .y(_0463_)
  );
  al_and3fft _1830_ (
    .a(_0437_),
    .b(_0462_),
    .c(_0463_),
    .y(_0464_)
  );
  al_oai21ftt _1831_ (
    .a(_0463_),
    .b(_0462_),
    .c(_0437_),
    .y(_0466_)
  );
  al_or3fft _1832_ (
    .a(_0436_),
    .b(_0466_),
    .c(_0464_),
    .y(_0467_)
  );
  al_ao21ftt _1833_ (
    .a(_0464_),
    .b(_0466_),
    .c(_0436_),
    .y(_0468_)
  );
  al_and3 _1834_ (
    .a(_0435_),
    .b(_0467_),
    .c(_0468_),
    .y(_0469_)
  );
  al_ao21 _1835_ (
    .a(_0467_),
    .b(_0468_),
    .c(_0435_),
    .y(_0470_)
  );
  al_nand2ft _1836_ (
    .a(_0469_),
    .b(_0470_),
    .y(_0471_)
  );
  al_ao21 _1837_ (
    .a(_0434_),
    .b(_0431_),
    .c(_0471_),
    .y(_0472_)
  );
  al_and3 _1838_ (
    .a(_0434_),
    .b(_0471_),
    .c(_0431_),
    .y(_0473_)
  );
  al_nand2ft _1839_ (
    .a(_0473_),
    .b(_0472_),
    .y(N6240)
  );
  al_inv _1840_ (
    .a(_0469_),
    .y(_0474_)
  );
  al_ao21 _1841_ (
    .a(_0436_),
    .b(_0466_),
    .c(_0464_),
    .y(_0475_)
  );
  al_nand2 _1842_ (
    .a(N528),
    .b(N188),
    .y(_0476_)
  );
  al_ao21 _1843_ (
    .a(_0438_),
    .b(_0461_),
    .c(_0460_),
    .y(_0477_)
  );
  al_nand2 _1844_ (
    .a(N511),
    .b(N205),
    .y(_0478_)
  );
  al_ao21ttf _1845_ (
    .a(_0440_),
    .b(_0457_),
    .c(_0456_),
    .y(_0479_)
  );
  al_nand2 _1846_ (
    .a(N494),
    .b(N222),
    .y(_0480_)
  );
  al_ao21ttf _1847_ (
    .a(_0442_),
    .b(_0452_),
    .c(_0451_),
    .y(_0481_)
  );
  al_nand2 _1848_ (
    .a(N477),
    .b(N239),
    .y(_0482_)
  );
  al_nand2 _1849_ (
    .a(N460),
    .b(N256),
    .y(_0483_)
  );
  al_ao21ttf _1850_ (
    .a(_0446_),
    .b(_0449_),
    .c(_0483_),
    .y(_0484_)
  );
  al_nand3ftt _1851_ (
    .a(_0483_),
    .b(_0446_),
    .c(_0449_),
    .y(_0486_)
  );
  al_nand3 _1852_ (
    .a(_0482_),
    .b(_0486_),
    .c(_0484_),
    .y(_0487_)
  );
  al_ao21 _1853_ (
    .a(_0486_),
    .b(_0484_),
    .c(_0482_),
    .y(_0488_)
  );
  al_nand3 _1854_ (
    .a(_0487_),
    .b(_0488_),
    .c(_0481_),
    .y(_0489_)
  );
  al_ao21 _1855_ (
    .a(_0487_),
    .b(_0488_),
    .c(_0481_),
    .y(_0490_)
  );
  al_and3 _1856_ (
    .a(_0480_),
    .b(_0489_),
    .c(_0490_),
    .y(_0491_)
  );
  al_ao21 _1857_ (
    .a(_0489_),
    .b(_0490_),
    .c(_0480_),
    .y(_0492_)
  );
  al_nand3ftt _1858_ (
    .a(_0491_),
    .b(_0492_),
    .c(_0479_),
    .y(_0493_)
  );
  al_ao21ftt _1859_ (
    .a(_0491_),
    .b(_0492_),
    .c(_0479_),
    .y(_0494_)
  );
  al_nand3 _1860_ (
    .a(_0478_),
    .b(_0493_),
    .c(_0494_),
    .y(_0495_)
  );
  al_ao21 _1861_ (
    .a(_0493_),
    .b(_0494_),
    .c(_0478_),
    .y(_0497_)
  );
  al_and3 _1862_ (
    .a(_0495_),
    .b(_0477_),
    .c(_0497_),
    .y(_0498_)
  );
  al_ao21 _1863_ (
    .a(_0495_),
    .b(_0497_),
    .c(_0477_),
    .y(_0499_)
  );
  al_nor3fft _1864_ (
    .a(_0476_),
    .b(_0499_),
    .c(_0498_),
    .y(_0500_)
  );
  al_oai21ftf _1865_ (
    .a(_0499_),
    .b(_0498_),
    .c(_0476_),
    .y(_0501_)
  );
  al_and3ftt _1866_ (
    .a(_0500_),
    .b(_0475_),
    .c(_0501_),
    .y(_0502_)
  );
  al_ao21ftt _1867_ (
    .a(_0500_),
    .b(_0501_),
    .c(_0475_),
    .y(_0503_)
  );
  al_nand2ft _1868_ (
    .a(_0502_),
    .b(_0503_),
    .y(_0504_)
  );
  al_ao21 _1869_ (
    .a(_0474_),
    .b(_0472_),
    .c(_0504_),
    .y(_0505_)
  );
  al_and3 _1870_ (
    .a(_0474_),
    .b(_0504_),
    .c(_0472_),
    .y(_0506_)
  );
  al_nand2ft _1871_ (
    .a(_0506_),
    .b(_0505_),
    .y(N6250)
  );
  al_inv _1872_ (
    .a(_0502_),
    .y(_0508_)
  );
  al_ao21 _1873_ (
    .a(_0476_),
    .b(_0499_),
    .c(_0498_),
    .y(_0509_)
  );
  al_nand2 _1874_ (
    .a(N528),
    .b(N205),
    .y(_0510_)
  );
  al_ao21ttf _1875_ (
    .a(_0478_),
    .b(_0494_),
    .c(_0493_),
    .y(_0511_)
  );
  al_nand2 _1876_ (
    .a(N511),
    .b(N222),
    .y(_0512_)
  );
  al_ao21ttf _1877_ (
    .a(_0480_),
    .b(_0490_),
    .c(_0489_),
    .y(_0513_)
  );
  al_nand2 _1878_ (
    .a(N494),
    .b(N239),
    .y(_0514_)
  );
  al_nand2 _1879_ (
    .a(N477),
    .b(N256),
    .y(_0515_)
  );
  al_ao21ttf _1880_ (
    .a(_0484_),
    .b(_0487_),
    .c(_0515_),
    .y(_0516_)
  );
  al_nand3ftt _1881_ (
    .a(_0515_),
    .b(_0484_),
    .c(_0487_),
    .y(_0518_)
  );
  al_and3 _1882_ (
    .a(_0514_),
    .b(_0518_),
    .c(_0516_),
    .y(_0519_)
  );
  al_ao21 _1883_ (
    .a(_0518_),
    .b(_0516_),
    .c(_0514_),
    .y(_0520_)
  );
  al_nand3ftt _1884_ (
    .a(_0519_),
    .b(_0520_),
    .c(_0513_),
    .y(_0521_)
  );
  al_ao21ftt _1885_ (
    .a(_0519_),
    .b(_0520_),
    .c(_0513_),
    .y(_0522_)
  );
  al_and3 _1886_ (
    .a(_0512_),
    .b(_0521_),
    .c(_0522_),
    .y(_0523_)
  );
  al_ao21 _1887_ (
    .a(_0521_),
    .b(_0522_),
    .c(_0512_),
    .y(_0524_)
  );
  al_nand3ftt _1888_ (
    .a(_0523_),
    .b(_0524_),
    .c(_0511_),
    .y(_0525_)
  );
  al_ao21ftt _1889_ (
    .a(_0523_),
    .b(_0524_),
    .c(_0511_),
    .y(_0526_)
  );
  al_nand3 _1890_ (
    .a(_0510_),
    .b(_0525_),
    .c(_0526_),
    .y(_0527_)
  );
  al_ao21 _1891_ (
    .a(_0525_),
    .b(_0526_),
    .c(_0510_),
    .y(_0529_)
  );
  al_and3 _1892_ (
    .a(_0527_),
    .b(_0529_),
    .c(_0509_),
    .y(_0530_)
  );
  al_ao21 _1893_ (
    .a(_0527_),
    .b(_0529_),
    .c(_0509_),
    .y(_0531_)
  );
  al_nand2ft _1894_ (
    .a(_0530_),
    .b(_0531_),
    .y(_0532_)
  );
  al_ao21 _1895_ (
    .a(_0508_),
    .b(_0505_),
    .c(_0532_),
    .y(_0533_)
  );
  al_and3 _1896_ (
    .a(_0508_),
    .b(_0532_),
    .c(_0505_),
    .y(_0534_)
  );
  al_nand2ft _1897_ (
    .a(_0534_),
    .b(_0533_),
    .y(N6260)
  );
  al_inv _1898_ (
    .a(_0530_),
    .y(_0535_)
  );
  al_ao21ttf _1899_ (
    .a(_0510_),
    .b(_0526_),
    .c(_0525_),
    .y(_0536_)
  );
  al_nand2 _1900_ (
    .a(N528),
    .b(N222),
    .y(_0537_)
  );
  al_nand2 _1901_ (
    .a(N511),
    .b(N239),
    .y(_0539_)
  );
  al_ao21ttf _1902_ (
    .a(_0514_),
    .b(_0518_),
    .c(_0516_),
    .y(_0540_)
  );
  al_ao21ftf _1903_ (
    .a(_1344_),
    .b(N494),
    .c(_0540_),
    .y(_0541_)
  );
  al_or3fft _1904_ (
    .a(N494),
    .b(N256),
    .c(_0540_),
    .y(_0542_)
  );
  al_and3 _1905_ (
    .a(_0539_),
    .b(_0541_),
    .c(_0542_),
    .y(_0543_)
  );
  al_ao21 _1906_ (
    .a(_0541_),
    .b(_0542_),
    .c(_0539_),
    .y(_0544_)
  );
  al_nand2ft _1907_ (
    .a(_0543_),
    .b(_0544_),
    .y(_0545_)
  );
  al_ao21ftt _1908_ (
    .a(_0523_),
    .b(_0521_),
    .c(_0545_),
    .y(_0546_)
  );
  al_nand3ftt _1909_ (
    .a(_0523_),
    .b(_0521_),
    .c(_0545_),
    .y(_0547_)
  );
  al_and3 _1910_ (
    .a(_0537_),
    .b(_0547_),
    .c(_0546_),
    .y(_0548_)
  );
  al_ao21 _1911_ (
    .a(_0547_),
    .b(_0546_),
    .c(_0537_),
    .y(_0550_)
  );
  al_or3fft _1912_ (
    .a(_0536_),
    .b(_0550_),
    .c(_0548_),
    .y(_0551_)
  );
  al_aoi21ftt _1913_ (
    .a(_0548_),
    .b(_0550_),
    .c(_0536_),
    .y(_0552_)
  );
  al_or2ft _1914_ (
    .a(_0551_),
    .b(_0552_),
    .y(_0553_)
  );
  al_ao21 _1915_ (
    .a(_0535_),
    .b(_0533_),
    .c(_0553_),
    .y(_0554_)
  );
  al_and3 _1916_ (
    .a(_0535_),
    .b(_0553_),
    .c(_0533_),
    .y(_0555_)
  );
  al_nand2ft _1917_ (
    .a(_0555_),
    .b(_0554_),
    .y(N6270)
  );
  al_ao21ttf _1918_ (
    .a(_0537_),
    .b(_0547_),
    .c(_0546_),
    .y(_0556_)
  );
  al_ao21ttf _1919_ (
    .a(_0539_),
    .b(_0542_),
    .c(_0541_),
    .y(_0557_)
  );
  al_ao21ftf _1920_ (
    .a(_1344_),
    .b(N511),
    .c(_0557_),
    .y(_0558_)
  );
  al_and3fft _1921_ (
    .a(_1344_),
    .b(_0557_),
    .c(N511),
    .y(_0560_)
  );
  al_nor2ft _1922_ (
    .a(_0558_),
    .b(_0560_),
    .y(_0561_)
  );
  al_ao21ftf _1923_ (
    .a(_0074_),
    .b(N528),
    .c(_0561_),
    .y(_0562_)
  );
  al_and3fft _1924_ (
    .a(_0074_),
    .b(_0561_),
    .c(N528),
    .y(_0563_)
  );
  al_or3fft _1925_ (
    .a(_0562_),
    .b(_0556_),
    .c(_0563_),
    .y(_0564_)
  );
  al_oa21ftf _1926_ (
    .a(_0562_),
    .b(_0563_),
    .c(_0556_),
    .y(_0565_)
  );
  al_nand2ft _1927_ (
    .a(_0565_),
    .b(_0564_),
    .y(_0566_)
  );
  al_ao21 _1928_ (
    .a(_0551_),
    .b(_0554_),
    .c(_0566_),
    .y(_0567_)
  );
  al_and3 _1929_ (
    .a(_0551_),
    .b(_0566_),
    .c(_0554_),
    .y(_0568_)
  );
  al_nand2ft _1930_ (
    .a(_0568_),
    .b(_0567_),
    .y(N6280)
  );
  al_nand2 _1931_ (
    .a(_0558_),
    .b(_0562_),
    .y(_0570_)
  );
  al_ao21ftf _1932_ (
    .a(_1344_),
    .b(N528),
    .c(_0570_),
    .y(_0571_)
  );
  al_and3fft _1933_ (
    .a(_1344_),
    .b(_0570_),
    .c(N528),
    .y(_0572_)
  );
  al_or2ft _1934_ (
    .a(_0571_),
    .b(_0572_),
    .y(_0573_)
  );
  al_ao21 _1935_ (
    .a(_0564_),
    .b(_0567_),
    .c(_0573_),
    .y(_0574_)
  );
  al_and2 _1936_ (
    .a(_0571_),
    .b(_0574_),
    .y(N6287)
  );
  al_and3 _1937_ (
    .a(_0564_),
    .b(_0573_),
    .c(_0567_),
    .y(_0575_)
  );
  al_nand2ft _1938_ (
    .a(_0575_),
    .b(_0574_),
    .y(N6288)
  );
  al_inv _1939_ (
    .a(_1076_),
    .y(N545)
  );
  al_nor3fft _1940_ (
    .a(_1312_),
    .b(_1313_),
    .c(_1220_),
    .y(_0576_)
  );
  al_nor2ft _1941_ (
    .a(_1315_),
    .b(_0576_),
    .y(N6150)
  );
  al_and2 _1942_ (
    .a(N290),
    .b(N18),
    .y(_1065_)
  );
  al_nand2 _1943_ (
    .a(N1),
    .b(N273),
    .y(_1076_)
  );
  al_and2 _1944_ (
    .a(N273),
    .b(N18),
    .y(_1087_)
  );
  al_ao21 _1945_ (
    .a(N1),
    .b(N290),
    .c(_1087_),
    .y(_1098_)
  );
  al_aoi21ftf _1946_ (
    .a(_1076_),
    .b(_1065_),
    .c(_1098_),
    .y(N1581)
  );
  al_and3 _1947_ (
    .a(N1),
    .b(N273),
    .c(_1065_),
    .y(_1118_)
  );
  al_and3 _1948_ (
    .a(N290),
    .b(N35),
    .c(_1087_),
    .y(_1129_)
  );
  al_ao21 _1949_ (
    .a(N273),
    .b(N35),
    .c(_1065_),
    .y(_1140_)
  );
  al_oai21ftf _1950_ (
    .a(_1140_),
    .b(_1129_),
    .c(_1118_),
    .y(_1151_)
  );
  al_and2 _1951_ (
    .a(N273),
    .b(N35),
    .y(_1162_)
  );
  al_and3fft _1952_ (
    .a(_1076_),
    .b(_1162_),
    .c(_1065_),
    .y(_1173_)
  );
  al_and2ft _1953_ (
    .a(_1173_),
    .b(_1151_),
    .y(_1184_)
  );
  al_aoi21ttf _1954_ (
    .a(N1),
    .b(N307),
    .c(_1184_),
    .y(_1195_)
  );
  al_or3fft _1955_ (
    .a(N1),
    .b(N307),
    .c(_1184_),
    .y(_1206_)
  );
  al_nand2ft _1956_ (
    .a(_1195_),
    .b(_1206_),
    .y(N1901)
  );
  al_nand2 _1957_ (
    .a(N1),
    .b(N324),
    .y(_1226_)
  );
  al_nand2 _1958_ (
    .a(N307),
    .b(N18),
    .y(_1237_)
  );
  al_and3 _1959_ (
    .a(N290),
    .b(N52),
    .c(_1162_),
    .y(_1248_)
  );
  al_nand2 _1960_ (
    .a(N290),
    .b(N35),
    .y(_1259_)
  );
  al_ao21ttf _1961_ (
    .a(N273),
    .b(N52),
    .c(_1259_),
    .y(_1270_)
  );
  al_oai21ftf _1962_ (
    .a(_1270_),
    .b(_1248_),
    .c(_1129_),
    .y(_1281_)
  );
  al_or3fft _1963_ (
    .a(_1270_),
    .b(_1129_),
    .c(_1248_),
    .y(_1292_)
  );
  al_and3 _1964_ (
    .a(_1237_),
    .b(_1281_),
    .c(_1292_),
    .y(_1303_)
  );
  al_ao21 _1965_ (
    .a(_1281_),
    .b(_1292_),
    .c(_1237_),
    .y(_1314_)
  );
  al_nand2ft _1966_ (
    .a(_1303_),
    .b(_1314_),
    .y(_1325_)
  );
  al_aoi21ftt _1967_ (
    .a(_1195_),
    .b(_1151_),
    .c(_1325_),
    .y(_1336_)
  );
  al_nand3ftt _1968_ (
    .a(_1195_),
    .b(_1151_),
    .c(_1325_),
    .y(_1347_)
  );
  al_nor3fft _1969_ (
    .a(_1226_),
    .b(_1347_),
    .c(_1336_),
    .y(_1358_)
  );
  al_oai21ftf _1970_ (
    .a(_1347_),
    .b(_1336_),
    .c(_1226_),
    .y(_1369_)
  );
  al_nand2ft _1971_ (
    .a(_1358_),
    .b(_1369_),
    .y(N2223)
  );
  al_nand2 _1972_ (
    .a(N1),
    .b(N341),
    .y(_1390_)
  );
  al_ao21 _1973_ (
    .a(_1226_),
    .b(_1347_),
    .c(_1336_),
    .y(_1401_)
  );
  al_nand2 _1974_ (
    .a(N324),
    .b(N18),
    .y(_1411_)
  );
  al_ao21ttf _1975_ (
    .a(_1237_),
    .b(_1292_),
    .c(_1281_),
    .y(_1422_)
  );
  al_nand2 _1976_ (
    .a(N307),
    .b(N35),
    .y(_1433_)
  );
  al_and2 _1977_ (
    .a(N273),
    .b(N52),
    .y(_0000_)
  );
  al_and3 _1978_ (
    .a(N290),
    .b(N69),
    .c(_0000_),
    .y(_0011_)
  );
  al_nand2 _1979_ (
    .a(N290),
    .b(N52),
    .y(_0022_)
  );
  al_ao21ttf _1980_ (
    .a(N273),
    .b(N69),
    .c(_0022_),
    .y(_0033_)
  );
  al_oai21ftf _1981_ (
    .a(_0033_),
    .b(_0011_),
    .c(_1248_),
    .y(_0044_)
  );
  al_or3fft _1982_ (
    .a(_0033_),
    .b(_1248_),
    .c(_0011_),
    .y(_0054_)
  );
  al_and3 _1983_ (
    .a(_1433_),
    .b(_0044_),
    .c(_0054_),
    .y(_0065_)
  );
  al_ao21 _1984_ (
    .a(_0044_),
    .b(_0054_),
    .c(_1433_),
    .y(_0076_)
  );
  al_nand3ftt _1985_ (
    .a(_0065_),
    .b(_1422_),
    .c(_0076_),
    .y(_0087_)
  );
  al_ao21ftt _1986_ (
    .a(_0065_),
    .b(_0076_),
    .c(_1422_),
    .y(_0098_)
  );
  al_and3 _1987_ (
    .a(_1411_),
    .b(_0087_),
    .c(_0098_),
    .y(_0109_)
  );
  al_ao21 _1988_ (
    .a(_0087_),
    .b(_0098_),
    .c(_1411_),
    .y(_0120_)
  );
  al_and3ftt _1989_ (
    .a(_0109_),
    .b(_0120_),
    .c(_1401_),
    .y(_0131_)
  );
  al_ao21ftt _1990_ (
    .a(_0109_),
    .b(_0120_),
    .c(_1401_),
    .y(_0141_)
  );
  al_nor3fft _1991_ (
    .a(_1390_),
    .b(_0141_),
    .c(_0131_),
    .y(_0152_)
  );
  al_oai21ftf _1992_ (
    .a(_0141_),
    .b(_0131_),
    .c(_1390_),
    .y(_0163_)
  );
  al_nand2ft _1993_ (
    .a(_0152_),
    .b(_0163_),
    .y(N2548)
  );
  al_nand2 _1994_ (
    .a(N1),
    .b(N358),
    .y(_0184_)
  );
  al_ao21 _1995_ (
    .a(_1390_),
    .b(_0141_),
    .c(_0131_),
    .y(_0195_)
  );
  al_nand2 _1996_ (
    .a(N341),
    .b(N18),
    .y(_0205_)
  );
  al_ao21ttf _1997_ (
    .a(_1411_),
    .b(_0098_),
    .c(_0087_),
    .y(_0216_)
  );
  al_nand2 _1998_ (
    .a(N324),
    .b(N35),
    .y(_0237_)
  );
  al_ao21ttf _1999_ (
    .a(_1433_),
    .b(_0054_),
    .c(_0044_),
    .y(_0238_)
  );
  al_nand2 _2000_ (
    .a(N307),
    .b(N52),
    .y(_0249_)
  );
  al_and2 _2001_ (
    .a(N273),
    .b(N69),
    .y(_0260_)
  );
  al_and3 _2002_ (
    .a(N290),
    .b(N86),
    .c(_0260_),
    .y(_0271_)
  );
  al_nand2 _2003_ (
    .a(N290),
    .b(N69),
    .y(_0281_)
  );
  al_ao21ttf _2004_ (
    .a(N273),
    .b(N86),
    .c(_0281_),
    .y(_0292_)
  );
  al_oai21ftf _2005_ (
    .a(_0292_),
    .b(_0271_),
    .c(_0011_),
    .y(_0303_)
  );
  al_or3fft _2006_ (
    .a(_0292_),
    .b(_0011_),
    .c(_0271_),
    .y(_0314_)
  );
  al_and3 _2007_ (
    .a(_0249_),
    .b(_0303_),
    .c(_0314_),
    .y(_0325_)
  );
  al_ao21 _2008_ (
    .a(_0303_),
    .b(_0314_),
    .c(_0249_),
    .y(_0335_)
  );
  al_nand3ftt _2009_ (
    .a(_0325_),
    .b(_0238_),
    .c(_0335_),
    .y(_0346_)
  );
  al_ao21ftt _2010_ (
    .a(_0325_),
    .b(_0335_),
    .c(_0238_),
    .y(_0357_)
  );
  al_and3 _2011_ (
    .a(_0237_),
    .b(_0346_),
    .c(_0357_),
    .y(_0368_)
  );
  al_ao21 _2012_ (
    .a(_0346_),
    .b(_0357_),
    .c(_0237_),
    .y(_0379_)
  );
  al_and3ftt _2013_ (
    .a(_0368_),
    .b(_0216_),
    .c(_0379_),
    .y(_0389_)
  );
  al_ao21ftt _2014_ (
    .a(_0368_),
    .b(_0379_),
    .c(_0216_),
    .y(_0400_)
  );
  al_nor3fft _2015_ (
    .a(_0205_),
    .b(_0400_),
    .c(_0389_),
    .y(_0411_)
  );
  al_oai21ftf _2016_ (
    .a(_0400_),
    .b(_0389_),
    .c(_0205_),
    .y(_0422_)
  );
  al_and3ftt _2017_ (
    .a(_0411_),
    .b(_0422_),
    .c(_0195_),
    .y(_0433_)
  );
  al_ao21ftt _2018_ (
    .a(_0411_),
    .b(_0422_),
    .c(_0195_),
    .y(_0443_)
  );
  al_nor3fft _2019_ (
    .a(_0184_),
    .b(_0443_),
    .c(_0433_),
    .y(_0454_)
  );
  al_oai21ftf _2020_ (
    .a(_0443_),
    .b(_0433_),
    .c(_0184_),
    .y(_0465_)
  );
  al_nand2ft _2021_ (
    .a(_0454_),
    .b(_0465_),
    .y(N2877)
  );
  al_nand2 _2022_ (
    .a(N1),
    .b(N375),
    .y(_0485_)
  );
  al_ao21 _2023_ (
    .a(_0184_),
    .b(_0443_),
    .c(_0433_),
    .y(_0496_)
  );
  al_nand2 _2024_ (
    .a(N358),
    .b(N18),
    .y(_0507_)
  );
  al_ao21 _2025_ (
    .a(_0205_),
    .b(_0400_),
    .c(_0389_),
    .y(_0517_)
  );
  al_nand2 _2026_ (
    .a(N341),
    .b(N35),
    .y(_0528_)
  );
  al_ao21ttf _2027_ (
    .a(_0237_),
    .b(_0357_),
    .c(_0346_),
    .y(_0538_)
  );
  al_nand2 _2028_ (
    .a(N324),
    .b(N52),
    .y(_0549_)
  );
  al_ao21ttf _2029_ (
    .a(_0249_),
    .b(_0314_),
    .c(_0303_),
    .y(_0559_)
  );
  al_nand2 _2030_ (
    .a(N307),
    .b(N69),
    .y(_0569_)
  );
  al_and2 _2031_ (
    .a(N273),
    .b(N86),
    .y(_0577_)
  );
  al_and3 _2032_ (
    .a(N290),
    .b(N103),
    .c(_0577_),
    .y(_0578_)
  );
  al_nand2 _2033_ (
    .a(N290),
    .b(N86),
    .y(_0579_)
  );
  al_ao21ttf _2034_ (
    .a(N273),
    .b(N103),
    .c(_0579_),
    .y(_0580_)
  );
  al_oai21ftf _2035_ (
    .a(_0580_),
    .b(_0578_),
    .c(_0271_),
    .y(_0581_)
  );
  al_or3fft _2036_ (
    .a(_0580_),
    .b(_0271_),
    .c(_0578_),
    .y(_0582_)
  );
  al_and3 _2037_ (
    .a(_0569_),
    .b(_0581_),
    .c(_0582_),
    .y(_0583_)
  );
  al_ao21 _2038_ (
    .a(_0581_),
    .b(_0582_),
    .c(_0569_),
    .y(_0584_)
  );
  al_nand3ftt _2039_ (
    .a(_0583_),
    .b(_0559_),
    .c(_0584_),
    .y(_0585_)
  );
  al_ao21ftt _2040_ (
    .a(_0583_),
    .b(_0584_),
    .c(_0559_),
    .y(_0586_)
  );
  al_and3 _2041_ (
    .a(_0549_),
    .b(_0585_),
    .c(_0586_),
    .y(_0587_)
  );
  al_ao21 _2042_ (
    .a(_0585_),
    .b(_0586_),
    .c(_0549_),
    .y(_0588_)
  );
  al_nand3ftt _2043_ (
    .a(_0587_),
    .b(_0538_),
    .c(_0588_),
    .y(_0589_)
  );
  al_ao21ftt _2044_ (
    .a(_0587_),
    .b(_0588_),
    .c(_0538_),
    .y(_0590_)
  );
  al_and3 _2045_ (
    .a(_0528_),
    .b(_0589_),
    .c(_0590_),
    .y(_0591_)
  );
  al_ao21 _2046_ (
    .a(_0589_),
    .b(_0590_),
    .c(_0528_),
    .y(_0592_)
  );
  al_and3ftt _2047_ (
    .a(_0591_),
    .b(_0592_),
    .c(_0517_),
    .y(_0593_)
  );
  al_ao21ftt _2048_ (
    .a(_0591_),
    .b(_0592_),
    .c(_0517_),
    .y(_0594_)
  );
  al_nor3fft _2049_ (
    .a(_0507_),
    .b(_0594_),
    .c(_0593_),
    .y(_0595_)
  );
  al_oai21ftf _2050_ (
    .a(_0594_),
    .b(_0593_),
    .c(_0507_),
    .y(_0596_)
  );
  al_and3ftt _2051_ (
    .a(_0595_),
    .b(_0596_),
    .c(_0496_),
    .y(_0597_)
  );
  al_ao21ftt _2052_ (
    .a(_0595_),
    .b(_0596_),
    .c(_0496_),
    .y(_0598_)
  );
  al_nor3fft _2053_ (
    .a(_0485_),
    .b(_0598_),
    .c(_0597_),
    .y(_0599_)
  );
  al_oai21ftf _2054_ (
    .a(_0598_),
    .b(_0597_),
    .c(_0485_),
    .y(_0600_)
  );
  al_nand2ft _2055_ (
    .a(_0599_),
    .b(_0600_),
    .y(N3211)
  );
  al_nand2 _2056_ (
    .a(N1),
    .b(N392),
    .y(_0601_)
  );
  al_ao21 _2057_ (
    .a(_0485_),
    .b(_0598_),
    .c(_0597_),
    .y(_0602_)
  );
  al_nand2 _2058_ (
    .a(N375),
    .b(N18),
    .y(_0603_)
  );
  al_ao21 _2059_ (
    .a(_0507_),
    .b(_0594_),
    .c(_0593_),
    .y(_0604_)
  );
  al_nand2 _2060_ (
    .a(N358),
    .b(N35),
    .y(_0605_)
  );
  al_ao21ttf _2061_ (
    .a(_0528_),
    .b(_0590_),
    .c(_0589_),
    .y(_0606_)
  );
  al_nand2 _2062_ (
    .a(N341),
    .b(N52),
    .y(_0607_)
  );
  al_ao21ttf _2063_ (
    .a(_0549_),
    .b(_0586_),
    .c(_0585_),
    .y(_0608_)
  );
  al_nand2 _2064_ (
    .a(N324),
    .b(N69),
    .y(_0609_)
  );
  al_ao21ttf _2065_ (
    .a(_0569_),
    .b(_0582_),
    .c(_0581_),
    .y(_0610_)
  );
  al_nand2 _2066_ (
    .a(N307),
    .b(N86),
    .y(_0611_)
  );
  al_and2 _2067_ (
    .a(N273),
    .b(N103),
    .y(_0612_)
  );
  al_and3 _2068_ (
    .a(N290),
    .b(N120),
    .c(_0612_),
    .y(_0613_)
  );
  al_nand2 _2069_ (
    .a(N290),
    .b(N103),
    .y(_0614_)
  );
  al_ao21ttf _2070_ (
    .a(N273),
    .b(N120),
    .c(_0614_),
    .y(_0615_)
  );
  al_oai21ftf _2071_ (
    .a(_0615_),
    .b(_0613_),
    .c(_0578_),
    .y(_0616_)
  );
  al_nand2 _2072_ (
    .a(N273),
    .b(N120),
    .y(_0617_)
  );
  al_nand3ftt _2073_ (
    .a(_0614_),
    .b(_0577_),
    .c(_0617_),
    .y(_0618_)
  );
  al_and3 _2074_ (
    .a(_0611_),
    .b(_0618_),
    .c(_0616_),
    .y(_0619_)
  );
  al_ao21 _2075_ (
    .a(_0618_),
    .b(_0616_),
    .c(_0611_),
    .y(_0620_)
  );
  al_nand3ftt _2076_ (
    .a(_0619_),
    .b(_0620_),
    .c(_0610_),
    .y(_0621_)
  );
  al_ao21ftt _2077_ (
    .a(_0619_),
    .b(_0620_),
    .c(_0610_),
    .y(_0622_)
  );
  al_and3 _2078_ (
    .a(_0609_),
    .b(_0621_),
    .c(_0622_),
    .y(_0623_)
  );
  al_ao21 _2079_ (
    .a(_0621_),
    .b(_0622_),
    .c(_0609_),
    .y(_0624_)
  );
  al_and3ftt _2080_ (
    .a(_0623_),
    .b(_0624_),
    .c(_0608_),
    .y(_0625_)
  );
  al_ao21ftt _2081_ (
    .a(_0623_),
    .b(_0624_),
    .c(_0608_),
    .y(_0626_)
  );
  al_nor3fft _2082_ (
    .a(_0607_),
    .b(_0626_),
    .c(_0625_),
    .y(_0627_)
  );
  al_oai21ftf _2083_ (
    .a(_0626_),
    .b(_0625_),
    .c(_0607_),
    .y(_0628_)
  );
  al_and3ftt _2084_ (
    .a(_0627_),
    .b(_0628_),
    .c(_0606_),
    .y(_0629_)
  );
  al_ao21ftt _2085_ (
    .a(_0627_),
    .b(_0628_),
    .c(_0606_),
    .y(_0630_)
  );
  al_nor3fft _2086_ (
    .a(_0605_),
    .b(_0630_),
    .c(_0629_),
    .y(_0631_)
  );
  al_oai21ftf _2087_ (
    .a(_0630_),
    .b(_0629_),
    .c(_0605_),
    .y(_0632_)
  );
  al_and3ftt _2088_ (
    .a(_0631_),
    .b(_0604_),
    .c(_0632_),
    .y(_0633_)
  );
  al_ao21ftt _2089_ (
    .a(_0631_),
    .b(_0632_),
    .c(_0604_),
    .y(_0634_)
  );
  al_nor3fft _2090_ (
    .a(_0603_),
    .b(_0634_),
    .c(_0633_),
    .y(_0635_)
  );
  al_oai21ftf _2091_ (
    .a(_0634_),
    .b(_0633_),
    .c(_0603_),
    .y(_0636_)
  );
  al_nand3ftt _2092_ (
    .a(_0635_),
    .b(_0602_),
    .c(_0636_),
    .y(_0637_)
  );
  al_ao21ftt _2093_ (
    .a(_0635_),
    .b(_0636_),
    .c(_0602_),
    .y(_0638_)
  );
  al_and3 _2094_ (
    .a(_0601_),
    .b(_0637_),
    .c(_0638_),
    .y(_0639_)
  );
  al_ao21 _2095_ (
    .a(_0637_),
    .b(_0638_),
    .c(_0601_),
    .y(_0640_)
  );
  al_nand2ft _2096_ (
    .a(_0639_),
    .b(_0640_),
    .y(N3552)
  );
  al_nand2 _2097_ (
    .a(N1),
    .b(N409),
    .y(_0641_)
  );
  al_ao21ttf _2098_ (
    .a(_0601_),
    .b(_0638_),
    .c(_0637_),
    .y(_0642_)
  );
  al_nand2 _2099_ (
    .a(N392),
    .b(N18),
    .y(_0643_)
  );
  al_ao21 _2100_ (
    .a(_0603_),
    .b(_0634_),
    .c(_0633_),
    .y(_0644_)
  );
  al_nand2 _2101_ (
    .a(N375),
    .b(N35),
    .y(_0645_)
  );
  al_ao21 _2102_ (
    .a(_0605_),
    .b(_0630_),
    .c(_0629_),
    .y(_0646_)
  );
  al_nand2 _2103_ (
    .a(N358),
    .b(N52),
    .y(_0647_)
  );
  al_ao21 _2104_ (
    .a(_0607_),
    .b(_0626_),
    .c(_0625_),
    .y(_0648_)
  );
  al_nand2 _2105_ (
    .a(N341),
    .b(N69),
    .y(_0649_)
  );
  al_ao21ttf _2106_ (
    .a(_0609_),
    .b(_0622_),
    .c(_0621_),
    .y(_0650_)
  );
  al_nand2 _2107_ (
    .a(N324),
    .b(N86),
    .y(_0651_)
  );
  al_ao21ttf _2108_ (
    .a(_0611_),
    .b(_0618_),
    .c(_0616_),
    .y(_0652_)
  );
  al_nand2 _2109_ (
    .a(N307),
    .b(N103),
    .y(_0653_)
  );
  al_and2 _2110_ (
    .a(N273),
    .b(N137),
    .y(_0654_)
  );
  al_and3 _2111_ (
    .a(N290),
    .b(N120),
    .c(_0654_),
    .y(_0655_)
  );
  al_nand2 _2112_ (
    .a(N290),
    .b(N120),
    .y(_0656_)
  );
  al_ao21ttf _2113_ (
    .a(N273),
    .b(N137),
    .c(_0656_),
    .y(_0657_)
  );
  al_oai21ftf _2114_ (
    .a(_0657_),
    .b(_0655_),
    .c(_0613_),
    .y(_0658_)
  );
  al_nand2 _2115_ (
    .a(N273),
    .b(N137),
    .y(_0659_)
  );
  al_nand3ftt _2116_ (
    .a(_0656_),
    .b(_0612_),
    .c(_0659_),
    .y(_0660_)
  );
  al_nand3 _2117_ (
    .a(_0653_),
    .b(_0660_),
    .c(_0658_),
    .y(_0661_)
  );
  al_ao21 _2118_ (
    .a(_0660_),
    .b(_0658_),
    .c(_0653_),
    .y(_0662_)
  );
  al_nand3 _2119_ (
    .a(_0661_),
    .b(_0652_),
    .c(_0662_),
    .y(_0663_)
  );
  al_ao21 _2120_ (
    .a(_0661_),
    .b(_0662_),
    .c(_0652_),
    .y(_0664_)
  );
  al_and3 _2121_ (
    .a(_0651_),
    .b(_0663_),
    .c(_0664_),
    .y(_0665_)
  );
  al_ao21 _2122_ (
    .a(_0663_),
    .b(_0664_),
    .c(_0651_),
    .y(_0666_)
  );
  al_and3ftt _2123_ (
    .a(_0665_),
    .b(_0650_),
    .c(_0666_),
    .y(_0667_)
  );
  al_ao21ftt _2124_ (
    .a(_0665_),
    .b(_0666_),
    .c(_0650_),
    .y(_0668_)
  );
  al_or3fft _2125_ (
    .a(_0649_),
    .b(_0668_),
    .c(_0667_),
    .y(_0669_)
  );
  al_oai21ftf _2126_ (
    .a(_0668_),
    .b(_0667_),
    .c(_0649_),
    .y(_0670_)
  );
  al_and3 _2127_ (
    .a(_0669_),
    .b(_0648_),
    .c(_0670_),
    .y(_0671_)
  );
  al_ao21 _2128_ (
    .a(_0669_),
    .b(_0670_),
    .c(_0648_),
    .y(_0672_)
  );
  al_nor3fft _2129_ (
    .a(_0647_),
    .b(_0672_),
    .c(_0671_),
    .y(_0673_)
  );
  al_oai21ftf _2130_ (
    .a(_0672_),
    .b(_0671_),
    .c(_0647_),
    .y(_0674_)
  );
  al_and3ftt _2131_ (
    .a(_0673_),
    .b(_0674_),
    .c(_0646_),
    .y(_0675_)
  );
  al_ao21ftt _2132_ (
    .a(_0673_),
    .b(_0674_),
    .c(_0646_),
    .y(_0676_)
  );
  al_nor3fft _2133_ (
    .a(_0645_),
    .b(_0676_),
    .c(_0675_),
    .y(_0677_)
  );
  al_oai21ftf _2134_ (
    .a(_0676_),
    .b(_0675_),
    .c(_0645_),
    .y(_0678_)
  );
  al_and3ftt _2135_ (
    .a(_0677_),
    .b(_0678_),
    .c(_0644_),
    .y(_0679_)
  );
  al_ao21ftt _2136_ (
    .a(_0677_),
    .b(_0678_),
    .c(_0644_),
    .y(_0680_)
  );
  al_nor3fft _2137_ (
    .a(_0643_),
    .b(_0680_),
    .c(_0679_),
    .y(_0681_)
  );
  al_oai21ftf _2138_ (
    .a(_0680_),
    .b(_0679_),
    .c(_0643_),
    .y(_0682_)
  );
  al_and3ftt _2139_ (
    .a(_0681_),
    .b(_0682_),
    .c(_0642_),
    .y(_0683_)
  );
  al_ao21ftt _2140_ (
    .a(_0681_),
    .b(_0682_),
    .c(_0642_),
    .y(_0684_)
  );
  al_nor3fft _2141_ (
    .a(_0641_),
    .b(_0684_),
    .c(_0683_),
    .y(_0685_)
  );
  al_oai21ftf _2142_ (
    .a(_0684_),
    .b(_0683_),
    .c(_0641_),
    .y(_0686_)
  );
  al_nand2ft _2143_ (
    .a(_0685_),
    .b(_0686_),
    .y(N3895)
  );
  al_nand2 _2144_ (
    .a(N1),
    .b(N426),
    .y(_0687_)
  );
  al_ao21 _2145_ (
    .a(_0641_),
    .b(_0684_),
    .c(_0683_),
    .y(_0688_)
  );
  al_nand2 _2146_ (
    .a(N409),
    .b(N18),
    .y(_0689_)
  );
  al_ao21 _2147_ (
    .a(_0643_),
    .b(_0680_),
    .c(_0679_),
    .y(_0690_)
  );
  al_nand2 _2148_ (
    .a(N392),
    .b(N35),
    .y(_0691_)
  );
  al_ao21 _2149_ (
    .a(_0645_),
    .b(_0676_),
    .c(_0675_),
    .y(_0692_)
  );
  al_nand2 _2150_ (
    .a(N375),
    .b(N52),
    .y(_0693_)
  );
  al_ao21 _2151_ (
    .a(_0647_),
    .b(_0672_),
    .c(_0671_),
    .y(_0694_)
  );
  al_nand2 _2152_ (
    .a(N358),
    .b(N69),
    .y(_0695_)
  );
  al_ao21 _2153_ (
    .a(_0649_),
    .b(_0668_),
    .c(_0667_),
    .y(_0696_)
  );
  al_nand2 _2154_ (
    .a(N341),
    .b(N86),
    .y(_0697_)
  );
  al_ao21ttf _2155_ (
    .a(_0651_),
    .b(_0664_),
    .c(_0663_),
    .y(_0698_)
  );
  al_nand2 _2156_ (
    .a(N324),
    .b(N103),
    .y(_0699_)
  );
  al_ao21ttf _2157_ (
    .a(_0653_),
    .b(_0660_),
    .c(_0658_),
    .y(_0700_)
  );
  al_nand2 _2158_ (
    .a(N307),
    .b(N120),
    .y(_0701_)
  );
  al_and3 _2159_ (
    .a(N290),
    .b(N154),
    .c(_0654_),
    .y(_0702_)
  );
  al_nand2 _2160_ (
    .a(N290),
    .b(N137),
    .y(_0703_)
  );
  al_ao21ttf _2161_ (
    .a(N273),
    .b(N154),
    .c(_0703_),
    .y(_0704_)
  );
  al_oai21ftf _2162_ (
    .a(_0704_),
    .b(_0702_),
    .c(_0655_),
    .y(_0705_)
  );
  al_nand2 _2163_ (
    .a(N273),
    .b(N154),
    .y(_0706_)
  );
  al_nand3fft _2164_ (
    .a(_0617_),
    .b(_0703_),
    .c(_0706_),
    .y(_0707_)
  );
  al_nand3 _2165_ (
    .a(_0701_),
    .b(_0707_),
    .c(_0705_),
    .y(_0708_)
  );
  al_ao21 _2166_ (
    .a(_0707_),
    .b(_0705_),
    .c(_0701_),
    .y(_0709_)
  );
  al_nand3 _2167_ (
    .a(_0708_),
    .b(_0700_),
    .c(_0709_),
    .y(_0710_)
  );
  al_ao21 _2168_ (
    .a(_0708_),
    .b(_0709_),
    .c(_0700_),
    .y(_0711_)
  );
  al_and3 _2169_ (
    .a(_0699_),
    .b(_0710_),
    .c(_0711_),
    .y(_0712_)
  );
  al_ao21 _2170_ (
    .a(_0710_),
    .b(_0711_),
    .c(_0699_),
    .y(_0713_)
  );
  al_nand3ftt _2171_ (
    .a(_0712_),
    .b(_0698_),
    .c(_0713_),
    .y(_0714_)
  );
  al_ao21ftt _2172_ (
    .a(_0712_),
    .b(_0713_),
    .c(_0698_),
    .y(_0715_)
  );
  al_and3 _2173_ (
    .a(_0697_),
    .b(_0714_),
    .c(_0715_),
    .y(_0716_)
  );
  al_ao21 _2174_ (
    .a(_0714_),
    .b(_0715_),
    .c(_0697_),
    .y(_0717_)
  );
  al_and3ftt _2175_ (
    .a(_0716_),
    .b(_0717_),
    .c(_0696_),
    .y(_0718_)
  );
  al_ao21ftt _2176_ (
    .a(_0716_),
    .b(_0717_),
    .c(_0696_),
    .y(_0719_)
  );
  al_or3fft _2177_ (
    .a(_0695_),
    .b(_0719_),
    .c(_0718_),
    .y(_0720_)
  );
  al_oai21ftf _2178_ (
    .a(_0719_),
    .b(_0718_),
    .c(_0695_),
    .y(_0721_)
  );
  al_and3 _2179_ (
    .a(_0720_),
    .b(_0694_),
    .c(_0721_),
    .y(_0722_)
  );
  al_ao21 _2180_ (
    .a(_0720_),
    .b(_0721_),
    .c(_0694_),
    .y(_0723_)
  );
  al_nor3fft _2181_ (
    .a(_0693_),
    .b(_0723_),
    .c(_0722_),
    .y(_0724_)
  );
  al_oai21ftf _2182_ (
    .a(_0723_),
    .b(_0722_),
    .c(_0693_),
    .y(_0725_)
  );
  al_and3ftt _2183_ (
    .a(_0724_),
    .b(_0725_),
    .c(_0692_),
    .y(_0726_)
  );
  al_ao21ftt _2184_ (
    .a(_0724_),
    .b(_0725_),
    .c(_0692_),
    .y(_0727_)
  );
  al_nor3fft _2185_ (
    .a(_0691_),
    .b(_0727_),
    .c(_0726_),
    .y(_0728_)
  );
  al_oai21ftf _2186_ (
    .a(_0727_),
    .b(_0726_),
    .c(_0691_),
    .y(_0729_)
  );
  al_and3ftt _2187_ (
    .a(_0728_),
    .b(_0729_),
    .c(_0690_),
    .y(_0730_)
  );
  al_ao21ftt _2188_ (
    .a(_0728_),
    .b(_0729_),
    .c(_0690_),
    .y(_0731_)
  );
  al_nor3fft _2189_ (
    .a(_0689_),
    .b(_0731_),
    .c(_0730_),
    .y(_0732_)
  );
  al_oai21ftf _2190_ (
    .a(_0731_),
    .b(_0730_),
    .c(_0689_),
    .y(_0733_)
  );
  al_and3ftt _2191_ (
    .a(_0732_),
    .b(_0733_),
    .c(_0688_),
    .y(_0734_)
  );
  al_ao21ftt _2192_ (
    .a(_0732_),
    .b(_0733_),
    .c(_0688_),
    .y(_0735_)
  );
  al_nor3fft _2193_ (
    .a(_0687_),
    .b(_0735_),
    .c(_0734_),
    .y(_0736_)
  );
  al_oai21ftf _2194_ (
    .a(_0735_),
    .b(_0734_),
    .c(_0687_),
    .y(_0737_)
  );
  al_nand2ft _2195_ (
    .a(_0736_),
    .b(_0737_),
    .y(N4241)
  );
  al_nand2 _2196_ (
    .a(N1),
    .b(N443),
    .y(_0738_)
  );
  al_ao21 _2197_ (
    .a(_0687_),
    .b(_0735_),
    .c(_0734_),
    .y(_0739_)
  );
  al_nand2 _2198_ (
    .a(N426),
    .b(N18),
    .y(_0740_)
  );
  al_ao21 _2199_ (
    .a(_0689_),
    .b(_0731_),
    .c(_0730_),
    .y(_0741_)
  );
  al_nand2 _2200_ (
    .a(N409),
    .b(N35),
    .y(_0742_)
  );
  al_ao21 _2201_ (
    .a(_0691_),
    .b(_0727_),
    .c(_0726_),
    .y(_0743_)
  );
  al_nand2 _2202_ (
    .a(N392),
    .b(N52),
    .y(_0744_)
  );
  al_ao21 _2203_ (
    .a(_0693_),
    .b(_0723_),
    .c(_0722_),
    .y(_0745_)
  );
  al_nand2 _2204_ (
    .a(N375),
    .b(N69),
    .y(_0746_)
  );
  al_ao21 _2205_ (
    .a(_0695_),
    .b(_0719_),
    .c(_0718_),
    .y(_0747_)
  );
  al_nand2 _2206_ (
    .a(N358),
    .b(N86),
    .y(_0748_)
  );
  al_ao21ttf _2207_ (
    .a(_0697_),
    .b(_0715_),
    .c(_0714_),
    .y(_0749_)
  );
  al_nand2 _2208_ (
    .a(N341),
    .b(N103),
    .y(_0750_)
  );
  al_ao21ttf _2209_ (
    .a(_0699_),
    .b(_0711_),
    .c(_0710_),
    .y(_0751_)
  );
  al_nand2 _2210_ (
    .a(N324),
    .b(N120),
    .y(_0752_)
  );
  al_ao21ttf _2211_ (
    .a(_0701_),
    .b(_0707_),
    .c(_0705_),
    .y(_0753_)
  );
  al_nand2 _2212_ (
    .a(N307),
    .b(N137),
    .y(_0754_)
  );
  al_and2 _2213_ (
    .a(N273),
    .b(N171),
    .y(_0755_)
  );
  al_and3 _2214_ (
    .a(N290),
    .b(N154),
    .c(_0755_),
    .y(_0756_)
  );
  al_nand2 _2215_ (
    .a(N290),
    .b(N154),
    .y(_0757_)
  );
  al_ao21ttf _2216_ (
    .a(N273),
    .b(N171),
    .c(_0757_),
    .y(_0758_)
  );
  al_oai21ftf _2217_ (
    .a(_0758_),
    .b(_0756_),
    .c(_0702_),
    .y(_0759_)
  );
  al_nand2 _2218_ (
    .a(N273),
    .b(N171),
    .y(_0760_)
  );
  al_nand3fft _2219_ (
    .a(_0659_),
    .b(_0757_),
    .c(_0760_),
    .y(_0761_)
  );
  al_nand3 _2220_ (
    .a(_0754_),
    .b(_0761_),
    .c(_0759_),
    .y(_0762_)
  );
  al_ao21 _2221_ (
    .a(_0761_),
    .b(_0759_),
    .c(_0754_),
    .y(_0763_)
  );
  al_nand3 _2222_ (
    .a(_0762_),
    .b(_0753_),
    .c(_0763_),
    .y(_0764_)
  );
  al_ao21 _2223_ (
    .a(_0762_),
    .b(_0763_),
    .c(_0753_),
    .y(_0765_)
  );
  al_and3 _2224_ (
    .a(_0752_),
    .b(_0764_),
    .c(_0765_),
    .y(_0766_)
  );
  al_ao21 _2225_ (
    .a(_0764_),
    .b(_0765_),
    .c(_0752_),
    .y(_0767_)
  );
  al_and3ftt _2226_ (
    .a(_0766_),
    .b(_0751_),
    .c(_0767_),
    .y(_0768_)
  );
  al_ao21ftt _2227_ (
    .a(_0766_),
    .b(_0767_),
    .c(_0751_),
    .y(_0769_)
  );
  al_nor3fft _2228_ (
    .a(_0750_),
    .b(_0769_),
    .c(_0768_),
    .y(_0770_)
  );
  al_oai21ftf _2229_ (
    .a(_0769_),
    .b(_0768_),
    .c(_0750_),
    .y(_0771_)
  );
  al_and3ftt _2230_ (
    .a(_0770_),
    .b(_0771_),
    .c(_0749_),
    .y(_0772_)
  );
  al_ao21ftt _2231_ (
    .a(_0770_),
    .b(_0771_),
    .c(_0749_),
    .y(_0773_)
  );
  al_nor3fft _2232_ (
    .a(_0748_),
    .b(_0773_),
    .c(_0772_),
    .y(_0774_)
  );
  al_oai21ftf _2233_ (
    .a(_0773_),
    .b(_0772_),
    .c(_0748_),
    .y(_0775_)
  );
  al_nor3fft _2234_ (
    .a(_0747_),
    .b(_0775_),
    .c(_0774_),
    .y(_0776_)
  );
  al_ao21ftt _2235_ (
    .a(_0774_),
    .b(_0775_),
    .c(_0747_),
    .y(_0777_)
  );
  al_or3fft _2236_ (
    .a(_0746_),
    .b(_0777_),
    .c(_0776_),
    .y(_0778_)
  );
  al_oai21ftf _2237_ (
    .a(_0777_),
    .b(_0776_),
    .c(_0746_),
    .y(_0779_)
  );
  al_and3 _2238_ (
    .a(_0745_),
    .b(_0778_),
    .c(_0779_),
    .y(_0780_)
  );
  al_ao21 _2239_ (
    .a(_0778_),
    .b(_0779_),
    .c(_0745_),
    .y(_0781_)
  );
  al_nor3fft _2240_ (
    .a(_0744_),
    .b(_0781_),
    .c(_0780_),
    .y(_0782_)
  );
  al_oai21ftf _2241_ (
    .a(_0781_),
    .b(_0780_),
    .c(_0744_),
    .y(_0783_)
  );
  al_nor3fft _2242_ (
    .a(_0743_),
    .b(_0783_),
    .c(_0782_),
    .y(_0784_)
  );
  al_ao21ftt _2243_ (
    .a(_0782_),
    .b(_0783_),
    .c(_0743_),
    .y(_0785_)
  );
  al_nor3fft _2244_ (
    .a(_0742_),
    .b(_0785_),
    .c(_0784_),
    .y(_0786_)
  );
  al_oai21ftf _2245_ (
    .a(_0785_),
    .b(_0784_),
    .c(_0742_),
    .y(_0787_)
  );
  al_nor3fft _2246_ (
    .a(_0741_),
    .b(_0787_),
    .c(_0786_),
    .y(_0788_)
  );
  al_ao21ftt _2247_ (
    .a(_0786_),
    .b(_0787_),
    .c(_0741_),
    .y(_0789_)
  );
  al_nor3fft _2248_ (
    .a(_0740_),
    .b(_0789_),
    .c(_0788_),
    .y(_0790_)
  );
  al_oai21ftf _2249_ (
    .a(_0789_),
    .b(_0788_),
    .c(_0740_),
    .y(_0791_)
  );
  al_nor3fft _2250_ (
    .a(_0739_),
    .b(_0791_),
    .c(_0790_),
    .y(_0792_)
  );
  al_ao21ftt _2251_ (
    .a(_0790_),
    .b(_0791_),
    .c(_0739_),
    .y(_0793_)
  );
  al_nor3fft _2252_ (
    .a(_0738_),
    .b(_0793_),
    .c(_0792_),
    .y(_0794_)
  );
  al_oai21ftf _2253_ (
    .a(_0793_),
    .b(_0792_),
    .c(_0738_),
    .y(_0795_)
  );
  al_nand2ft _2254_ (
    .a(_0794_),
    .b(_0795_),
    .y(N4591)
  );
  al_nand2 _2255_ (
    .a(N1),
    .b(N460),
    .y(_0796_)
  );
  al_ao21 _2256_ (
    .a(_0738_),
    .b(_0793_),
    .c(_0792_),
    .y(_0797_)
  );
  al_nand2 _2257_ (
    .a(N443),
    .b(N18),
    .y(_0798_)
  );
  al_ao21 _2258_ (
    .a(_0740_),
    .b(_0789_),
    .c(_0788_),
    .y(_0799_)
  );
  al_nand2 _2259_ (
    .a(N426),
    .b(N35),
    .y(_0800_)
  );
  al_ao21 _2260_ (
    .a(_0742_),
    .b(_0785_),
    .c(_0784_),
    .y(_0801_)
  );
  al_nand2 _2261_ (
    .a(N409),
    .b(N52),
    .y(_0802_)
  );
  al_ao21 _2262_ (
    .a(_0744_),
    .b(_0781_),
    .c(_0780_),
    .y(_0803_)
  );
  al_nand2 _2263_ (
    .a(N392),
    .b(N69),
    .y(_0804_)
  );
  al_ao21 _2264_ (
    .a(_0746_),
    .b(_0777_),
    .c(_0776_),
    .y(_0805_)
  );
  al_nand2 _2265_ (
    .a(N375),
    .b(N86),
    .y(_0806_)
  );
  al_ao21 _2266_ (
    .a(_0748_),
    .b(_0773_),
    .c(_0772_),
    .y(_0807_)
  );
  al_nand2 _2267_ (
    .a(N358),
    .b(N103),
    .y(_0808_)
  );
  al_ao21 _2268_ (
    .a(_0750_),
    .b(_0769_),
    .c(_0768_),
    .y(_0809_)
  );
  al_nand2 _2269_ (
    .a(N341),
    .b(N120),
    .y(_0810_)
  );
  al_ao21ttf _2270_ (
    .a(_0752_),
    .b(_0765_),
    .c(_0764_),
    .y(_0811_)
  );
  al_nand2 _2271_ (
    .a(N324),
    .b(N137),
    .y(_0812_)
  );
  al_ao21ttf _2272_ (
    .a(_0754_),
    .b(_0761_),
    .c(_0759_),
    .y(_0813_)
  );
  al_nand2 _2273_ (
    .a(N307),
    .b(N154),
    .y(_0814_)
  );
  al_and3 _2274_ (
    .a(N290),
    .b(N188),
    .c(_0755_),
    .y(_0815_)
  );
  al_nand2 _2275_ (
    .a(N290),
    .b(N171),
    .y(_0816_)
  );
  al_ao21ttf _2276_ (
    .a(N273),
    .b(N188),
    .c(_0816_),
    .y(_0817_)
  );
  al_oai21ftf _2277_ (
    .a(_0817_),
    .b(_0815_),
    .c(_0756_),
    .y(_0818_)
  );
  al_nand2 _2278_ (
    .a(N273),
    .b(N188),
    .y(_0819_)
  );
  al_nand3fft _2279_ (
    .a(_0706_),
    .b(_0816_),
    .c(_0819_),
    .y(_0820_)
  );
  al_nand3 _2280_ (
    .a(_0814_),
    .b(_0820_),
    .c(_0818_),
    .y(_0821_)
  );
  al_ao21 _2281_ (
    .a(_0820_),
    .b(_0818_),
    .c(_0814_),
    .y(_0822_)
  );
  al_nand3 _2282_ (
    .a(_0821_),
    .b(_0813_),
    .c(_0822_),
    .y(_0823_)
  );
  al_ao21 _2283_ (
    .a(_0821_),
    .b(_0822_),
    .c(_0813_),
    .y(_0824_)
  );
  al_and3 _2284_ (
    .a(_0812_),
    .b(_0823_),
    .c(_0824_),
    .y(_0825_)
  );
  al_ao21 _2285_ (
    .a(_0823_),
    .b(_0824_),
    .c(_0812_),
    .y(_0826_)
  );
  al_and3ftt _2286_ (
    .a(_0825_),
    .b(_0826_),
    .c(_0811_),
    .y(_0827_)
  );
  al_ao21ftt _2287_ (
    .a(_0825_),
    .b(_0826_),
    .c(_0811_),
    .y(_0828_)
  );
  al_nor3fft _2288_ (
    .a(_0810_),
    .b(_0828_),
    .c(_0827_),
    .y(_0829_)
  );
  al_oai21ftf _2289_ (
    .a(_0828_),
    .b(_0827_),
    .c(_0810_),
    .y(_0830_)
  );
  al_and3ftt _2290_ (
    .a(_0829_),
    .b(_0809_),
    .c(_0830_),
    .y(_0831_)
  );
  al_ao21ftt _2291_ (
    .a(_0829_),
    .b(_0830_),
    .c(_0809_),
    .y(_0832_)
  );
  al_nor3fft _2292_ (
    .a(_0808_),
    .b(_0832_),
    .c(_0831_),
    .y(_0833_)
  );
  al_oai21ftf _2293_ (
    .a(_0832_),
    .b(_0831_),
    .c(_0808_),
    .y(_0834_)
  );
  al_and3ftt _2294_ (
    .a(_0833_),
    .b(_0834_),
    .c(_0807_),
    .y(_0835_)
  );
  al_ao21ftt _2295_ (
    .a(_0833_),
    .b(_0834_),
    .c(_0807_),
    .y(_0836_)
  );
  al_nor3fft _2296_ (
    .a(_0806_),
    .b(_0836_),
    .c(_0835_),
    .y(_0837_)
  );
  al_oai21ftf _2297_ (
    .a(_0836_),
    .b(_0835_),
    .c(_0806_),
    .y(_0838_)
  );
  al_and3ftt _2298_ (
    .a(_0837_),
    .b(_0838_),
    .c(_0805_),
    .y(_0839_)
  );
  al_ao21ftt _2299_ (
    .a(_0837_),
    .b(_0838_),
    .c(_0805_),
    .y(_0840_)
  );
  al_or3fft _2300_ (
    .a(_0804_),
    .b(_0840_),
    .c(_0839_),
    .y(_0841_)
  );
  al_oai21ftf _2301_ (
    .a(_0840_),
    .b(_0839_),
    .c(_0804_),
    .y(_0842_)
  );
  al_and3 _2302_ (
    .a(_0803_),
    .b(_0841_),
    .c(_0842_),
    .y(_0843_)
  );
  al_ao21 _2303_ (
    .a(_0841_),
    .b(_0842_),
    .c(_0803_),
    .y(_0844_)
  );
  al_nor3fft _2304_ (
    .a(_0802_),
    .b(_0844_),
    .c(_0843_),
    .y(_0845_)
  );
  al_oai21ftf _2305_ (
    .a(_0844_),
    .b(_0843_),
    .c(_0802_),
    .y(_0846_)
  );
  al_and3ftt _2306_ (
    .a(_0845_),
    .b(_0846_),
    .c(_0801_),
    .y(_0847_)
  );
  al_ao21ftt _2307_ (
    .a(_0845_),
    .b(_0846_),
    .c(_0801_),
    .y(_0848_)
  );
  al_or3fft _2308_ (
    .a(_0800_),
    .b(_0848_),
    .c(_0847_),
    .y(_0849_)
  );
  al_oai21ftf _2309_ (
    .a(_0848_),
    .b(_0847_),
    .c(_0800_),
    .y(_0850_)
  );
  al_and3 _2310_ (
    .a(_0849_),
    .b(_0799_),
    .c(_0850_),
    .y(_0851_)
  );
  al_ao21 _2311_ (
    .a(_0849_),
    .b(_0850_),
    .c(_0799_),
    .y(_0852_)
  );
  al_nor3fft _2312_ (
    .a(_0798_),
    .b(_0852_),
    .c(_0851_),
    .y(_0853_)
  );
  al_oai21ftf _2313_ (
    .a(_0852_),
    .b(_0851_),
    .c(_0798_),
    .y(_0854_)
  );
  al_and3ftt _2314_ (
    .a(_0853_),
    .b(_0854_),
    .c(_0797_),
    .y(_0855_)
  );
  al_ao21ftt _2315_ (
    .a(_0853_),
    .b(_0854_),
    .c(_0797_),
    .y(_0856_)
  );
  al_nor3fft _2316_ (
    .a(_0796_),
    .b(_0856_),
    .c(_0855_),
    .y(_0857_)
  );
  al_oai21ftf _2317_ (
    .a(_0856_),
    .b(_0855_),
    .c(_0796_),
    .y(_0858_)
  );
  al_nand2ft _2318_ (
    .a(_0857_),
    .b(_0858_),
    .y(N4946)
  );
  al_nand2 _2319_ (
    .a(N1),
    .b(N477),
    .y(_0859_)
  );
  al_ao21 _2320_ (
    .a(_0796_),
    .b(_0856_),
    .c(_0855_),
    .y(_0860_)
  );
  al_nand2 _2321_ (
    .a(N460),
    .b(N18),
    .y(_0861_)
  );
  al_ao21 _2322_ (
    .a(_0798_),
    .b(_0852_),
    .c(_0851_),
    .y(_0862_)
  );
  al_nand2 _2323_ (
    .a(N443),
    .b(N35),
    .y(_0863_)
  );
  al_ao21 _2324_ (
    .a(_0800_),
    .b(_0848_),
    .c(_0847_),
    .y(_0864_)
  );
  al_nand2 _2325_ (
    .a(N426),
    .b(N52),
    .y(_0865_)
  );
  al_ao21 _2326_ (
    .a(_0802_),
    .b(_0844_),
    .c(_0843_),
    .y(_0866_)
  );
  al_nand2 _2327_ (
    .a(N409),
    .b(N69),
    .y(_0867_)
  );
  al_ao21 _2328_ (
    .a(_0804_),
    .b(_0840_),
    .c(_0839_),
    .y(_0868_)
  );
  al_nand2 _2329_ (
    .a(N392),
    .b(N86),
    .y(_0869_)
  );
  al_ao21 _2330_ (
    .a(_0806_),
    .b(_0836_),
    .c(_0835_),
    .y(_0870_)
  );
  al_nand2 _2331_ (
    .a(N375),
    .b(N103),
    .y(_0871_)
  );
  al_ao21 _2332_ (
    .a(_0808_),
    .b(_0832_),
    .c(_0831_),
    .y(_0872_)
  );
  al_nand2 _2333_ (
    .a(N358),
    .b(N120),
    .y(_0873_)
  );
  al_ao21 _2334_ (
    .a(_0810_),
    .b(_0828_),
    .c(_0827_),
    .y(_0874_)
  );
  al_nand2 _2335_ (
    .a(N341),
    .b(N137),
    .y(_0875_)
  );
  al_ao21ttf _2336_ (
    .a(_0812_),
    .b(_0824_),
    .c(_0823_),
    .y(_0876_)
  );
  al_nand2 _2337_ (
    .a(N324),
    .b(N154),
    .y(_0877_)
  );
  al_ao21ttf _2338_ (
    .a(_0814_),
    .b(_0820_),
    .c(_0818_),
    .y(_0878_)
  );
  al_nand2 _2339_ (
    .a(N307),
    .b(N171),
    .y(_0879_)
  );
  al_and2 _2340_ (
    .a(N273),
    .b(N205),
    .y(_0880_)
  );
  al_and3 _2341_ (
    .a(N290),
    .b(N188),
    .c(_0880_),
    .y(_0881_)
  );
  al_nand2 _2342_ (
    .a(N290),
    .b(N188),
    .y(_0882_)
  );
  al_ao21ttf _2343_ (
    .a(N273),
    .b(N205),
    .c(_0882_),
    .y(_0883_)
  );
  al_oai21ftf _2344_ (
    .a(_0883_),
    .b(_0881_),
    .c(_0815_),
    .y(_0884_)
  );
  al_nand2 _2345_ (
    .a(N273),
    .b(N205),
    .y(_0885_)
  );
  al_nand3fft _2346_ (
    .a(_0760_),
    .b(_0882_),
    .c(_0885_),
    .y(_0886_)
  );
  al_nand3 _2347_ (
    .a(_0879_),
    .b(_0886_),
    .c(_0884_),
    .y(_0887_)
  );
  al_ao21 _2348_ (
    .a(_0886_),
    .b(_0884_),
    .c(_0879_),
    .y(_0888_)
  );
  al_nand3 _2349_ (
    .a(_0887_),
    .b(_0878_),
    .c(_0888_),
    .y(_0889_)
  );
  al_ao21 _2350_ (
    .a(_0887_),
    .b(_0888_),
    .c(_0878_),
    .y(_0890_)
  );
  al_and3 _2351_ (
    .a(_0877_),
    .b(_0889_),
    .c(_0890_),
    .y(_0891_)
  );
  al_ao21 _2352_ (
    .a(_0889_),
    .b(_0890_),
    .c(_0877_),
    .y(_0892_)
  );
  al_and3ftt _2353_ (
    .a(_0891_),
    .b(_0892_),
    .c(_0876_),
    .y(_0893_)
  );
  al_ao21ftt _2354_ (
    .a(_0891_),
    .b(_0892_),
    .c(_0876_),
    .y(_0894_)
  );
  al_nor3fft _2355_ (
    .a(_0875_),
    .b(_0894_),
    .c(_0893_),
    .y(_0895_)
  );
  al_oai21ftf _2356_ (
    .a(_0894_),
    .b(_0893_),
    .c(_0875_),
    .y(_0896_)
  );
  al_and3ftt _2357_ (
    .a(_0895_),
    .b(_0874_),
    .c(_0896_),
    .y(_0897_)
  );
  al_ao21ftt _2358_ (
    .a(_0895_),
    .b(_0896_),
    .c(_0874_),
    .y(_0898_)
  );
  al_nor3fft _2359_ (
    .a(_0873_),
    .b(_0898_),
    .c(_0897_),
    .y(_0899_)
  );
  al_oai21ftf _2360_ (
    .a(_0898_),
    .b(_0897_),
    .c(_0873_),
    .y(_0900_)
  );
  al_and3ftt _2361_ (
    .a(_0899_),
    .b(_0872_),
    .c(_0900_),
    .y(_0901_)
  );
  al_ao21ftt _2362_ (
    .a(_0899_),
    .b(_0900_),
    .c(_0872_),
    .y(_0902_)
  );
  al_nor3fft _2363_ (
    .a(_0871_),
    .b(_0902_),
    .c(_0901_),
    .y(_0903_)
  );
  al_oai21ftf _2364_ (
    .a(_0902_),
    .b(_0901_),
    .c(_0871_),
    .y(_0904_)
  );
  al_nand3ftt _2365_ (
    .a(_0903_),
    .b(_0870_),
    .c(_0904_),
    .y(_0905_)
  );
  al_ao21ftt _2366_ (
    .a(_0903_),
    .b(_0904_),
    .c(_0870_),
    .y(_0906_)
  );
  al_nand3 _2367_ (
    .a(_0869_),
    .b(_0905_),
    .c(_0906_),
    .y(_0907_)
  );
  al_ao21 _2368_ (
    .a(_0905_),
    .b(_0906_),
    .c(_0869_),
    .y(_0908_)
  );
  al_and3 _2369_ (
    .a(_0907_),
    .b(_0868_),
    .c(_0908_),
    .y(_0909_)
  );
  al_ao21 _2370_ (
    .a(_0907_),
    .b(_0908_),
    .c(_0868_),
    .y(_0910_)
  );
  al_or3fft _2371_ (
    .a(_0867_),
    .b(_0910_),
    .c(_0909_),
    .y(_0911_)
  );
  al_oai21ftf _2372_ (
    .a(_0910_),
    .b(_0909_),
    .c(_0867_),
    .y(_0912_)
  );
  al_and3 _2373_ (
    .a(_0911_),
    .b(_0866_),
    .c(_0912_),
    .y(_0913_)
  );
  al_ao21 _2374_ (
    .a(_0911_),
    .b(_0912_),
    .c(_0866_),
    .y(_0914_)
  );
  al_or3fft _2375_ (
    .a(_0865_),
    .b(_0914_),
    .c(_0913_),
    .y(_0915_)
  );
  al_oai21ftf _2376_ (
    .a(_0914_),
    .b(_0913_),
    .c(_0865_),
    .y(_0916_)
  );
  al_and3 _2377_ (
    .a(_0915_),
    .b(_0864_),
    .c(_0916_),
    .y(_0917_)
  );
  al_ao21 _2378_ (
    .a(_0915_),
    .b(_0916_),
    .c(_0864_),
    .y(_0918_)
  );
  al_or3fft _2379_ (
    .a(_0863_),
    .b(_0918_),
    .c(_0917_),
    .y(_0919_)
  );
  al_oai21ftf _2380_ (
    .a(_0918_),
    .b(_0917_),
    .c(_0863_),
    .y(_0920_)
  );
  al_and3 _2381_ (
    .a(_0919_),
    .b(_0862_),
    .c(_0920_),
    .y(_0921_)
  );
  al_ao21 _2382_ (
    .a(_0919_),
    .b(_0920_),
    .c(_0862_),
    .y(_0922_)
  );
  al_nor3fft _2383_ (
    .a(_0861_),
    .b(_0922_),
    .c(_0921_),
    .y(_0923_)
  );
  al_oai21ftf _2384_ (
    .a(_0922_),
    .b(_0921_),
    .c(_0861_),
    .y(_0924_)
  );
  al_and3ftt _2385_ (
    .a(_0923_),
    .b(_0924_),
    .c(_0860_),
    .y(_0925_)
  );
  al_ao21ftt _2386_ (
    .a(_0923_),
    .b(_0924_),
    .c(_0860_),
    .y(_0926_)
  );
  al_nor3fft _2387_ (
    .a(_0859_),
    .b(_0926_),
    .c(_0925_),
    .y(_0927_)
  );
  al_oai21ftf _2388_ (
    .a(_0926_),
    .b(_0925_),
    .c(_0859_),
    .y(_0928_)
  );
  al_nand2ft _2389_ (
    .a(_0927_),
    .b(_0928_),
    .y(N5308)
  );
  al_nand2 _2390_ (
    .a(N1),
    .b(N494),
    .y(_0929_)
  );
  al_ao21 _2391_ (
    .a(_0859_),
    .b(_0926_),
    .c(_0925_),
    .y(_0930_)
  );
  al_nand2 _2392_ (
    .a(N477),
    .b(N18),
    .y(_0931_)
  );
  al_ao21 _2393_ (
    .a(_0861_),
    .b(_0922_),
    .c(_0921_),
    .y(_0932_)
  );
  al_nand2 _2394_ (
    .a(N460),
    .b(N35),
    .y(_0933_)
  );
  al_ao21 _2395_ (
    .a(_0863_),
    .b(_0918_),
    .c(_0917_),
    .y(_0934_)
  );
  al_nand2 _2396_ (
    .a(N443),
    .b(N52),
    .y(_0935_)
  );
  al_ao21 _2397_ (
    .a(_0865_),
    .b(_0914_),
    .c(_0913_),
    .y(_0936_)
  );
  al_nand2 _2398_ (
    .a(N426),
    .b(N69),
    .y(_0937_)
  );
  al_ao21 _2399_ (
    .a(_0867_),
    .b(_0910_),
    .c(_0909_),
    .y(_0938_)
  );
  al_nand2 _2400_ (
    .a(N409),
    .b(N86),
    .y(_0939_)
  );
  al_ao21ttf _2401_ (
    .a(_0869_),
    .b(_0906_),
    .c(_0905_),
    .y(_0940_)
  );
  al_nand2 _2402_ (
    .a(N392),
    .b(N103),
    .y(_0941_)
  );
  al_ao21 _2403_ (
    .a(_0871_),
    .b(_0902_),
    .c(_0901_),
    .y(_0942_)
  );
  al_nand2 _2404_ (
    .a(N375),
    .b(N120),
    .y(_0943_)
  );
  al_ao21 _2405_ (
    .a(_0873_),
    .b(_0898_),
    .c(_0897_),
    .y(_0944_)
  );
  al_nand2 _2406_ (
    .a(N358),
    .b(N137),
    .y(_0945_)
  );
  al_ao21 _2407_ (
    .a(_0875_),
    .b(_0894_),
    .c(_0893_),
    .y(_0946_)
  );
  al_nand2 _2408_ (
    .a(N341),
    .b(N154),
    .y(_0947_)
  );
  al_ao21ttf _2409_ (
    .a(_0877_),
    .b(_0890_),
    .c(_0889_),
    .y(_0948_)
  );
  al_nand2 _2410_ (
    .a(N324),
    .b(N171),
    .y(_0949_)
  );
  al_ao21ttf _2411_ (
    .a(_0879_),
    .b(_0886_),
    .c(_0884_),
    .y(_0950_)
  );
  al_nand2 _2412_ (
    .a(N307),
    .b(N188),
    .y(_0951_)
  );
  al_and3 _2413_ (
    .a(N290),
    .b(N222),
    .c(_0880_),
    .y(_0952_)
  );
  al_nand2 _2414_ (
    .a(N290),
    .b(N205),
    .y(_0953_)
  );
  al_ao21ttf _2415_ (
    .a(N273),
    .b(N222),
    .c(_0953_),
    .y(_0954_)
  );
  al_oai21ftf _2416_ (
    .a(_0954_),
    .b(_0952_),
    .c(_0881_),
    .y(_0955_)
  );
  al_nand2 _2417_ (
    .a(N273),
    .b(N222),
    .y(_0956_)
  );
  al_nand3fft _2418_ (
    .a(_0819_),
    .b(_0953_),
    .c(_0956_),
    .y(_0957_)
  );
  al_nand3 _2419_ (
    .a(_0951_),
    .b(_0957_),
    .c(_0955_),
    .y(_0958_)
  );
  al_ao21 _2420_ (
    .a(_0957_),
    .b(_0955_),
    .c(_0951_),
    .y(_0959_)
  );
  al_nand3 _2421_ (
    .a(_0958_),
    .b(_0950_),
    .c(_0959_),
    .y(_0960_)
  );
  al_ao21 _2422_ (
    .a(_0958_),
    .b(_0959_),
    .c(_0950_),
    .y(_0961_)
  );
  al_and3 _2423_ (
    .a(_0949_),
    .b(_0960_),
    .c(_0961_),
    .y(_0962_)
  );
  al_ao21 _2424_ (
    .a(_0960_),
    .b(_0961_),
    .c(_0949_),
    .y(_0963_)
  );
  al_and3ftt _2425_ (
    .a(_0962_),
    .b(_0948_),
    .c(_0963_),
    .y(_0964_)
  );
  al_ao21ftt _2426_ (
    .a(_0962_),
    .b(_0963_),
    .c(_0948_),
    .y(_0965_)
  );
  al_nor3fft _2427_ (
    .a(_0947_),
    .b(_0965_),
    .c(_0964_),
    .y(_0966_)
  );
  al_oai21ftf _2428_ (
    .a(_0965_),
    .b(_0964_),
    .c(_0947_),
    .y(_0967_)
  );
  al_and3ftt _2429_ (
    .a(_0966_),
    .b(_0946_),
    .c(_0967_),
    .y(_0968_)
  );
  al_ao21ftt _2430_ (
    .a(_0966_),
    .b(_0967_),
    .c(_0946_),
    .y(_0969_)
  );
  al_nor3fft _2431_ (
    .a(_0945_),
    .b(_0969_),
    .c(_0968_),
    .y(_0970_)
  );
  al_oai21ftf _2432_ (
    .a(_0969_),
    .b(_0968_),
    .c(_0945_),
    .y(_0971_)
  );
  al_nand3ftt _2433_ (
    .a(_0970_),
    .b(_0944_),
    .c(_0971_),
    .y(_0972_)
  );
  al_ao21ftt _2434_ (
    .a(_0970_),
    .b(_0971_),
    .c(_0944_),
    .y(_0973_)
  );
  al_nand3 _2435_ (
    .a(_0943_),
    .b(_0972_),
    .c(_0973_),
    .y(_0974_)
  );
  al_ao21 _2436_ (
    .a(_0972_),
    .b(_0973_),
    .c(_0943_),
    .y(_0975_)
  );
  al_and3 _2437_ (
    .a(_0974_),
    .b(_0942_),
    .c(_0975_),
    .y(_0976_)
  );
  al_ao21 _2438_ (
    .a(_0974_),
    .b(_0975_),
    .c(_0942_),
    .y(_0977_)
  );
  al_or3fft _2439_ (
    .a(_0941_),
    .b(_0977_),
    .c(_0976_),
    .y(_0978_)
  );
  al_oai21ftf _2440_ (
    .a(_0977_),
    .b(_0976_),
    .c(_0941_),
    .y(_0979_)
  );
  al_and3 _2441_ (
    .a(_0978_),
    .b(_0940_),
    .c(_0979_),
    .y(_0980_)
  );
  al_ao21 _2442_ (
    .a(_0978_),
    .b(_0979_),
    .c(_0940_),
    .y(_0981_)
  );
  al_nor3fft _2443_ (
    .a(_0939_),
    .b(_0981_),
    .c(_0980_),
    .y(_0982_)
  );
  al_oai21ftf _2444_ (
    .a(_0981_),
    .b(_0980_),
    .c(_0939_),
    .y(_0983_)
  );
  al_nand3ftt _2445_ (
    .a(_0982_),
    .b(_0983_),
    .c(_0938_),
    .y(_0984_)
  );
  al_ao21ftt _2446_ (
    .a(_0982_),
    .b(_0983_),
    .c(_0938_),
    .y(_0985_)
  );
  al_nand3 _2447_ (
    .a(_0937_),
    .b(_0984_),
    .c(_0985_),
    .y(_0986_)
  );
  al_ao21 _2448_ (
    .a(_0984_),
    .b(_0985_),
    .c(_0937_),
    .y(_0987_)
  );
  al_and3 _2449_ (
    .a(_0986_),
    .b(_0936_),
    .c(_0987_),
    .y(_0988_)
  );
  al_ao21 _2450_ (
    .a(_0986_),
    .b(_0987_),
    .c(_0936_),
    .y(_0989_)
  );
  al_nor3fft _2451_ (
    .a(_0935_),
    .b(_0989_),
    .c(_0988_),
    .y(_0990_)
  );
  al_oai21ftf _2452_ (
    .a(_0989_),
    .b(_0988_),
    .c(_0935_),
    .y(_0991_)
  );
  al_nand3ftt _2453_ (
    .a(_0990_),
    .b(_0991_),
    .c(_0934_),
    .y(_0992_)
  );
  al_ao21ftt _2454_ (
    .a(_0990_),
    .b(_0991_),
    .c(_0934_),
    .y(_0993_)
  );
  al_nand3 _2455_ (
    .a(_0933_),
    .b(_0992_),
    .c(_0993_),
    .y(_0994_)
  );
  al_ao21 _2456_ (
    .a(_0992_),
    .b(_0993_),
    .c(_0933_),
    .y(_0995_)
  );
  al_and3 _2457_ (
    .a(_0994_),
    .b(_0932_),
    .c(_0995_),
    .y(_0996_)
  );
  al_ao21 _2458_ (
    .a(_0994_),
    .b(_0995_),
    .c(_0932_),
    .y(_0997_)
  );
  al_nor3fft _2459_ (
    .a(_0931_),
    .b(_0997_),
    .c(_0996_),
    .y(_0998_)
  );
  al_oai21ftf _2460_ (
    .a(_0997_),
    .b(_0996_),
    .c(_0931_),
    .y(_0999_)
  );
  al_and3ftt _2461_ (
    .a(_0998_),
    .b(_0999_),
    .c(_0930_),
    .y(_1000_)
  );
  al_ao21ftt _2462_ (
    .a(_0998_),
    .b(_0999_),
    .c(_0930_),
    .y(_1001_)
  );
  al_nor3fft _2463_ (
    .a(_0929_),
    .b(_1001_),
    .c(_1000_),
    .y(_1002_)
  );
  al_oai21ftf _2464_ (
    .a(_1001_),
    .b(_1000_),
    .c(_0929_),
    .y(_1003_)
  );
  al_nand2ft _2465_ (
    .a(_1002_),
    .b(_1003_),
    .y(N5672)
  );
  al_nand2 _2466_ (
    .a(N1),
    .b(N511),
    .y(_1004_)
  );
  al_ao21 _2467_ (
    .a(_0929_),
    .b(_1001_),
    .c(_1000_),
    .y(_1005_)
  );
  al_nand2 _2468_ (
    .a(N494),
    .b(N18),
    .y(_1006_)
  );
  al_ao21 _2469_ (
    .a(_0931_),
    .b(_0997_),
    .c(_0996_),
    .y(_1007_)
  );
  al_nand2 _2470_ (
    .a(N477),
    .b(N35),
    .y(_1008_)
  );
  al_ao21ttf _2471_ (
    .a(_0933_),
    .b(_0993_),
    .c(_0992_),
    .y(_1009_)
  );
  al_nand2 _2472_ (
    .a(N460),
    .b(N52),
    .y(_1010_)
  );
  al_ao21 _2473_ (
    .a(_0935_),
    .b(_0989_),
    .c(_0988_),
    .y(_1011_)
  );
  al_nand2 _2474_ (
    .a(N443),
    .b(N69),
    .y(_1012_)
  );
  al_ao21ttf _2475_ (
    .a(_0937_),
    .b(_0985_),
    .c(_0984_),
    .y(_1013_)
  );
  al_nand2 _2476_ (
    .a(N426),
    .b(N86),
    .y(_1014_)
  );
  al_ao21 _2477_ (
    .a(_0939_),
    .b(_0981_),
    .c(_0980_),
    .y(_1015_)
  );
  al_nand2 _2478_ (
    .a(N409),
    .b(N103),
    .y(_1016_)
  );
  al_ao21 _2479_ (
    .a(_0941_),
    .b(_0977_),
    .c(_0976_),
    .y(_1017_)
  );
  al_nand2 _2480_ (
    .a(N392),
    .b(N120),
    .y(_1018_)
  );
  al_ao21ttf _2481_ (
    .a(_0943_),
    .b(_0973_),
    .c(_0972_),
    .y(_1019_)
  );
  al_nand2 _2482_ (
    .a(N375),
    .b(N137),
    .y(_1020_)
  );
  al_ao21 _2483_ (
    .a(_0945_),
    .b(_0969_),
    .c(_0968_),
    .y(_1021_)
  );
  al_nand2 _2484_ (
    .a(N358),
    .b(N154),
    .y(_1022_)
  );
  al_ao21 _2485_ (
    .a(_0947_),
    .b(_0965_),
    .c(_0964_),
    .y(_1023_)
  );
  al_nand2 _2486_ (
    .a(N341),
    .b(N171),
    .y(_1024_)
  );
  al_ao21ttf _2487_ (
    .a(_0949_),
    .b(_0961_),
    .c(_0960_),
    .y(_1025_)
  );
  al_nand2 _2488_ (
    .a(N324),
    .b(N188),
    .y(_1026_)
  );
  al_aoi21ttf _2489_ (
    .a(_0951_),
    .b(_0957_),
    .c(_0955_),
    .y(_1027_)
  );
  al_nand2 _2490_ (
    .a(N307),
    .b(N205),
    .y(_1028_)
  );
  al_and2 _2491_ (
    .a(N290),
    .b(N239),
    .y(_1029_)
  );
  al_nand3 _2492_ (
    .a(N273),
    .b(N222),
    .c(_1029_),
    .y(_1030_)
  );
  al_nand2 _2493_ (
    .a(N290),
    .b(N222),
    .y(_1031_)
  );
  al_ao21ttf _2494_ (
    .a(N273),
    .b(N239),
    .c(_1031_),
    .y(_1032_)
  );
  al_ao21 _2495_ (
    .a(_1032_),
    .b(_1030_),
    .c(_0952_),
    .y(_1033_)
  );
  al_nand2 _2496_ (
    .a(N273),
    .b(N239),
    .y(_1034_)
  );
  al_nand3fft _2497_ (
    .a(_0885_),
    .b(_1031_),
    .c(_1034_),
    .y(_1035_)
  );
  al_and3 _2498_ (
    .a(_1028_),
    .b(_1035_),
    .c(_1033_),
    .y(_1036_)
  );
  al_ao21 _2499_ (
    .a(_1035_),
    .b(_1033_),
    .c(_1028_),
    .y(_1037_)
  );
  al_nand3fft _2500_ (
    .a(_1036_),
    .b(_1027_),
    .c(_1037_),
    .y(_1038_)
  );
  al_ao21ttf _2501_ (
    .a(_0951_),
    .b(_0957_),
    .c(_0955_),
    .y(_1039_)
  );
  al_nand3 _2502_ (
    .a(_1028_),
    .b(_1035_),
    .c(_1033_),
    .y(_1040_)
  );
  al_ao21 _2503_ (
    .a(_1040_),
    .b(_1037_),
    .c(_1039_),
    .y(_1041_)
  );
  al_and3 _2504_ (
    .a(_1026_),
    .b(_1038_),
    .c(_1041_),
    .y(_1042_)
  );
  al_ao21 _2505_ (
    .a(_1038_),
    .b(_1041_),
    .c(_1026_),
    .y(_1043_)
  );
  al_and3ftt _2506_ (
    .a(_1042_),
    .b(_1025_),
    .c(_1043_),
    .y(_1044_)
  );
  al_nand3 _2507_ (
    .a(_1026_),
    .b(_1038_),
    .c(_1041_),
    .y(_1045_)
  );
  al_ao21 _2508_ (
    .a(_1045_),
    .b(_1043_),
    .c(_1025_),
    .y(_1046_)
  );
  al_nor3fft _2509_ (
    .a(_1024_),
    .b(_1046_),
    .c(_1044_),
    .y(_1047_)
  );
  al_nand3ftt _2510_ (
    .a(_1042_),
    .b(_1025_),
    .c(_1043_),
    .y(_1048_)
  );
  al_ao21 _2511_ (
    .a(_1046_),
    .b(_1048_),
    .c(_1024_),
    .y(_1049_)
  );
  al_and3ftt _2512_ (
    .a(_1047_),
    .b(_1023_),
    .c(_1049_),
    .y(_1050_)
  );
  al_nand3 _2513_ (
    .a(_1024_),
    .b(_1046_),
    .c(_1048_),
    .y(_1051_)
  );
  al_ao21 _2514_ (
    .a(_1051_),
    .b(_1049_),
    .c(_1023_),
    .y(_1052_)
  );
  al_nor3fft _2515_ (
    .a(_1022_),
    .b(_1052_),
    .c(_1050_),
    .y(_1053_)
  );
  al_nand3ftt _2516_ (
    .a(_1047_),
    .b(_1023_),
    .c(_1049_),
    .y(_1054_)
  );
  al_ao21 _2517_ (
    .a(_1052_),
    .b(_1054_),
    .c(_1022_),
    .y(_1055_)
  );
  al_and3ftt _2518_ (
    .a(_1053_),
    .b(_1021_),
    .c(_1055_),
    .y(_1056_)
  );
  al_nand3 _2519_ (
    .a(_1022_),
    .b(_1052_),
    .c(_1054_),
    .y(_1057_)
  );
  al_ao21 _2520_ (
    .a(_1057_),
    .b(_1055_),
    .c(_1021_),
    .y(_1058_)
  );
  al_nor3fft _2521_ (
    .a(_1020_),
    .b(_1058_),
    .c(_1056_),
    .y(_1059_)
  );
  al_nand3ftt _2522_ (
    .a(_1053_),
    .b(_1021_),
    .c(_1055_),
    .y(_1060_)
  );
  al_ao21 _2523_ (
    .a(_1058_),
    .b(_1060_),
    .c(_1020_),
    .y(_1061_)
  );
  al_and3ftt _2524_ (
    .a(_1059_),
    .b(_1061_),
    .c(_1019_),
    .y(_1062_)
  );
  al_nand3 _2525_ (
    .a(_1020_),
    .b(_1058_),
    .c(_1060_),
    .y(_1063_)
  );
  al_ao21 _2526_ (
    .a(_1063_),
    .b(_1061_),
    .c(_1019_),
    .y(_1064_)
  );
  al_nor3fft _2527_ (
    .a(_1018_),
    .b(_1064_),
    .c(_1062_),
    .y(_1066_)
  );
  al_nand3ftt _2528_ (
    .a(_1059_),
    .b(_1061_),
    .c(_1019_),
    .y(_1067_)
  );
  al_ao21 _2529_ (
    .a(_1064_),
    .b(_1067_),
    .c(_1018_),
    .y(_1068_)
  );
  al_and3ftt _2530_ (
    .a(_1066_),
    .b(_1017_),
    .c(_1068_),
    .y(_1069_)
  );
  al_nand3 _2531_ (
    .a(_1018_),
    .b(_1064_),
    .c(_1067_),
    .y(_1070_)
  );
  al_ao21 _2532_ (
    .a(_1070_),
    .b(_1068_),
    .c(_1017_),
    .y(_1071_)
  );
  al_nor3fft _2533_ (
    .a(_1016_),
    .b(_1071_),
    .c(_1069_),
    .y(_1072_)
  );
  al_nand3ftt _2534_ (
    .a(_1066_),
    .b(_1017_),
    .c(_1068_),
    .y(_1073_)
  );
  al_ao21 _2535_ (
    .a(_1071_),
    .b(_1073_),
    .c(_1016_),
    .y(_1074_)
  );
  al_and3ftt _2536_ (
    .a(_1072_),
    .b(_1074_),
    .c(_1015_),
    .y(_1075_)
  );
  al_nand3 _2537_ (
    .a(_1016_),
    .b(_1071_),
    .c(_1073_),
    .y(_1077_)
  );
  al_ao21 _2538_ (
    .a(_1077_),
    .b(_1074_),
    .c(_1015_),
    .y(_1078_)
  );
  al_nor3fft _2539_ (
    .a(_1014_),
    .b(_1078_),
    .c(_1075_),
    .y(_1079_)
  );
  al_nand3ftt _2540_ (
    .a(_1072_),
    .b(_1074_),
    .c(_1015_),
    .y(_1080_)
  );
  al_ao21 _2541_ (
    .a(_1078_),
    .b(_1080_),
    .c(_1014_),
    .y(_1081_)
  );
  al_and3ftt _2542_ (
    .a(_1079_),
    .b(_1081_),
    .c(_1013_),
    .y(_1082_)
  );
  al_nand3 _2543_ (
    .a(_1014_),
    .b(_1078_),
    .c(_1080_),
    .y(_1083_)
  );
  al_ao21 _2544_ (
    .a(_1083_),
    .b(_1081_),
    .c(_1013_),
    .y(_1084_)
  );
  al_nor3fft _2545_ (
    .a(_1012_),
    .b(_1084_),
    .c(_1082_),
    .y(_1085_)
  );
  al_nand3ftt _2546_ (
    .a(_1079_),
    .b(_1081_),
    .c(_1013_),
    .y(_1086_)
  );
  al_ao21 _2547_ (
    .a(_1084_),
    .b(_1086_),
    .c(_1012_),
    .y(_1088_)
  );
  al_and3ftt _2548_ (
    .a(_1085_),
    .b(_1088_),
    .c(_1011_),
    .y(_1089_)
  );
  al_nand3 _2549_ (
    .a(_1012_),
    .b(_1084_),
    .c(_1086_),
    .y(_1090_)
  );
  al_ao21 _2550_ (
    .a(_1090_),
    .b(_1088_),
    .c(_1011_),
    .y(_1091_)
  );
  al_nor3fft _2551_ (
    .a(_1010_),
    .b(_1091_),
    .c(_1089_),
    .y(_1092_)
  );
  al_nand3ftt _2552_ (
    .a(_1085_),
    .b(_1088_),
    .c(_1011_),
    .y(_1093_)
  );
  al_ao21 _2553_ (
    .a(_1091_),
    .b(_1093_),
    .c(_1010_),
    .y(_1094_)
  );
  al_and3ftt _2554_ (
    .a(_1092_),
    .b(_1094_),
    .c(_1009_),
    .y(_1095_)
  );
  al_nand3 _2555_ (
    .a(_1010_),
    .b(_1091_),
    .c(_1093_),
    .y(_1096_)
  );
  al_ao21 _2556_ (
    .a(_1096_),
    .b(_1094_),
    .c(_1009_),
    .y(_1097_)
  );
  al_nor3fft _2557_ (
    .a(_1008_),
    .b(_1097_),
    .c(_1095_),
    .y(_1099_)
  );
  al_nand3ftt _2558_ (
    .a(_1092_),
    .b(_1094_),
    .c(_1009_),
    .y(_1100_)
  );
  al_ao21 _2559_ (
    .a(_1097_),
    .b(_1100_),
    .c(_1008_),
    .y(_1101_)
  );
  al_nand3ftt _2560_ (
    .a(_1099_),
    .b(_1101_),
    .c(_1007_),
    .y(_1102_)
  );
  al_nand3 _2561_ (
    .a(_1008_),
    .b(_1097_),
    .c(_1100_),
    .y(_1103_)
  );
  al_ao21 _2562_ (
    .a(_1103_),
    .b(_1101_),
    .c(_1007_),
    .y(_1104_)
  );
  al_nand3 _2563_ (
    .a(_1006_),
    .b(_1104_),
    .c(_1102_),
    .y(_1105_)
  );
  al_ao21 _2564_ (
    .a(_1104_),
    .b(_1102_),
    .c(_1006_),
    .y(_1106_)
  );
  al_and3 _2565_ (
    .a(_1105_),
    .b(_1106_),
    .c(_1005_),
    .y(_1107_)
  );
  al_ao21 _2566_ (
    .a(_1105_),
    .b(_1106_),
    .c(_1005_),
    .y(_1108_)
  );
  al_nor3fft _2567_ (
    .a(_1004_),
    .b(_1108_),
    .c(_1107_),
    .y(_1109_)
  );
  al_oai21ftf _2568_ (
    .a(_1108_),
    .b(_1107_),
    .c(_1004_),
    .y(_1110_)
  );
  al_nand2ft _2569_ (
    .a(_1109_),
    .b(_1110_),
    .y(N5971)
  );
  al_nand2 _2570_ (
    .a(N1),
    .b(N528),
    .y(_1111_)
  );
  al_aoi21 _2571_ (
    .a(_1004_),
    .b(_1108_),
    .c(_1107_),
    .y(_1112_)
  );
  al_nand2 _2572_ (
    .a(N511),
    .b(N18),
    .y(_1113_)
  );
  al_and3ftt _2573_ (
    .a(_1099_),
    .b(_1101_),
    .c(_1007_),
    .y(_1114_)
  );
  al_ao21 _2574_ (
    .a(_1006_),
    .b(_1104_),
    .c(_1114_),
    .y(_1115_)
  );
  al_nand2 _2575_ (
    .a(N494),
    .b(N35),
    .y(_1116_)
  );
  al_ao21 _2576_ (
    .a(_1008_),
    .b(_1097_),
    .c(_1095_),
    .y(_1117_)
  );
  al_nand2 _2577_ (
    .a(N477),
    .b(N52),
    .y(_1119_)
  );
  al_ao21 _2578_ (
    .a(_1010_),
    .b(_1091_),
    .c(_1089_),
    .y(_1120_)
  );
  al_nand2 _2579_ (
    .a(N460),
    .b(N69),
    .y(_1121_)
  );
  al_ao21 _2580_ (
    .a(_1012_),
    .b(_1084_),
    .c(_1082_),
    .y(_1122_)
  );
  al_nand2 _2581_ (
    .a(N443),
    .b(N86),
    .y(_1123_)
  );
  al_ao21 _2582_ (
    .a(_1014_),
    .b(_1078_),
    .c(_1075_),
    .y(_1124_)
  );
  al_nand2 _2583_ (
    .a(N426),
    .b(N103),
    .y(_1125_)
  );
  al_ao21 _2584_ (
    .a(_1016_),
    .b(_1071_),
    .c(_1069_),
    .y(_1126_)
  );
  al_nand2 _2585_ (
    .a(N409),
    .b(N120),
    .y(_1127_)
  );
  al_ao21 _2586_ (
    .a(_1018_),
    .b(_1064_),
    .c(_1062_),
    .y(_1128_)
  );
  al_nand2 _2587_ (
    .a(N392),
    .b(N137),
    .y(_1130_)
  );
  al_ao21 _2588_ (
    .a(_1020_),
    .b(_1058_),
    .c(_1056_),
    .y(_1131_)
  );
  al_nand2 _2589_ (
    .a(N375),
    .b(N154),
    .y(_1132_)
  );
  al_ao21 _2590_ (
    .a(_1022_),
    .b(_1052_),
    .c(_1050_),
    .y(_1133_)
  );
  al_nand2 _2591_ (
    .a(N358),
    .b(N171),
    .y(_1134_)
  );
  al_ao21 _2592_ (
    .a(_1024_),
    .b(_1046_),
    .c(_1044_),
    .y(_1135_)
  );
  al_nand2 _2593_ (
    .a(N341),
    .b(N188),
    .y(_1136_)
  );
  al_and3ftt _2594_ (
    .a(_1036_),
    .b(_1039_),
    .c(_1037_),
    .y(_1137_)
  );
  al_ao21 _2595_ (
    .a(_1026_),
    .b(_1041_),
    .c(_1137_),
    .y(_1138_)
  );
  al_nand2 _2596_ (
    .a(N324),
    .b(N205),
    .y(_1139_)
  );
  al_ao21ttf _2597_ (
    .a(_1028_),
    .b(_1035_),
    .c(_1033_),
    .y(_1141_)
  );
  al_nand2 _2598_ (
    .a(N307),
    .b(N222),
    .y(_1142_)
  );
  al_nand3fft _2599_ (
    .a(N256),
    .b(_0956_),
    .c(_1029_),
    .y(_1143_)
  );
  al_nand2 _2600_ (
    .a(N273),
    .b(N256),
    .y(_1144_)
  );
  al_nand3ftt _2601_ (
    .a(N222),
    .b(N290),
    .c(N239),
    .y(_1145_)
  );
  al_mux2h _2602_ (
    .a(_1145_),
    .b(_1029_),
    .s(_1144_),
    .y(_1146_)
  );
  al_nand3 _2603_ (
    .a(_1142_),
    .b(_1143_),
    .c(_1146_),
    .y(_1147_)
  );
  al_ao21 _2604_ (
    .a(_1143_),
    .b(_1146_),
    .c(_1142_),
    .y(_1148_)
  );
  al_nand3 _2605_ (
    .a(_1147_),
    .b(_1148_),
    .c(_1141_),
    .y(_1149_)
  );
  al_ao21 _2606_ (
    .a(_1147_),
    .b(_1148_),
    .c(_1141_),
    .y(_1150_)
  );
  al_and3 _2607_ (
    .a(_1139_),
    .b(_1149_),
    .c(_1150_),
    .y(_1152_)
  );
  al_ao21 _2608_ (
    .a(_1149_),
    .b(_1150_),
    .c(_1139_),
    .y(_1153_)
  );
  al_nand3ftt _2609_ (
    .a(_1152_),
    .b(_1153_),
    .c(_1138_),
    .y(_1154_)
  );
  al_aoi21 _2610_ (
    .a(_1026_),
    .b(_1041_),
    .c(_1137_),
    .y(_1155_)
  );
  al_ao21ftf _2611_ (
    .a(_1152_),
    .b(_1153_),
    .c(_1155_),
    .y(_1156_)
  );
  al_nand3 _2612_ (
    .a(_1136_),
    .b(_1154_),
    .c(_1156_),
    .y(_1157_)
  );
  al_ao21 _2613_ (
    .a(_1154_),
    .b(_1156_),
    .c(_1136_),
    .y(_1158_)
  );
  al_nand3 _2614_ (
    .a(_1157_),
    .b(_1158_),
    .c(_1135_),
    .y(_1159_)
  );
  al_ao21 _2615_ (
    .a(_1157_),
    .b(_1158_),
    .c(_1135_),
    .y(_1160_)
  );
  al_and3 _2616_ (
    .a(_1134_),
    .b(_1159_),
    .c(_1160_),
    .y(_1161_)
  );
  al_ao21 _2617_ (
    .a(_1159_),
    .b(_1160_),
    .c(_1134_),
    .y(_1163_)
  );
  al_nand3ftt _2618_ (
    .a(_1161_),
    .b(_1163_),
    .c(_1133_),
    .y(_1164_)
  );
  al_nand3 _2619_ (
    .a(_1134_),
    .b(_1159_),
    .c(_1160_),
    .y(_1165_)
  );
  al_ao21 _2620_ (
    .a(_1165_),
    .b(_1163_),
    .c(_1133_),
    .y(_1166_)
  );
  al_and3 _2621_ (
    .a(_1132_),
    .b(_1164_),
    .c(_1166_),
    .y(_1167_)
  );
  al_ao21 _2622_ (
    .a(_1164_),
    .b(_1166_),
    .c(_1132_),
    .y(_1168_)
  );
  al_nand3ftt _2623_ (
    .a(_1167_),
    .b(_1168_),
    .c(_1131_),
    .y(_1169_)
  );
  al_nand3 _2624_ (
    .a(_1132_),
    .b(_1164_),
    .c(_1166_),
    .y(_1170_)
  );
  al_ao21 _2625_ (
    .a(_1170_),
    .b(_1168_),
    .c(_1131_),
    .y(_1171_)
  );
  al_and3 _2626_ (
    .a(_1130_),
    .b(_1169_),
    .c(_1171_),
    .y(_1172_)
  );
  al_ao21 _2627_ (
    .a(_1169_),
    .b(_1171_),
    .c(_1130_),
    .y(_1174_)
  );
  al_nand3ftt _2628_ (
    .a(_1172_),
    .b(_1174_),
    .c(_1128_),
    .y(_1175_)
  );
  al_nand3 _2629_ (
    .a(_1130_),
    .b(_1169_),
    .c(_1171_),
    .y(_1176_)
  );
  al_ao21 _2630_ (
    .a(_1176_),
    .b(_1174_),
    .c(_1128_),
    .y(_1177_)
  );
  al_and3 _2631_ (
    .a(_1127_),
    .b(_1175_),
    .c(_1177_),
    .y(_1178_)
  );
  al_ao21 _2632_ (
    .a(_1175_),
    .b(_1177_),
    .c(_1127_),
    .y(_1179_)
  );
  al_nand3ftt _2633_ (
    .a(_1178_),
    .b(_1179_),
    .c(_1126_),
    .y(_1180_)
  );
  al_nand3 _2634_ (
    .a(_1127_),
    .b(_1175_),
    .c(_1177_),
    .y(_1181_)
  );
  al_ao21 _2635_ (
    .a(_1181_),
    .b(_1179_),
    .c(_1126_),
    .y(_1182_)
  );
  al_and3 _2636_ (
    .a(_1125_),
    .b(_1180_),
    .c(_1182_),
    .y(_1183_)
  );
  al_ao21 _2637_ (
    .a(_1180_),
    .b(_1182_),
    .c(_1125_),
    .y(_1185_)
  );
  al_nand3ftt _2638_ (
    .a(_1183_),
    .b(_1185_),
    .c(_1124_),
    .y(_1186_)
  );
  al_nand3 _2639_ (
    .a(_1125_),
    .b(_1180_),
    .c(_1182_),
    .y(_1187_)
  );
  al_ao21 _2640_ (
    .a(_1187_),
    .b(_1185_),
    .c(_1124_),
    .y(_1188_)
  );
  al_and3 _2641_ (
    .a(_1123_),
    .b(_1186_),
    .c(_1188_),
    .y(_1189_)
  );
  al_ao21 _2642_ (
    .a(_1186_),
    .b(_1188_),
    .c(_1123_),
    .y(_1190_)
  );
  al_nand3ftt _2643_ (
    .a(_1189_),
    .b(_1190_),
    .c(_1122_),
    .y(_1191_)
  );
  al_nand3 _2644_ (
    .a(_1123_),
    .b(_1186_),
    .c(_1188_),
    .y(_1192_)
  );
  al_ao21 _2645_ (
    .a(_1192_),
    .b(_1190_),
    .c(_1122_),
    .y(_1193_)
  );
  al_and3 _2646_ (
    .a(_1121_),
    .b(_1191_),
    .c(_1193_),
    .y(_1194_)
  );
  al_ao21 _2647_ (
    .a(_1191_),
    .b(_1193_),
    .c(_1121_),
    .y(_1196_)
  );
  al_nand3ftt _2648_ (
    .a(_1194_),
    .b(_1196_),
    .c(_1120_),
    .y(_1197_)
  );
  al_nand3 _2649_ (
    .a(_1121_),
    .b(_1191_),
    .c(_1193_),
    .y(_1198_)
  );
  al_ao21 _2650_ (
    .a(_1198_),
    .b(_1196_),
    .c(_1120_),
    .y(_1199_)
  );
  al_and3 _2651_ (
    .a(_1119_),
    .b(_1197_),
    .c(_1199_),
    .y(_1200_)
  );
  al_ao21 _2652_ (
    .a(_1197_),
    .b(_1199_),
    .c(_1119_),
    .y(_1201_)
  );
  al_and3ftt _2653_ (
    .a(_1200_),
    .b(_1201_),
    .c(_1117_),
    .y(_1202_)
  );
  al_aoi21 _2654_ (
    .a(_1008_),
    .b(_1097_),
    .c(_1095_),
    .y(_1203_)
  );
  al_nand3 _2655_ (
    .a(_1119_),
    .b(_1197_),
    .c(_1199_),
    .y(_1204_)
  );
  al_ao21ttf _2656_ (
    .a(_1204_),
    .b(_1201_),
    .c(_1203_),
    .y(_1205_)
  );
  al_nor3fft _2657_ (
    .a(_1116_),
    .b(_1205_),
    .c(_1202_),
    .y(_1207_)
  );
  al_nand3ftt _2658_ (
    .a(_1200_),
    .b(_1201_),
    .c(_1117_),
    .y(_1208_)
  );
  al_ao21 _2659_ (
    .a(_1205_),
    .b(_1208_),
    .c(_1116_),
    .y(_1209_)
  );
  al_nand3ftt _2660_ (
    .a(_1207_),
    .b(_1209_),
    .c(_1115_),
    .y(_1210_)
  );
  al_aoi21 _2661_ (
    .a(_1006_),
    .b(_1104_),
    .c(_1114_),
    .y(_1211_)
  );
  al_nand3 _2662_ (
    .a(_1116_),
    .b(_1205_),
    .c(_1208_),
    .y(_1212_)
  );
  al_ao21ttf _2663_ (
    .a(_1212_),
    .b(_1209_),
    .c(_1211_),
    .y(_1213_)
  );
  al_nand3 _2664_ (
    .a(_1113_),
    .b(_1213_),
    .c(_1210_),
    .y(_1214_)
  );
  al_ao21 _2665_ (
    .a(_1213_),
    .b(_1210_),
    .c(_1113_),
    .y(_1215_)
  );
  al_nor3fft _2666_ (
    .a(_1214_),
    .b(_1215_),
    .c(_1112_),
    .y(_1216_)
  );
  al_ao21ttf _2667_ (
    .a(_1214_),
    .b(_1215_),
    .c(_1112_),
    .y(_1217_)
  );
  al_nor3fft _2668_ (
    .a(_1111_),
    .b(_1217_),
    .c(_1216_),
    .y(_1218_)
  );
  al_oai21ftf _2669_ (
    .a(_1217_),
    .b(_1216_),
    .c(_1111_),
    .y(_1219_)
  );
  al_nand2ft _2670_ (
    .a(_1218_),
    .b(_1219_),
    .y(N6123)
  );
  al_aoi21 _2671_ (
    .a(_1111_),
    .b(_1217_),
    .c(_1216_),
    .y(_1220_)
  );
  al_nand2 _2672_ (
    .a(N528),
    .b(N18),
    .y(_1221_)
  );
  al_and3ftt _2673_ (
    .a(_1207_),
    .b(_1209_),
    .c(_1115_),
    .y(_1222_)
  );
  al_ao21 _2674_ (
    .a(_1113_),
    .b(_1213_),
    .c(_1222_),
    .y(_1223_)
  );
  al_nand2 _2675_ (
    .a(N511),
    .b(N35),
    .y(_1224_)
  );
  al_ao21 _2676_ (
    .a(_1116_),
    .b(_1205_),
    .c(_1202_),
    .y(_1225_)
  );
  al_nand2 _2677_ (
    .a(N494),
    .b(N52),
    .y(_1227_)
  );
  al_ao21ttf _2678_ (
    .a(_1119_),
    .b(_1199_),
    .c(_1197_),
    .y(_1228_)
  );
  al_nand2 _2679_ (
    .a(N477),
    .b(N69),
    .y(_1229_)
  );
  al_ao21ttf _2680_ (
    .a(_1121_),
    .b(_1193_),
    .c(_1191_),
    .y(_1230_)
  );
  al_nand2 _2681_ (
    .a(N460),
    .b(N86),
    .y(_1231_)
  );
  al_ao21ttf _2682_ (
    .a(_1123_),
    .b(_1188_),
    .c(_1186_),
    .y(_1232_)
  );
  al_nand2 _2683_ (
    .a(N443),
    .b(N103),
    .y(_1233_)
  );
  al_ao21ttf _2684_ (
    .a(_1125_),
    .b(_1182_),
    .c(_1180_),
    .y(_1234_)
  );
  al_nand2 _2685_ (
    .a(N426),
    .b(N120),
    .y(_1235_)
  );
  al_ao21ttf _2686_ (
    .a(_1127_),
    .b(_1177_),
    .c(_1175_),
    .y(_1236_)
  );
  al_nand2 _2687_ (
    .a(N409),
    .b(N137),
    .y(_1238_)
  );
  al_ao21ttf _2688_ (
    .a(_1130_),
    .b(_1171_),
    .c(_1169_),
    .y(_1239_)
  );
  al_nand2 _2689_ (
    .a(N392),
    .b(N154),
    .y(_1240_)
  );
  al_ao21ttf _2690_ (
    .a(_1132_),
    .b(_1166_),
    .c(_1164_),
    .y(_1241_)
  );
  al_nand2 _2691_ (
    .a(N375),
    .b(N171),
    .y(_1242_)
  );
  al_ao21ttf _2692_ (
    .a(_1134_),
    .b(_1160_),
    .c(_1159_),
    .y(_1243_)
  );
  al_nand2 _2693_ (
    .a(N358),
    .b(N188),
    .y(_1244_)
  );
  al_ao21ttf _2694_ (
    .a(_1136_),
    .b(_1156_),
    .c(_1154_),
    .y(_1245_)
  );
  al_nand2 _2695_ (
    .a(N341),
    .b(N205),
    .y(_1246_)
  );
  al_ao21ttf _2696_ (
    .a(_1139_),
    .b(_1150_),
    .c(_1149_),
    .y(_1247_)
  );
  al_nand2 _2697_ (
    .a(N324),
    .b(N222),
    .y(_1249_)
  );
  al_ao21ttf _2698_ (
    .a(_1142_),
    .b(_1143_),
    .c(_1146_),
    .y(_1250_)
  );
  al_and2 _2699_ (
    .a(N290),
    .b(N256),
    .y(_1251_)
  );
  al_nand2 _2700_ (
    .a(N307),
    .b(N239),
    .y(_1252_)
  );
  al_nand3 _2701_ (
    .a(_1034_),
    .b(_1251_),
    .c(_1252_),
    .y(_1253_)
  );
  al_ao21 _2702_ (
    .a(_1034_),
    .b(_1251_),
    .c(_1252_),
    .y(_1254_)
  );
  al_nand3 _2703_ (
    .a(_1254_),
    .b(_1253_),
    .c(_1250_),
    .y(_1255_)
  );
  al_ao21 _2704_ (
    .a(_1253_),
    .b(_1254_),
    .c(_1250_),
    .y(_1256_)
  );
  al_nand3 _2705_ (
    .a(_1249_),
    .b(_1255_),
    .c(_1256_),
    .y(_1257_)
  );
  al_ao21 _2706_ (
    .a(_1255_),
    .b(_1256_),
    .c(_1249_),
    .y(_1258_)
  );
  al_nand3 _2707_ (
    .a(_1257_),
    .b(_1258_),
    .c(_1247_),
    .y(_1260_)
  );
  al_ao21 _2708_ (
    .a(_1257_),
    .b(_1258_),
    .c(_1247_),
    .y(_1261_)
  );
  al_nand3 _2709_ (
    .a(_1246_),
    .b(_1260_),
    .c(_1261_),
    .y(_1262_)
  );
  al_ao21 _2710_ (
    .a(_1260_),
    .b(_1261_),
    .c(_1246_),
    .y(_1263_)
  );
  al_nand3 _2711_ (
    .a(_1262_),
    .b(_1263_),
    .c(_1245_),
    .y(_1264_)
  );
  al_ao21 _2712_ (
    .a(_1262_),
    .b(_1263_),
    .c(_1245_),
    .y(_1265_)
  );
  al_and3 _2713_ (
    .a(_1244_),
    .b(_1264_),
    .c(_1265_),
    .y(_1266_)
  );
  al_ao21 _2714_ (
    .a(_1264_),
    .b(_1265_),
    .c(_1244_),
    .y(_1267_)
  );
  al_nand3ftt _2715_ (
    .a(_1266_),
    .b(_1267_),
    .c(_1243_),
    .y(_1268_)
  );
  al_ao21ftt _2716_ (
    .a(_1266_),
    .b(_1267_),
    .c(_1243_),
    .y(_1269_)
  );
  al_and3 _2717_ (
    .a(_1242_),
    .b(_1268_),
    .c(_1269_),
    .y(_1271_)
  );
  al_ao21 _2718_ (
    .a(_1268_),
    .b(_1269_),
    .c(_1242_),
    .y(_1272_)
  );
  al_nand3ftt _2719_ (
    .a(_1271_),
    .b(_1272_),
    .c(_1241_),
    .y(_1273_)
  );
  al_ao21ftt _2720_ (
    .a(_1271_),
    .b(_1272_),
    .c(_1241_),
    .y(_1274_)
  );
  al_and3 _2721_ (
    .a(_1240_),
    .b(_1273_),
    .c(_1274_),
    .y(_1275_)
  );
  al_ao21 _2722_ (
    .a(_1273_),
    .b(_1274_),
    .c(_1240_),
    .y(_1276_)
  );
  al_nand3ftt _2723_ (
    .a(_1275_),
    .b(_1276_),
    .c(_1239_),
    .y(_1277_)
  );
  al_ao21ftt _2724_ (
    .a(_1275_),
    .b(_1276_),
    .c(_1239_),
    .y(_1278_)
  );
  al_and3 _2725_ (
    .a(_1238_),
    .b(_1277_),
    .c(_1278_),
    .y(_1279_)
  );
  al_ao21 _2726_ (
    .a(_1277_),
    .b(_1278_),
    .c(_1238_),
    .y(_1280_)
  );
  al_nand3ftt _2727_ (
    .a(_1279_),
    .b(_1280_),
    .c(_1236_),
    .y(_1282_)
  );
  al_ao21ftt _2728_ (
    .a(_1279_),
    .b(_1280_),
    .c(_1236_),
    .y(_1283_)
  );
  al_and3 _2729_ (
    .a(_1235_),
    .b(_1282_),
    .c(_1283_),
    .y(_1284_)
  );
  al_ao21 _2730_ (
    .a(_1282_),
    .b(_1283_),
    .c(_1235_),
    .y(_1285_)
  );
  al_nand3ftt _2731_ (
    .a(_1284_),
    .b(_1285_),
    .c(_1234_),
    .y(_1286_)
  );
  al_ao21ftt _2732_ (
    .a(_1284_),
    .b(_1285_),
    .c(_1234_),
    .y(_1287_)
  );
  al_and3 _2733_ (
    .a(_1233_),
    .b(_1286_),
    .c(_1287_),
    .y(_1288_)
  );
  al_ao21 _2734_ (
    .a(_1286_),
    .b(_1287_),
    .c(_1233_),
    .y(_1289_)
  );
  al_nand3ftt _2735_ (
    .a(_1288_),
    .b(_1289_),
    .c(_1232_),
    .y(_1290_)
  );
  al_ao21ftt _2736_ (
    .a(_1288_),
    .b(_1289_),
    .c(_1232_),
    .y(_1291_)
  );
  al_and3 _2737_ (
    .a(_1231_),
    .b(_1290_),
    .c(_1291_),
    .y(_1293_)
  );
  al_ao21 _2738_ (
    .a(_1290_),
    .b(_1291_),
    .c(_1231_),
    .y(_1294_)
  );
  al_nand3ftt _2739_ (
    .a(_1293_),
    .b(_1294_),
    .c(_1230_),
    .y(_1295_)
  );
  al_ao21ftt _2740_ (
    .a(_1293_),
    .b(_1294_),
    .c(_1230_),
    .y(_1296_)
  );
  al_and3 _2741_ (
    .a(_1229_),
    .b(_1295_),
    .c(_1296_),
    .y(_1297_)
  );
  al_ao21 _2742_ (
    .a(_1295_),
    .b(_1296_),
    .c(_1229_),
    .y(_1298_)
  );
  al_nand3ftt _2743_ (
    .a(_1297_),
    .b(_1298_),
    .c(_1228_),
    .y(_1299_)
  );
  al_ao21ftt _2744_ (
    .a(_1297_),
    .b(_1298_),
    .c(_1228_),
    .y(_1300_)
  );
  al_and3 _2745_ (
    .a(_1227_),
    .b(_1299_),
    .c(_1300_),
    .y(_1301_)
  );
  al_ao21 _2746_ (
    .a(_1299_),
    .b(_1300_),
    .c(_1227_),
    .y(_1302_)
  );
  al_nand3ftt _2747_ (
    .a(_1301_),
    .b(_1302_),
    .c(_1225_),
    .y(_1304_)
  );
  al_ao21ftt _2748_ (
    .a(_1301_),
    .b(_1302_),
    .c(_1225_),
    .y(_1305_)
  );
  al_and3 _2749_ (
    .a(_1224_),
    .b(_1304_),
    .c(_1305_),
    .y(_1306_)
  );
  al_ao21 _2750_ (
    .a(_1304_),
    .b(_1305_),
    .c(_1224_),
    .y(_1307_)
  );
  al_nand3ftt _2751_ (
    .a(_1306_),
    .b(_1307_),
    .c(_1223_),
    .y(_1308_)
  );
  al_aoi21 _2752_ (
    .a(_1113_),
    .b(_1213_),
    .c(_1222_),
    .y(_1309_)
  );
  al_nand3 _2753_ (
    .a(_1224_),
    .b(_1304_),
    .c(_1305_),
    .y(_1310_)
  );
  al_ao21ttf _2754_ (
    .a(_1310_),
    .b(_1307_),
    .c(_1309_),
    .y(_1311_)
  );
  al_nand3 _2755_ (
    .a(_1221_),
    .b(_1311_),
    .c(_1308_),
    .y(_1312_)
  );
  al_ao21 _2756_ (
    .a(_1311_),
    .b(_1308_),
    .c(_1221_),
    .y(_1313_)
  );
  al_ao21ttf _2757_ (
    .a(_1312_),
    .b(_1313_),
    .c(_1220_),
    .y(_1315_)
  );
  al_ao21ttf _2758_ (
    .a(_1221_),
    .b(_1311_),
    .c(_1308_),
    .y(_1316_)
  );
  al_nand2 _2759_ (
    .a(N528),
    .b(N35),
    .y(_1317_)
  );
  al_aoi21ttf _2760_ (
    .a(_1224_),
    .b(_1305_),
    .c(_1304_),
    .y(_1318_)
  );
  al_nand2 _2761_ (
    .a(N511),
    .b(N52),
    .y(_1319_)
  );
  al_aoi21ttf _2762_ (
    .a(_1227_),
    .b(_1300_),
    .c(_1299_),
    .y(_1320_)
  );
  al_nand2 _2763_ (
    .a(N494),
    .b(N69),
    .y(_1321_)
  );
  al_aoi21ttf _2764_ (
    .a(_1229_),
    .b(_1296_),
    .c(_1295_),
    .y(_1322_)
  );
  al_nand2 _2765_ (
    .a(N477),
    .b(N86),
    .y(_1323_)
  );
  al_aoi21ttf _2766_ (
    .a(_1231_),
    .b(_1291_),
    .c(_1290_),
    .y(_1324_)
  );
  al_nand2 _2767_ (
    .a(N460),
    .b(N103),
    .y(_1326_)
  );
  al_aoi21ttf _2768_ (
    .a(_1233_),
    .b(_1287_),
    .c(_1286_),
    .y(_1327_)
  );
  al_nand2 _2769_ (
    .a(N443),
    .b(N120),
    .y(_1328_)
  );
  al_aoi21ttf _2770_ (
    .a(_1235_),
    .b(_1283_),
    .c(_1282_),
    .y(_1329_)
  );
  al_nand2 _2771_ (
    .a(N426),
    .b(N137),
    .y(_1330_)
  );
  al_aoi21ttf _2772_ (
    .a(_1238_),
    .b(_1278_),
    .c(_1277_),
    .y(_1331_)
  );
  al_nand2 _2773_ (
    .a(N409),
    .b(N154),
    .y(_1332_)
  );
  al_aoi21ttf _2774_ (
    .a(_1240_),
    .b(_1274_),
    .c(_1273_),
    .y(_1333_)
  );
  al_nand2 _2775_ (
    .a(N392),
    .b(N171),
    .y(_1334_)
  );
  al_aoi21ttf _2776_ (
    .a(_1242_),
    .b(_1269_),
    .c(_1268_),
    .y(_1335_)
  );
  al_nand2 _2777_ (
    .a(N375),
    .b(N188),
    .y(_1337_)
  );
  al_ao21ttf _2778_ (
    .a(_1244_),
    .b(_1265_),
    .c(_1264_),
    .y(_1338_)
  );
  al_nand2 _2779_ (
    .a(N358),
    .b(N205),
    .y(_1339_)
  );
  al_ao21ttf _2780_ (
    .a(_1246_),
    .b(_1261_),
    .c(_1260_),
    .y(_1340_)
  );
  al_nand2 _2781_ (
    .a(N341),
    .b(N222),
    .y(_1341_)
  );
  al_ao21ttf _2782_ (
    .a(_1249_),
    .b(_1256_),
    .c(_1255_),
    .y(_1342_)
  );
  al_nand2 _2783_ (
    .a(N324),
    .b(N239),
    .y(_1343_)
  );
  al_inv _2784_ (
    .a(N256),
    .y(_1344_)
  );
  al_ao21ttf _2785_ (
    .a(_1034_),
    .b(_1252_),
    .c(_1251_),
    .y(_1345_)
  );
  al_ao21ftf _2786_ (
    .a(_1344_),
    .b(N307),
    .c(_1345_),
    .y(_1346_)
  );
  al_or3fft _2787_ (
    .a(N307),
    .b(N256),
    .c(_1345_),
    .y(_1348_)
  );
  al_nand3 _2788_ (
    .a(_1343_),
    .b(_1346_),
    .c(_1348_),
    .y(_1349_)
  );
  al_ao21 _2789_ (
    .a(_1346_),
    .b(_1348_),
    .c(_1343_),
    .y(_1350_)
  );
  al_nand3 _2790_ (
    .a(_1349_),
    .b(_1350_),
    .c(_1342_),
    .y(_1351_)
  );
  al_ao21 _2791_ (
    .a(_1349_),
    .b(_1350_),
    .c(_1342_),
    .y(_1352_)
  );
  al_nand3 _2792_ (
    .a(_1341_),
    .b(_1351_),
    .c(_1352_),
    .y(_1353_)
  );
  al_ao21 _2793_ (
    .a(_1351_),
    .b(_1352_),
    .c(_1341_),
    .y(_1354_)
  );
  al_nand3 _2794_ (
    .a(_1353_),
    .b(_1354_),
    .c(_1340_),
    .y(_1355_)
  );
  al_ao21 _2795_ (
    .a(_1353_),
    .b(_1354_),
    .c(_1340_),
    .y(_1356_)
  );
  al_nand3 _2796_ (
    .a(_1339_),
    .b(_1355_),
    .c(_1356_),
    .y(_1357_)
  );
  al_ao21 _2797_ (
    .a(_1355_),
    .b(_1356_),
    .c(_1339_),
    .y(_1359_)
  );
  al_nand3 _2798_ (
    .a(_1357_),
    .b(_1359_),
    .c(_1338_),
    .y(_1360_)
  );
  al_ao21 _2799_ (
    .a(_1357_),
    .b(_1359_),
    .c(_1338_),
    .y(_1361_)
  );
  al_nand3 _2800_ (
    .a(_1337_),
    .b(_1360_),
    .c(_1361_),
    .y(_1362_)
  );
  al_ao21 _2801_ (
    .a(_1360_),
    .b(_1361_),
    .c(_1337_),
    .y(_1363_)
  );
  al_or3fft _2802_ (
    .a(_1362_),
    .b(_1363_),
    .c(_1335_),
    .y(_1364_)
  );
  al_ao21ttf _2803_ (
    .a(_1362_),
    .b(_1363_),
    .c(_1335_),
    .y(_1365_)
  );
  al_nand3 _2804_ (
    .a(_1334_),
    .b(_1365_),
    .c(_1364_),
    .y(_1366_)
  );
  al_ao21 _2805_ (
    .a(_1365_),
    .b(_1364_),
    .c(_1334_),
    .y(_1367_)
  );
  al_or3fft _2806_ (
    .a(_1366_),
    .b(_1367_),
    .c(_1333_),
    .y(_1368_)
  );
  al_ao21ttf _2807_ (
    .a(_1366_),
    .b(_1367_),
    .c(_1333_),
    .y(_1370_)
  );
  al_nand3 _2808_ (
    .a(_1332_),
    .b(_1370_),
    .c(_1368_),
    .y(_1371_)
  );
  al_ao21 _2809_ (
    .a(_1370_),
    .b(_1368_),
    .c(_1332_),
    .y(_1372_)
  );
  al_or3fft _2810_ (
    .a(_1371_),
    .b(_1372_),
    .c(_1331_),
    .y(_1373_)
  );
  al_ao21ttf _2811_ (
    .a(_1371_),
    .b(_1372_),
    .c(_1331_),
    .y(_1374_)
  );
  al_nand3 _2812_ (
    .a(_1330_),
    .b(_1374_),
    .c(_1373_),
    .y(_1375_)
  );
  al_ao21 _2813_ (
    .a(_1374_),
    .b(_1373_),
    .c(_1330_),
    .y(_1376_)
  );
  al_or3fft _2814_ (
    .a(_1375_),
    .b(_1376_),
    .c(_1329_),
    .y(_1377_)
  );
  al_ao21ttf _2815_ (
    .a(_1375_),
    .b(_1376_),
    .c(_1329_),
    .y(_1378_)
  );
  al_nand3 _2816_ (
    .a(_1328_),
    .b(_1378_),
    .c(_1377_),
    .y(_1379_)
  );
  al_ao21 _2817_ (
    .a(_1378_),
    .b(_1377_),
    .c(_1328_),
    .y(_1380_)
  );
  al_or3fft _2818_ (
    .a(_1379_),
    .b(_1380_),
    .c(_1327_),
    .y(_1381_)
  );
  al_ao21ttf _2819_ (
    .a(_1379_),
    .b(_1380_),
    .c(_1327_),
    .y(_1382_)
  );
  al_nand3 _2820_ (
    .a(_1326_),
    .b(_1382_),
    .c(_1381_),
    .y(_1383_)
  );
  al_ao21 _2821_ (
    .a(_1382_),
    .b(_1381_),
    .c(_1326_),
    .y(_1384_)
  );
  al_or3fft _2822_ (
    .a(_1383_),
    .b(_1384_),
    .c(_1324_),
    .y(_1385_)
  );
  al_ao21ttf _2823_ (
    .a(_1383_),
    .b(_1384_),
    .c(_1324_),
    .y(_1386_)
  );
  al_nand3 _2824_ (
    .a(_1323_),
    .b(_1386_),
    .c(_1385_),
    .y(_1387_)
  );
  al_ao21 _2825_ (
    .a(_1386_),
    .b(_1385_),
    .c(_1323_),
    .y(_1388_)
  );
  al_or3fft _2826_ (
    .a(_1387_),
    .b(_1388_),
    .c(_1322_),
    .y(_1389_)
  );
  al_ao21ttf _2827_ (
    .a(_1387_),
    .b(_1388_),
    .c(_1322_),
    .y(_1391_)
  );
  al_nand3 _2828_ (
    .a(_1321_),
    .b(_1391_),
    .c(_1389_),
    .y(_1392_)
  );
  al_ao21 _2829_ (
    .a(_1391_),
    .b(_1389_),
    .c(_1321_),
    .y(_1393_)
  );
  al_or3fft _2830_ (
    .a(_1392_),
    .b(_1393_),
    .c(_1320_),
    .y(_1394_)
  );
  al_ao21ttf _2831_ (
    .a(_1392_),
    .b(_1393_),
    .c(_1320_),
    .y(_1395_)
  );
  al_nand3 _2832_ (
    .a(_1319_),
    .b(_1395_),
    .c(_1394_),
    .y(_1396_)
  );
  al_ao21 _2833_ (
    .a(_1395_),
    .b(_1394_),
    .c(_1319_),
    .y(_1397_)
  );
  al_or3fft _2834_ (
    .a(_1396_),
    .b(_1397_),
    .c(_1318_),
    .y(_1398_)
  );
  al_ao21ttf _2835_ (
    .a(_1396_),
    .b(_1397_),
    .c(_1318_),
    .y(_1399_)
  );
  al_and3 _2836_ (
    .a(_1317_),
    .b(_1399_),
    .c(_1398_),
    .y(_1400_)
  );
  al_ao21 _2837_ (
    .a(_1399_),
    .b(_1398_),
    .c(_1317_),
    .y(_1402_)
  );
  al_and3ftt _2838_ (
    .a(_1400_),
    .b(_1402_),
    .c(_1316_),
    .y(_1403_)
  );
  al_ao21ftt _2839_ (
    .a(_1400_),
    .b(_1402_),
    .c(_1316_),
    .y(_1404_)
  );
  al_nand3ftt _2840_ (
    .a(_1403_),
    .b(_1315_),
    .c(_1404_),
    .y(_1405_)
  );
  al_oa21ftf _2841_ (
    .a(_1404_),
    .b(_1403_),
    .c(_1315_),
    .y(_1406_)
  );
  al_or2ft _2842_ (
    .a(_1405_),
    .b(_1406_),
    .y(N6160)
  );
  al_ao21 _2843_ (
    .a(_1404_),
    .b(_1315_),
    .c(_1403_),
    .y(_1407_)
  );
  al_ao21ttf _2844_ (
    .a(_1317_),
    .b(_1399_),
    .c(_1398_),
    .y(_1408_)
  );
  al_nand2 _2845_ (
    .a(N528),
    .b(N52),
    .y(_1409_)
  );
  al_ao21ttf _2846_ (
    .a(_1319_),
    .b(_1395_),
    .c(_1394_),
    .y(_1410_)
  );
  al_nand2 _2847_ (
    .a(N511),
    .b(N69),
    .y(_1412_)
  );
  al_ao21ttf _2848_ (
    .a(_1321_),
    .b(_1391_),
    .c(_1389_),
    .y(_1413_)
  );
  al_nand2 _2849_ (
    .a(N494),
    .b(N86),
    .y(_1414_)
  );
  al_ao21ttf _2850_ (
    .a(_1323_),
    .b(_1386_),
    .c(_1385_),
    .y(_1415_)
  );
  al_nand2 _2851_ (
    .a(N477),
    .b(N103),
    .y(_1416_)
  );
  al_ao21ttf _2852_ (
    .a(_1326_),
    .b(_1382_),
    .c(_1381_),
    .y(_1417_)
  );
  al_nand2 _2853_ (
    .a(N460),
    .b(N120),
    .y(_1418_)
  );
  al_ao21ttf _2854_ (
    .a(_1328_),
    .b(_1378_),
    .c(_1377_),
    .y(_1419_)
  );
  al_nand2 _2855_ (
    .a(N443),
    .b(N137),
    .y(_1420_)
  );
  al_ao21ttf _2856_ (
    .a(_1330_),
    .b(_1374_),
    .c(_1373_),
    .y(_1421_)
  );
  al_nand2 _2857_ (
    .a(N426),
    .b(N154),
    .y(_1423_)
  );
  al_ao21ttf _2858_ (
    .a(_1332_),
    .b(_1370_),
    .c(_1368_),
    .y(_1424_)
  );
  al_nand2 _2859_ (
    .a(N409),
    .b(N171),
    .y(_1425_)
  );
  al_ao21ttf _2860_ (
    .a(_1334_),
    .b(_1365_),
    .c(_1364_),
    .y(_1426_)
  );
  al_nand2 _2861_ (
    .a(N392),
    .b(N188),
    .y(_1427_)
  );
  al_ao21ttf _2862_ (
    .a(_1337_),
    .b(_1361_),
    .c(_1360_),
    .y(_1428_)
  );
  al_nand2 _2863_ (
    .a(N375),
    .b(N205),
    .y(_1429_)
  );
  al_ao21ttf _2864_ (
    .a(_1339_),
    .b(_1356_),
    .c(_1355_),
    .y(_1430_)
  );
  al_nand2 _2865_ (
    .a(N358),
    .b(N222),
    .y(_1431_)
  );
  al_ao21ttf _2866_ (
    .a(_1341_),
    .b(_1352_),
    .c(_1351_),
    .y(_1432_)
  );
  al_nand2 _2867_ (
    .a(N341),
    .b(N239),
    .y(_1434_)
  );
  al_ao21ttf _2868_ (
    .a(_1343_),
    .b(_1348_),
    .c(_1346_),
    .y(_1435_)
  );
  al_ao21ftf _2869_ (
    .a(_1344_),
    .b(N324),
    .c(_1435_),
    .y(_1436_)
  );
  al_or3fft _2870_ (
    .a(N324),
    .b(N256),
    .c(_1435_),
    .y(_1437_)
  );
  al_nand3 _2871_ (
    .a(_1434_),
    .b(_1436_),
    .c(_1437_),
    .y(_1438_)
  );
  al_ao21 _2872_ (
    .a(_1436_),
    .b(_1437_),
    .c(_1434_),
    .y(_1439_)
  );
  al_nand3 _2873_ (
    .a(_1438_),
    .b(_1439_),
    .c(_1432_),
    .y(_1440_)
  );
  al_ao21 _2874_ (
    .a(_1438_),
    .b(_1439_),
    .c(_1432_),
    .y(_1441_)
  );
  al_nand3 _2875_ (
    .a(_1431_),
    .b(_1440_),
    .c(_1441_),
    .y(_1442_)
  );
  al_ao21 _2876_ (
    .a(_1440_),
    .b(_1441_),
    .c(_1431_),
    .y(_1443_)
  );
  al_nand3 _2877_ (
    .a(_1442_),
    .b(_1443_),
    .c(_1430_),
    .y(_0001_)
  );
  al_ao21 _2878_ (
    .a(_1442_),
    .b(_1443_),
    .c(_1430_),
    .y(_0002_)
  );
  al_nand3 _2879_ (
    .a(_1429_),
    .b(_0001_),
    .c(_0002_),
    .y(_0003_)
  );
  al_ao21 _2880_ (
    .a(_0001_),
    .b(_0002_),
    .c(_1429_),
    .y(_0004_)
  );
  al_nand3 _2881_ (
    .a(_0003_),
    .b(_0004_),
    .c(_1428_),
    .y(_0005_)
  );
  al_ao21 _2882_ (
    .a(_0003_),
    .b(_0004_),
    .c(_1428_),
    .y(_0006_)
  );
  al_nand3 _2883_ (
    .a(_1427_),
    .b(_0005_),
    .c(_0006_),
    .y(_0007_)
  );
  al_ao21 _2884_ (
    .a(_0005_),
    .b(_0006_),
    .c(_1427_),
    .y(_0008_)
  );
  al_nand3 _2885_ (
    .a(_0007_),
    .b(_0008_),
    .c(_1426_),
    .y(_0009_)
  );
  al_ao21 _2886_ (
    .a(_0007_),
    .b(_0008_),
    .c(_1426_),
    .y(_0010_)
  );
  al_nand3 _2887_ (
    .a(_1425_),
    .b(_0009_),
    .c(_0010_),
    .y(_0012_)
  );
  al_ao21 _2888_ (
    .a(_0009_),
    .b(_0010_),
    .c(_1425_),
    .y(_0013_)
  );
  al_nand3 _2889_ (
    .a(_0012_),
    .b(_0013_),
    .c(_1424_),
    .y(_0014_)
  );
  al_ao21 _2890_ (
    .a(_0012_),
    .b(_0013_),
    .c(_1424_),
    .y(_0015_)
  );
  al_nand3 _2891_ (
    .a(_1423_),
    .b(_0014_),
    .c(_0015_),
    .y(_0016_)
  );
  al_ao21 _2892_ (
    .a(_0014_),
    .b(_0015_),
    .c(_1423_),
    .y(_0017_)
  );
  al_nand3 _2893_ (
    .a(_0016_),
    .b(_0017_),
    .c(_1421_),
    .y(_0018_)
  );
  al_ao21 _2894_ (
    .a(_0016_),
    .b(_0017_),
    .c(_1421_),
    .y(_0019_)
  );
  al_nand3 _2895_ (
    .a(_1420_),
    .b(_0018_),
    .c(_0019_),
    .y(_0020_)
  );
  al_ao21 _2896_ (
    .a(_0018_),
    .b(_0019_),
    .c(_1420_),
    .y(_0021_)
  );
  al_nand3 _2897_ (
    .a(_0020_),
    .b(_0021_),
    .c(_1419_),
    .y(_0023_)
  );
  al_ao21 _2898_ (
    .a(_0020_),
    .b(_0021_),
    .c(_1419_),
    .y(_0024_)
  );
  al_nand3 _2899_ (
    .a(_1418_),
    .b(_0023_),
    .c(_0024_),
    .y(_0025_)
  );
  al_ao21 _2900_ (
    .a(_0023_),
    .b(_0024_),
    .c(_1418_),
    .y(_0026_)
  );
  al_nand3 _2901_ (
    .a(_0025_),
    .b(_0026_),
    .c(_1417_),
    .y(_0027_)
  );
  al_ao21 _2902_ (
    .a(_0025_),
    .b(_0026_),
    .c(_1417_),
    .y(_0028_)
  );
  al_nand3 _2903_ (
    .a(_1416_),
    .b(_0027_),
    .c(_0028_),
    .y(_0029_)
  );
  al_ao21 _2904_ (
    .a(_0027_),
    .b(_0028_),
    .c(_1416_),
    .y(_0030_)
  );
  al_nand3 _2905_ (
    .a(_0029_),
    .b(_0030_),
    .c(_1415_),
    .y(_0031_)
  );
  al_ao21 _2906_ (
    .a(_0029_),
    .b(_0030_),
    .c(_1415_),
    .y(_0032_)
  );
  al_nand3 _2907_ (
    .a(_1414_),
    .b(_0031_),
    .c(_0032_),
    .y(_0034_)
  );
  al_ao21 _2908_ (
    .a(_0031_),
    .b(_0032_),
    .c(_1414_),
    .y(_0035_)
  );
  al_nand3 _2909_ (
    .a(_0034_),
    .b(_0035_),
    .c(_1413_),
    .y(_0036_)
  );
  al_ao21 _2910_ (
    .a(_0034_),
    .b(_0035_),
    .c(_1413_),
    .y(_0037_)
  );
  al_nand3 _2911_ (
    .a(_1412_),
    .b(_0036_),
    .c(_0037_),
    .y(_0038_)
  );
  al_ao21 _2912_ (
    .a(_0036_),
    .b(_0037_),
    .c(_1412_),
    .y(_0039_)
  );
  al_nand3 _2913_ (
    .a(_0038_),
    .b(_0039_),
    .c(_1410_),
    .y(_0040_)
  );
  al_ao21 _2914_ (
    .a(_0038_),
    .b(_0039_),
    .c(_1410_),
    .y(_0041_)
  );
  al_and3 _2915_ (
    .a(_1409_),
    .b(_0040_),
    .c(_0041_),
    .y(_0042_)
  );
  al_ao21 _2916_ (
    .a(_0040_),
    .b(_0041_),
    .c(_1409_),
    .y(_0043_)
  );
  al_and3ftt _2917_ (
    .a(_0042_),
    .b(_0043_),
    .c(_1408_),
    .y(_0045_)
  );
  al_ao21ftt _2918_ (
    .a(_0042_),
    .b(_0043_),
    .c(_1408_),
    .y(_0046_)
  );
  al_nand3ftt _2919_ (
    .a(_0045_),
    .b(_0046_),
    .c(_1407_),
    .y(_0047_)
  );
  assign N6141 = N6150;
endmodule
