
module s38417(GND, VDD, CK, g1249, g16297, g16355, g16399, g16437, g16496, g1943, g24734, g25420, g25435, g25442, g25489, g26104, g26135, g26149, g2637, g27380, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, g3231, g3232, g3233, g3234, g3993, g4088, g4090, g4200, g4321, g4323, g4450, g4590, g51, g5388, g5437, g5472, g5511, g5549, g5555, g5595, g5612, g5629, g563, g5637, g5648, g5657, g5686, g5695, g5738, g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518, g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944, g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334, g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012, g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249, g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266, g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire _1886_;
  wire _1887_;
  wire _1888_;
  wire _1889_;
  wire _1890_;
  wire _1891_;
  wire _1892_;
  wire _1893_;
  wire _1894_;
  wire _1895_;
  wire _1896_;
  wire _1897_;
  wire _1898_;
  wire _1899_;
  wire _1900_;
  wire _1901_;
  wire _1902_;
  wire _1903_;
  wire _1904_;
  wire _1905_;
  wire _1906_;
  wire _1907_;
  wire _1908_;
  wire _1909_;
  wire _1910_;
  wire _1911_;
  wire _1912_;
  wire _1913_;
  wire _1914_;
  wire _1915_;
  wire _1916_;
  wire _1917_;
  wire _1918_;
  wire _1919_;
  wire _1920_;
  wire _1921_;
  wire _1922_;
  wire _1923_;
  wire _1924_;
  wire _1925_;
  wire _1926_;
  wire _1927_;
  wire _1928_;
  wire _1929_;
  wire _1930_;
  wire _1931_;
  wire _1932_;
  wire _1933_;
  wire _1934_;
  wire _1935_;
  wire _1936_;
  wire _1937_;
  wire _1938_;
  wire _1939_;
  wire _1940_;
  wire _1941_;
  wire _1942_;
  wire _1943_;
  wire _1944_;
  wire _1945_;
  wire _1946_;
  wire _1947_;
  wire _1948_;
  wire _1949_;
  wire _1950_;
  wire _1951_;
  wire _1952_;
  wire _1953_;
  wire _1954_;
  wire _1955_;
  wire _1956_;
  wire _1957_;
  wire _1958_;
  wire _1959_;
  wire _1960_;
  wire _1961_;
  wire _1962_;
  wire _1963_;
  wire _1964_;
  wire _1965_;
  wire _1966_;
  wire _1967_;
  wire _1968_;
  wire _1969_;
  wire _1970_;
  wire _1971_;
  wire _1972_;
  wire _1973_;
  wire _1974_;
  wire _1975_;
  wire _1976_;
  wire _1977_;
  wire _1978_;
  wire _1979_;
  wire _1980_;
  wire _1981_;
  wire _1982_;
  wire _1983_;
  wire _1984_;
  wire _1985_;
  wire _1986_;
  wire _1987_;
  wire _1988_;
  wire _1989_;
  wire _1990_;
  wire _1991_;
  wire _1992_;
  wire _1993_;
  wire _1994_;
  wire _1995_;
  wire _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  wire _2002_;
  wire _2003_;
  wire _2004_;
  wire _2005_;
  wire _2006_;
  wire _2007_;
  wire _2008_;
  wire _2009_;
  wire _2010_;
  wire _2011_;
  wire _2012_;
  wire _2013_;
  wire _2014_;
  wire _2015_;
  wire _2016_;
  wire _2017_;
  wire _2018_;
  wire _2019_;
  wire _2020_;
  wire _2021_;
  wire _2022_;
  wire _2023_;
  wire _2024_;
  wire _2025_;
  wire _2026_;
  wire _2027_;
  wire _2028_;
  wire _2029_;
  wire _2030_;
  wire _2031_;
  wire _2032_;
  wire _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire _2039_;
  wire _2040_;
  wire _2041_;
  wire _2042_;
  wire _2043_;
  wire _2044_;
  wire _2045_;
  wire _2046_;
  wire _2047_;
  wire _2048_;
  wire _2049_;
  wire _2050_;
  wire _2051_;
  wire _2052_;
  wire _2053_;
  wire _2054_;
  wire _2055_;
  wire _2056_;
  wire _2057_;
  wire _2058_;
  wire _2059_;
  wire _2060_;
  wire _2061_;
  wire _2062_;
  wire _2063_;
  wire _2064_;
  wire _2065_;
  wire _2066_;
  wire _2067_;
  wire _2068_;
  wire _2069_;
  wire _2070_;
  wire _2071_;
  wire _2072_;
  wire _2073_;
  wire _2074_;
  wire _2075_;
  wire _2076_;
  wire _2077_;
  wire _2078_;
  wire _2079_;
  wire _2080_;
  wire _2081_;
  wire _2082_;
  wire _2083_;
  wire _2084_;
  wire _2085_;
  wire _2086_;
  wire _2087_;
  wire _2088_;
  wire _2089_;
  wire _2090_;
  wire _2091_;
  wire _2092_;
  wire _2093_;
  wire _2094_;
  wire _2095_;
  wire _2096_;
  wire _2097_;
  wire _2098_;
  wire _2099_;
  wire _2100_;
  wire _2101_;
  wire _2102_;
  wire _2103_;
  wire _2104_;
  wire _2105_;
  wire _2106_;
  wire _2107_;
  wire _2108_;
  wire _2109_;
  wire _2110_;
  wire _2111_;
  wire _2112_;
  wire _2113_;
  wire _2114_;
  wire _2115_;
  wire _2116_;
  wire _2117_;
  wire _2118_;
  wire _2119_;
  wire _2120_;
  wire _2121_;
  wire _2122_;
  wire _2123_;
  wire _2124_;
  wire _2125_;
  wire _2126_;
  wire _2127_;
  wire _2128_;
  wire _2129_;
  wire _2130_;
  wire _2131_;
  wire _2132_;
  wire _2133_;
  wire _2134_;
  wire _2135_;
  wire _2136_;
  wire _2137_;
  wire _2138_;
  wire _2139_;
  wire _2140_;
  wire _2141_;
  wire _2142_;
  wire _2143_;
  wire _2144_;
  wire _2145_;
  wire _2146_;
  wire _2147_;
  wire _2148_;
  wire _2149_;
  wire _2150_;
  wire _2151_;
  wire _2152_;
  wire _2153_;
  wire _2154_;
  wire _2155_;
  wire _2156_;
  wire _2157_;
  wire _2158_;
  wire _2159_;
  wire _2160_;
  wire _2161_;
  wire _2162_;
  wire _2163_;
  wire _2164_;
  wire _2165_;
  wire _2166_;
  wire _2167_;
  wire _2168_;
  wire _2169_;
  wire _2170_;
  wire _2171_;
  wire _2172_;
  wire _2173_;
  wire _2174_;
  wire _2175_;
  wire _2176_;
  wire _2177_;
  wire _2178_;
  wire _2179_;
  wire _2180_;
  wire _2181_;
  wire _2182_;
  wire _2183_;
  wire _2184_;
  wire _2185_;
  wire _2186_;
  wire _2187_;
  wire _2188_;
  wire _2189_;
  wire _2190_;
  wire _2191_;
  wire _2192_;
  wire _2193_;
  wire _2194_;
  wire _2195_;
  wire _2196_;
  wire _2197_;
  wire _2198_;
  wire _2199_;
  wire _2200_;
  wire _2201_;
  wire _2202_;
  wire _2203_;
  wire _2204_;
  wire _2205_;
  wire _2206_;
  wire _2207_;
  wire _2208_;
  wire _2209_;
  wire _2210_;
  wire _2211_;
  wire _2212_;
  wire _2213_;
  wire _2214_;
  wire _2215_;
  wire _2216_;
  wire _2217_;
  wire _2218_;
  wire _2219_;
  wire _2220_;
  wire _2221_;
  wire _2222_;
  wire _2223_;
  wire _2224_;
  wire _2225_;
  wire _2226_;
  wire _2227_;
  wire _2228_;
  wire _2229_;
  wire _2230_;
  wire _2231_;
  wire _2232_;
  wire _2233_;
  wire _2234_;
  wire _2235_;
  wire _2236_;
  wire _2237_;
  wire _2238_;
  wire _2239_;
  wire _2240_;
  wire _2241_;
  wire _2242_;
  wire _2243_;
  wire _2244_;
  wire _2245_;
  wire _2246_;
  wire _2247_;
  wire _2248_;
  wire _2249_;
  wire _2250_;
  wire _2251_;
  wire _2252_;
  wire _2253_;
  wire _2254_;
  wire _2255_;
  wire _2256_;
  wire _2257_;
  wire _2258_;
  wire _2259_;
  wire _2260_;
  wire _2261_;
  wire _2262_;
  wire _2263_;
  wire _2264_;
  wire _2265_;
  wire _2266_;
  wire _2267_;
  wire _2268_;
  wire _2269_;
  wire _2270_;
  wire _2271_;
  wire _2272_;
  wire _2273_;
  wire _2274_;
  wire _2275_;
  wire _2276_;
  wire _2277_;
  wire _2278_;
  wire _2279_;
  wire _2280_;
  wire _2281_;
  wire _2282_;
  wire _2283_;
  wire _2284_;
  wire _2285_;
  wire _2286_;
  wire _2287_;
  wire _2288_;
  wire _2289_;
  wire _2290_;
  wire _2291_;
  wire _2292_;
  wire _2293_;
  wire _2294_;
  wire _2295_;
  wire _2296_;
  wire _2297_;
  wire _2298_;
  wire _2299_;
  wire _2300_;
  wire _2301_;
  wire _2302_;
  wire _2303_;
  wire _2304_;
  wire _2305_;
  wire _2306_;
  wire _2307_;
  wire _2308_;
  wire _2309_;
  wire _2310_;
  wire _2311_;
  wire _2312_;
  wire _2313_;
  wire _2314_;
  wire _2315_;
  wire _2316_;
  wire _2317_;
  wire _2318_;
  wire _2319_;
  wire _2320_;
  wire _2321_;
  wire _2322_;
  wire _2323_;
  wire _2324_;
  wire _2325_;
  wire _2326_;
  wire _2327_;
  wire _2328_;
  wire _2329_;
  wire _2330_;
  wire _2331_;
  wire _2332_;
  wire _2333_;
  wire _2334_;
  wire _2335_;
  wire _2336_;
  wire _2337_;
  wire _2338_;
  wire _2339_;
  wire _2340_;
  wire _2341_;
  wire _2342_;
  wire _2343_;
  wire _2344_;
  wire _2345_;
  wire _2346_;
  wire _2347_;
  wire _2348_;
  wire _2349_;
  wire _2350_;
  wire _2351_;
  wire _2352_;
  wire _2353_;
  wire _2354_;
  wire _2355_;
  wire _2356_;
  wire _2357_;
  wire _2358_;
  wire _2359_;
  wire _2360_;
  wire _2361_;
  wire _2362_;
  wire _2363_;
  wire _2364_;
  wire _2365_;
  wire _2366_;
  wire _2367_;
  wire _2368_;
  wire _2369_;
  wire _2370_;
  wire _2371_;
  wire _2372_;
  wire _2373_;
  wire _2374_;
  wire _2375_;
  wire _2376_;
  wire _2377_;
  wire _2378_;
  wire _2379_;
  wire _2380_;
  wire _2381_;
  wire _2382_;
  wire _2383_;
  wire _2384_;
  wire _2385_;
  wire _2386_;
  wire _2387_;
  wire _2388_;
  wire _2389_;
  wire _2390_;
  wire _2391_;
  wire _2392_;
  wire _2393_;
  wire _2394_;
  wire _2395_;
  wire _2396_;
  wire _2397_;
  wire _2398_;
  wire _2399_;
  wire _2400_;
  wire _2401_;
  wire _2402_;
  wire _2403_;
  wire _2404_;
  wire _2405_;
  wire _2406_;
  wire _2407_;
  wire _2408_;
  wire _2409_;
  wire _2410_;
  wire _2411_;
  wire _2412_;
  wire _2413_;
  wire _2414_;
  wire _2415_;
  wire _2416_;
  wire _2417_;
  wire _2418_;
  wire _2419_;
  wire _2420_;
  wire _2421_;
  wire _2422_;
  wire _2423_;
  wire _2424_;
  wire _2425_;
  wire _2426_;
  wire _2427_;
  wire _2428_;
  wire _2429_;
  wire _2430_;
  wire _2431_;
  wire _2432_;
  wire _2433_;
  wire _2434_;
  wire _2435_;
  wire _2436_;
  wire _2437_;
  wire _2438_;
  wire _2439_;
  wire _2440_;
  wire _2441_;
  wire _2442_;
  wire _2443_;
  wire _2444_;
  wire _2445_;
  wire _2446_;
  wire _2447_;
  wire _2448_;
  wire _2449_;
  wire _2450_;
  wire _2451_;
  wire _2452_;
  wire _2453_;
  wire _2454_;
  wire _2455_;
  wire _2456_;
  wire _2457_;
  wire _2458_;
  wire _2459_;
  wire _2460_;
  wire _2461_;
  wire _2462_;
  wire _2463_;
  wire _2464_;
  wire _2465_;
  wire _2466_;
  wire _2467_;
  wire _2468_;
  wire _2469_;
  wire _2470_;
  wire _2471_;
  wire _2472_;
  wire _2473_;
  wire _2474_;
  wire _2475_;
  wire _2476_;
  wire _2477_;
  wire _2478_;
  wire _2479_;
  wire _2480_;
  wire _2481_;
  wire _2482_;
  wire _2483_;
  wire _2484_;
  wire _2485_;
  wire _2486_;
  wire _2487_;
  wire _2488_;
  wire _2489_;
  wire _2490_;
  wire _2491_;
  wire _2492_;
  wire _2493_;
  wire _2494_;
  wire _2495_;
  wire _2496_;
  wire _2497_;
  wire _2498_;
  wire _2499_;
  wire _2500_;
  wire _2501_;
  wire _2502_;
  wire _2503_;
  wire _2504_;
  wire _2505_;
  wire _2506_;
  wire _2507_;
  wire _2508_;
  wire _2509_;
  wire _2510_;
  wire _2511_;
  wire _2512_;
  wire _2513_;
  wire _2514_;
  wire _2515_;
  wire _2516_;
  wire _2517_;
  wire _2518_;
  wire _2519_;
  wire _2520_;
  wire _2521_;
  wire _2522_;
  wire _2523_;
  wire _2524_;
  wire _2525_;
  wire _2526_;
  wire _2527_;
  wire _2528_;
  wire _2529_;
  wire _2530_;
  wire _2531_;
  wire _2532_;
  wire _2533_;
  wire _2534_;
  wire _2535_;
  wire _2536_;
  wire _2537_;
  wire _2538_;
  wire _2539_;
  wire _2540_;
  wire _2541_;
  wire _2542_;
  wire _2543_;
  wire _2544_;
  wire _2545_;
  wire _2546_;
  wire _2547_;
  wire _2548_;
  wire _2549_;
  wire _2550_;
  wire _2551_;
  wire _2552_;
  wire _2553_;
  wire _2554_;
  wire _2555_;
  wire _2556_;
  wire _2557_;
  wire _2558_;
  wire _2559_;
  wire _2560_;
  wire _2561_;
  wire _2562_;
  wire _2563_;
  wire _2564_;
  wire _2565_;
  wire _2566_;
  wire _2567_;
  wire _2568_;
  wire _2569_;
  wire _2570_;
  wire _2571_;
  wire _2572_;
  wire _2573_;
  wire _2574_;
  wire _2575_;
  wire _2576_;
  wire _2577_;
  wire _2578_;
  wire _2579_;
  wire _2580_;
  wire _2581_;
  wire _2582_;
  wire _2583_;
  wire _2584_;
  wire _2585_;
  wire _2586_;
  wire _2587_;
  wire _2588_;
  wire _2589_;
  wire _2590_;
  wire _2591_;
  wire _2592_;
  wire _2593_;
  wire _2594_;
  wire _2595_;
  wire _2596_;
  wire _2597_;
  wire _2598_;
  wire _2599_;
  wire _2600_;
  wire _2601_;
  wire _2602_;
  wire _2603_;
  wire _2604_;
  wire _2605_;
  wire _2606_;
  wire _2607_;
  wire _2608_;
  wire _2609_;
  wire _2610_;
  wire _2611_;
  wire _2612_;
  wire _2613_;
  wire _2614_;
  wire _2615_;
  wire _2616_;
  wire _2617_;
  wire _2618_;
  wire _2619_;
  wire _2620_;
  wire _2621_;
  wire _2622_;
  wire _2623_;
  wire _2624_;
  wire _2625_;
  wire _2626_;
  wire _2627_;
  wire _2628_;
  wire _2629_;
  wire _2630_;
  wire _2631_;
  wire _2632_;
  wire _2633_;
  wire _2634_;
  wire _2635_;
  wire _2636_;
  wire _2637_;
  wire _2638_;
  wire _2639_;
  wire _2640_;
  wire _2641_;
  wire _2642_;
  wire _2643_;
  wire _2644_;
  wire _2645_;
  wire _2646_;
  wire _2647_;
  wire _2648_;
  wire _2649_;
  wire _2650_;
  wire _2651_;
  wire _2652_;
  wire _2653_;
  wire _2654_;
  wire _2655_;
  wire _2656_;
  wire _2657_;
  wire _2658_;
  wire _2659_;
  wire _2660_;
  wire _2661_;
  wire _2662_;
  wire _2663_;
  wire _2664_;
  wire _2665_;
  wire _2666_;
  wire _2667_;
  wire _2668_;
  wire _2669_;
  wire _2670_;
  wire _2671_;
  wire _2672_;
  wire _2673_;
  wire _2674_;
  wire _2675_;
  wire _2676_;
  wire _2677_;
  wire _2678_;
  wire _2679_;
  wire _2680_;
  wire _2681_;
  wire _2682_;
  wire _2683_;
  wire _2684_;
  wire _2685_;
  wire _2686_;
  wire _2687_;
  wire _2688_;
  wire _2689_;
  wire _2690_;
  wire _2691_;
  wire _2692_;
  wire _2693_;
  wire _2694_;
  wire _2695_;
  wire _2696_;
  wire _2697_;
  wire _2698_;
  wire _2699_;
  wire _2700_;
  wire _2701_;
  wire _2702_;
  wire _2703_;
  wire _2704_;
  wire _2705_;
  wire _2706_;
  wire _2707_;
  wire _2708_;
  wire _2709_;
  wire _2710_;
  wire _2711_;
  wire _2712_;
  wire _2713_;
  wire _2714_;
  wire _2715_;
  wire _2716_;
  wire _2717_;
  wire _2718_;
  wire _2719_;
  wire _2720_;
  wire _2721_;
  wire _2722_;
  wire _2723_;
  wire _2724_;
  wire _2725_;
  wire _2726_;
  wire _2727_;
  wire _2728_;
  wire _2729_;
  wire _2730_;
  wire _2731_;
  wire _2732_;
  wire _2733_;
  wire _2734_;
  wire _2735_;
  wire _2736_;
  wire _2737_;
  wire _2738_;
  wire _2739_;
  wire _2740_;
  wire _2741_;
  wire _2742_;
  wire _2743_;
  wire _2744_;
  wire _2745_;
  wire _2746_;
  wire _2747_;
  wire _2748_;
  wire _2749_;
  wire _2750_;
  wire _2751_;
  wire _2752_;
  wire _2753_;
  wire _2754_;
  wire _2755_;
  wire _2756_;
  wire _2757_;
  wire _2758_;
  wire _2759_;
  wire _2760_;
  wire _2761_;
  wire _2762_;
  wire _2763_;
  wire _2764_;
  wire _2765_;
  wire _2766_;
  wire _2767_;
  wire _2768_;
  wire _2769_;
  wire _2770_;
  wire _2771_;
  wire _2772_;
  wire _2773_;
  wire _2774_;
  wire _2775_;
  wire _2776_;
  wire _2777_;
  wire _2778_;
  wire _2779_;
  wire _2780_;
  wire _2781_;
  wire _2782_;
  wire _2783_;
  wire _2784_;
  wire _2785_;
  wire _2786_;
  wire _2787_;
  wire _2788_;
  wire _2789_;
  wire _2790_;
  wire _2791_;
  wire _2792_;
  wire _2793_;
  wire _2794_;
  wire _2795_;
  wire _2796_;
  wire _2797_;
  wire _2798_;
  wire _2799_;
  wire _2800_;
  wire _2801_;
  wire _2802_;
  wire _2803_;
  wire _2804_;
  wire _2805_;
  wire _2806_;
  wire _2807_;
  wire _2808_;
  wire _2809_;
  wire _2810_;
  wire _2811_;
  wire _2812_;
  wire _2813_;
  wire _2814_;
  wire _2815_;
  wire _2816_;
  wire _2817_;
  wire _2818_;
  wire _2819_;
  wire _2820_;
  wire _2821_;
  wire _2822_;
  wire _2823_;
  wire _2824_;
  wire _2825_;
  wire _2826_;
  wire _2827_;
  wire _2828_;
  wire _2829_;
  wire _2830_;
  wire _2831_;
  wire _2832_;
  wire _2833_;
  wire _2834_;
  wire _2835_;
  wire _2836_;
  wire _2837_;
  wire _2838_;
  wire _2839_;
  wire _2840_;
  wire _2841_;
  wire _2842_;
  wire _2843_;
  wire _2844_;
  wire _2845_;
  wire _2846_;
  wire _2847_;
  wire _2848_;
  wire _2849_;
  wire _2850_;
  wire _2851_;
  wire _2852_;
  wire _2853_;
  wire _2854_;
  wire _2855_;
  wire _2856_;
  wire _2857_;
  wire _2858_;
  wire _2859_;
  wire _2860_;
  wire _2861_;
  wire _2862_;
  wire _2863_;
  wire _2864_;
  wire _2865_;
  wire _2866_;
  wire _2867_;
  wire _2868_;
  wire _2869_;
  wire _2870_;
  wire _2871_;
  wire _2872_;
  wire _2873_;
  wire _2874_;
  wire _2875_;
  wire _2876_;
  wire _2877_;
  wire _2878_;
  wire _2879_;
  wire _2880_;
  wire _2881_;
  wire _2882_;
  wire _2883_;
  wire _2884_;
  wire _2885_;
  wire _2886_;
  wire _2887_;
  wire _2888_;
  wire _2889_;
  wire _2890_;
  wire _2891_;
  wire _2892_;
  wire _2893_;
  wire _2894_;
  wire _2895_;
  wire _2896_;
  wire _2897_;
  wire _2898_;
  wire _2899_;
  wire _2900_;
  wire _2901_;
  wire _2902_;
  wire _2903_;
  wire _2904_;
  wire _2905_;
  wire _2906_;
  wire _2907_;
  wire _2908_;
  wire _2909_;
  wire _2910_;
  wire _2911_;
  wire _2912_;
  wire _2913_;
  wire _2914_;
  wire _2915_;
  wire _2916_;
  wire _2917_;
  wire _2918_;
  wire _2919_;
  wire _2920_;
  wire _2921_;
  wire _2922_;
  wire _2923_;
  wire _2924_;
  wire _2925_;
  wire _2926_;
  wire _2927_;
  wire _2928_;
  wire _2929_;
  wire _2930_;
  wire _2931_;
  wire _2932_;
  wire _2933_;
  wire _2934_;
  wire _2935_;
  wire _2936_;
  wire _2937_;
  wire _2938_;
  wire _2939_;
  wire _2940_;
  wire _2941_;
  wire _2942_;
  wire _2943_;
  wire _2944_;
  wire _2945_;
  wire _2946_;
  wire _2947_;
  wire _2948_;
  wire _2949_;
  wire _2950_;
  wire _2951_;
  wire _2952_;
  wire _2953_;
  wire _2954_;
  wire _2955_;
  wire _2956_;
  wire _2957_;
  wire _2958_;
  wire _2959_;
  wire _2960_;
  wire _2961_;
  wire _2962_;
  wire _2963_;
  wire _2964_;
  wire _2965_;
  wire _2966_;
  wire _2967_;
  wire _2968_;
  wire _2969_;
  wire _2970_;
  wire _2971_;
  wire _2972_;
  wire _2973_;
  wire _2974_;
  wire _2975_;
  wire _2976_;
  wire _2977_;
  wire _2978_;
  wire _2979_;
  wire _2980_;
  wire _2981_;
  wire _2982_;
  wire _2983_;
  wire _2984_;
  wire _2985_;
  wire _2986_;
  wire _2987_;
  wire _2988_;
  wire _2989_;
  wire _2990_;
  wire _2991_;
  wire _2992_;
  wire _2993_;
  wire _2994_;
  wire _2995_;
  wire _2996_;
  wire _2997_;
  wire _2998_;
  wire _2999_;
  wire _3000_;
  wire _3001_;
  wire _3002_;
  wire _3003_;
  wire _3004_;
  wire _3005_;
  wire _3006_;
  wire _3007_;
  wire _3008_;
  wire _3009_;
  wire _3010_;
  wire _3011_;
  wire _3012_;
  wire _3013_;
  wire _3014_;
  wire _3015_;
  wire _3016_;
  wire _3017_;
  wire _3018_;
  wire _3019_;
  wire _3020_;
  wire _3021_;
  wire _3022_;
  wire _3023_;
  wire _3024_;
  wire _3025_;
  wire _3026_;
  wire _3027_;
  wire _3028_;
  wire _3029_;
  wire _3030_;
  wire _3031_;
  wire _3032_;
  wire _3033_;
  wire _3034_;
  wire _3035_;
  wire _3036_;
  wire _3037_;
  wire _3038_;
  wire _3039_;
  wire _3040_;
  wire _3041_;
  wire _3042_;
  wire _3043_;
  wire _3044_;
  wire _3045_;
  wire _3046_;
  wire _3047_;
  wire _3048_;
  wire _3049_;
  wire _3050_;
  wire _3051_;
  wire _3052_;
  wire _3053_;
  wire _3054_;
  wire _3055_;
  wire _3056_;
  wire _3057_;
  wire _3058_;
  wire _3059_;
  wire _3060_;
  wire _3061_;
  wire _3062_;
  wire _3063_;
  wire _3064_;
  wire _3065_;
  wire _3066_;
  wire _3067_;
  wire _3068_;
  wire _3069_;
  wire _3070_;
  wire _3071_;
  wire _3072_;
  wire _3073_;
  wire _3074_;
  wire _3075_;
  wire _3076_;
  wire _3077_;
  wire _3078_;
  wire _3079_;
  wire _3080_;
  wire _3081_;
  wire _3082_;
  wire _3083_;
  wire _3084_;
  wire _3085_;
  wire _3086_;
  wire _3087_;
  wire _3088_;
  wire _3089_;
  wire _3090_;
  wire _3091_;
  wire _3092_;
  wire _3093_;
  wire _3094_;
  wire _3095_;
  wire _3096_;
  wire _3097_;
  wire _3098_;
  wire _3099_;
  wire _3100_;
  wire _3101_;
  wire _3102_;
  wire _3103_;
  wire _3104_;
  wire _3105_;
  wire _3106_;
  wire _3107_;
  wire _3108_;
  wire _3109_;
  wire _3110_;
  wire _3111_;
  wire _3112_;
  wire _3113_;
  wire _3114_;
  wire _3115_;
  wire _3116_;
  wire _3117_;
  wire _3118_;
  wire _3119_;
  wire _3120_;
  wire _3121_;
  wire _3122_;
  wire _3123_;
  wire _3124_;
  wire _3125_;
  wire _3126_;
  wire _3127_;
  wire _3128_;
  wire _3129_;
  wire _3130_;
  wire _3131_;
  wire _3132_;
  wire _3133_;
  wire _3134_;
  wire _3135_;
  wire _3136_;
  wire _3137_;
  wire _3138_;
  wire _3139_;
  wire _3140_;
  wire _3141_;
  wire _3142_;
  wire _3143_;
  wire _3144_;
  wire _3145_;
  wire _3146_;
  wire _3147_;
  wire _3148_;
  wire _3149_;
  wire _3150_;
  wire _3151_;
  wire _3152_;
  wire _3153_;
  wire _3154_;
  wire _3155_;
  wire _3156_;
  wire _3157_;
  wire _3158_;
  wire _3159_;
  wire _3160_;
  wire _3161_;
  wire _3162_;
  wire _3163_;
  wire _3164_;
  wire _3165_;
  wire _3166_;
  wire _3167_;
  wire _3168_;
  wire _3169_;
  wire _3170_;
  wire _3171_;
  wire _3172_;
  wire _3173_;
  wire _3174_;
  wire _3175_;
  wire _3176_;
  wire _3177_;
  wire _3178_;
  wire _3179_;
  wire _3180_;
  wire _3181_;
  wire _3182_;
  wire _3183_;
  wire _3184_;
  wire _3185_;
  wire _3186_;
  wire _3187_;
  wire _3188_;
  wire _3189_;
  wire _3190_;
  wire _3191_;
  wire _3192_;
  wire _3193_;
  wire _3194_;
  wire _3195_;
  wire _3196_;
  wire _3197_;
  wire _3198_;
  wire _3199_;
  wire _3200_;
  wire _3201_;
  wire _3202_;
  wire _3203_;
  wire _3204_;
  wire _3205_;
  wire _3206_;
  wire _3207_;
  wire _3208_;
  wire _3209_;
  wire _3210_;
  wire _3211_;
  wire _3212_;
  wire _3213_;
  wire _3214_;
  wire _3215_;
  wire _3216_;
  wire _3217_;
  wire _3218_;
  wire _3219_;
  wire _3220_;
  wire _3221_;
  wire _3222_;
  wire _3223_;
  wire _3224_;
  wire _3225_;
  wire _3226_;
  wire _3227_;
  wire _3228_;
  wire _3229_;
  wire _3230_;
  wire _3231_;
  wire _3232_;
  wire _3233_;
  wire _3234_;
  wire _3235_;
  wire _3236_;
  wire _3237_;
  wire _3238_;
  wire _3239_;
  wire _3240_;
  wire _3241_;
  wire _3242_;
  wire _3243_;
  wire _3244_;
  wire _3245_;
  wire _3246_;
  wire _3247_;
  wire _3248_;
  wire _3249_;
  wire _3250_;
  wire _3251_;
  wire _3252_;
  wire _3253_;
  wire _3254_;
  wire _3255_;
  wire _3256_;
  wire _3257_;
  wire _3258_;
  wire _3259_;
  wire _3260_;
  wire _3261_;
  wire _3262_;
  wire _3263_;
  wire _3264_;
  wire _3265_;
  wire _3266_;
  wire _3267_;
  wire _3268_;
  wire _3269_;
  wire _3270_;
  wire _3271_;
  wire _3272_;
  wire _3273_;
  wire _3274_;
  wire _3275_;
  wire _3276_;
  wire _3277_;
  wire _3278_;
  wire _3279_;
  wire _3280_;
  wire _3281_;
  wire _3282_;
  wire _3283_;
  wire _3284_;
  wire _3285_;
  wire _3286_;
  wire _3287_;
  wire _3288_;
  wire _3289_;
  wire _3290_;
  wire _3291_;
  wire _3292_;
  wire _3293_;
  wire _3294_;
  wire _3295_;
  wire _3296_;
  wire _3297_;
  wire _3298_;
  wire _3299_;
  wire _3300_;
  wire _3301_;
  wire _3302_;
  wire _3303_;
  wire _3304_;
  wire _3305_;
  wire _3306_;
  wire _3307_;
  wire _3308_;
  wire _3309_;
  wire _3310_;
  wire _3311_;
  wire _3312_;
  wire _3313_;
  wire _3314_;
  wire _3315_;
  wire _3316_;
  wire _3317_;
  wire _3318_;
  wire _3319_;
  wire _3320_;
  wire _3321_;
  wire _3322_;
  wire _3323_;
  wire _3324_;
  wire _3325_;
  wire _3326_;
  wire _3327_;
  wire _3328_;
  wire _3329_;
  wire _3330_;
  wire _3331_;
  wire _3332_;
  wire _3333_;
  wire _3334_;
  wire _3335_;
  wire _3336_;
  wire _3337_;
  wire _3338_;
  wire _3339_;
  wire _3340_;
  wire _3341_;
  wire _3342_;
  wire _3343_;
  wire _3344_;
  wire _3345_;
  wire _3346_;
  wire _3347_;
  wire _3348_;
  wire _3349_;
  wire _3350_;
  wire _3351_;
  wire _3352_;
  wire _3353_;
  wire _3354_;
  wire _3355_;
  wire _3356_;
  wire _3357_;
  wire _3358_;
  wire _3359_;
  wire _3360_;
  wire _3361_;
  wire _3362_;
  wire _3363_;
  wire _3364_;
  wire _3365_;
  wire _3366_;
  wire _3367_;
  wire _3368_;
  wire _3369_;
  wire _3370_;
  wire _3371_;
  wire _3372_;
  wire _3373_;
  wire _3374_;
  wire _3375_;
  wire _3376_;
  wire _3377_;
  wire _3378_;
  wire _3379_;
  wire _3380_;
  wire _3381_;
  wire _3382_;
  wire _3383_;
  wire _3384_;
  wire _3385_;
  wire _3386_;
  wire _3387_;
  wire _3388_;
  wire _3389_;
  wire _3390_;
  wire _3391_;
  wire _3392_;
  wire _3393_;
  wire _3394_;
  wire _3395_;
  wire _3396_;
  wire _3397_;
  wire _3398_;
  wire _3399_;
  wire _3400_;
  wire _3401_;
  wire _3402_;
  wire _3403_;
  wire _3404_;
  wire _3405_;
  wire _3406_;
  wire _3407_;
  wire _3408_;
  wire _3409_;
  wire _3410_;
  wire _3411_;
  wire _3412_;
  wire _3413_;
  wire _3414_;
  wire _3415_;
  wire _3416_;
  wire _3417_;
  wire _3418_;
  wire _3419_;
  wire _3420_;
  wire _3421_;
  wire _3422_;
  wire _3423_;
  wire _3424_;
  wire _3425_;
  wire _3426_;
  wire _3427_;
  wire _3428_;
  wire _3429_;
  wire _3430_;
  wire _3431_;
  wire _3432_;
  wire _3433_;
  wire _3434_;
  wire _3435_;
  wire _3436_;
  wire _3437_;
  wire _3438_;
  wire _3439_;
  wire _3440_;
  wire _3441_;
  wire _3442_;
  wire _3443_;
  wire _3444_;
  wire _3445_;
  wire _3446_;
  wire _3447_;
  wire _3448_;
  wire _3449_;
  wire _3450_;
  wire _3451_;
  wire _3452_;
  wire _3453_;
  wire _3454_;
  wire _3455_;
  wire _3456_;
  wire _3457_;
  wire _3458_;
  wire _3459_;
  wire _3460_;
  wire _3461_;
  wire _3462_;
  wire _3463_;
  wire _3464_;
  wire _3465_;
  wire _3466_;
  wire _3467_;
  wire _3468_;
  wire _3469_;
  wire _3470_;
  wire _3471_;
  wire _3472_;
  wire _3473_;
  wire _3474_;
  wire _3475_;
  wire _3476_;
  wire _3477_;
  wire _3478_;
  wire _3479_;
  wire _3480_;
  wire _3481_;
  wire _3482_;
  wire _3483_;
  wire _3484_;
  wire _3485_;
  wire _3486_;
  wire _3487_;
  wire _3488_;
  wire _3489_;
  wire _3490_;
  wire _3491_;
  wire _3492_;
  wire _3493_;
  wire _3494_;
  wire _3495_;
  wire _3496_;
  wire _3497_;
  wire _3498_;
  wire _3499_;
  wire _3500_;
  wire _3501_;
  wire _3502_;
  wire _3503_;
  wire _3504_;
  wire _3505_;
  wire _3506_;
  wire _3507_;
  wire _3508_;
  wire _3509_;
  wire _3510_;
  wire _3511_;
  wire _3512_;
  wire _3513_;
  wire _3514_;
  wire _3515_;
  wire _3516_;
  wire _3517_;
  wire _3518_;
  wire _3519_;
  wire _3520_;
  wire _3521_;
  wire _3522_;
  wire _3523_;
  wire _3524_;
  wire _3525_;
  wire _3526_;
  wire _3527_;
  wire _3528_;
  wire _3529_;
  wire _3530_;
  wire _3531_;
  wire _3532_;
  wire _3533_;
  wire _3534_;
  wire _3535_;
  wire _3536_;
  wire _3537_;
  wire _3538_;
  wire _3539_;
  wire _3540_;
  wire _3541_;
  wire _3542_;
  wire _3543_;
  wire _3544_;
  wire _3545_;
  wire _3546_;
  wire _3547_;
  wire _3548_;
  wire _3549_;
  wire _3550_;
  wire _3551_;
  wire _3552_;
  wire _3553_;
  wire _3554_;
  wire _3555_;
  wire _3556_;
  wire _3557_;
  wire _3558_;
  wire _3559_;
  wire _3560_;
  wire _3561_;
  wire _3562_;
  wire _3563_;
  wire _3564_;
  wire _3565_;
  wire _3566_;
  wire _3567_;
  wire _3568_;
  wire _3569_;
  wire _3570_;
  wire _3571_;
  wire _3572_;
  wire _3573_;
  wire _3574_;
  wire _3575_;
  wire _3576_;
  wire _3577_;
  wire _3578_;
  wire _3579_;
  wire _3580_;
  wire _3581_;
  wire _3582_;
  wire _3583_;
  wire _3584_;
  wire _3585_;
  wire _3586_;
  wire _3587_;
  wire _3588_;
  wire _3589_;
  wire _3590_;
  wire _3591_;
  input CK;
  wire \DFF_0.CK ;
  wire \DFF_0.D ;
  wire \DFF_0.Q ;
  wire \DFF_1.CK ;
  wire \DFF_1.D ;
  wire \DFF_1.Q ;
  wire \DFF_10.CK ;
  wire \DFF_10.D ;
  wire \DFF_10.Q ;
  wire \DFF_100.CK ;
  wire \DFF_100.D ;
  wire \DFF_100.Q ;
  wire \DFF_1000.CK ;
  wire \DFF_1000.D ;
  wire \DFF_1000.Q ;
  wire \DFF_1001.CK ;
  wire \DFF_1001.D ;
  wire \DFF_1001.Q ;
  wire \DFF_1002.CK ;
  wire \DFF_1002.D ;
  wire \DFF_1002.Q ;
  wire \DFF_1003.CK ;
  wire \DFF_1003.D ;
  wire \DFF_1003.Q ;
  wire \DFF_1004.CK ;
  wire \DFF_1004.D ;
  wire \DFF_1004.Q ;
  wire \DFF_1005.CK ;
  wire \DFF_1005.D ;
  wire \DFF_1005.Q ;
  wire \DFF_1006.CK ;
  wire \DFF_1006.D ;
  wire \DFF_1006.Q ;
  wire \DFF_1007.CK ;
  wire \DFF_1007.D ;
  wire \DFF_1007.Q ;
  wire \DFF_1008.CK ;
  wire \DFF_1008.D ;
  wire \DFF_1008.Q ;
  wire \DFF_1009.CK ;
  wire \DFF_1009.D ;
  wire \DFF_1009.Q ;
  wire \DFF_101.CK ;
  wire \DFF_101.D ;
  wire \DFF_101.Q ;
  wire \DFF_1010.CK ;
  wire \DFF_1010.D ;
  wire \DFF_1010.Q ;
  wire \DFF_1011.CK ;
  wire \DFF_1011.D ;
  wire \DFF_1011.Q ;
  wire \DFF_1012.CK ;
  wire \DFF_1012.D ;
  wire \DFF_1012.Q ;
  wire \DFF_1013.CK ;
  wire \DFF_1013.D ;
  wire \DFF_1013.Q ;
  wire \DFF_1014.CK ;
  wire \DFF_1014.D ;
  wire \DFF_1014.Q ;
  wire \DFF_1015.CK ;
  wire \DFF_1015.D ;
  wire \DFF_1015.Q ;
  wire \DFF_1016.CK ;
  wire \DFF_1016.D ;
  wire \DFF_1016.Q ;
  wire \DFF_1017.CK ;
  wire \DFF_1017.D ;
  wire \DFF_1017.Q ;
  wire \DFF_1018.CK ;
  wire \DFF_1019.CK ;
  wire \DFF_102.CK ;
  wire \DFF_102.D ;
  wire \DFF_102.Q ;
  wire \DFF_1020.CK ;
  wire \DFF_1021.CK ;
  wire \DFF_1022.CK ;
  wire \DFF_1023.CK ;
  wire \DFF_1024.CK ;
  wire \DFF_1025.CK ;
  wire \DFF_1026.CK ;
  wire \DFF_1027.CK ;
  wire \DFF_1028.CK ;
  wire \DFF_1028.D ;
  wire \DFF_1028.Q ;
  wire \DFF_1029.CK ;
  wire \DFF_1029.D ;
  wire \DFF_1029.Q ;
  wire \DFF_103.CK ;
  wire \DFF_103.D ;
  wire \DFF_103.Q ;
  wire \DFF_1030.CK ;
  wire \DFF_1030.D ;
  wire \DFF_1030.Q ;
  wire \DFF_1031.CK ;
  wire \DFF_1031.D ;
  wire \DFF_1031.Q ;
  wire \DFF_1032.CK ;
  wire \DFF_1032.D ;
  wire \DFF_1032.Q ;
  wire \DFF_1033.CK ;
  wire \DFF_1033.D ;
  wire \DFF_1033.Q ;
  wire \DFF_1034.CK ;
  wire \DFF_1034.D ;
  wire \DFF_1034.Q ;
  wire \DFF_1035.CK ;
  wire \DFF_1035.D ;
  wire \DFF_1035.Q ;
  wire \DFF_1036.CK ;
  wire \DFF_1036.D ;
  wire \DFF_1036.Q ;
  wire \DFF_1037.CK ;
  wire \DFF_1037.D ;
  wire \DFF_1037.Q ;
  wire \DFF_1038.CK ;
  wire \DFF_1038.D ;
  wire \DFF_1038.Q ;
  wire \DFF_1039.CK ;
  wire \DFF_1039.D ;
  wire \DFF_1039.Q ;
  wire \DFF_104.CK ;
  wire \DFF_104.D ;
  wire \DFF_104.Q ;
  wire \DFF_1040.CK ;
  wire \DFF_1040.D ;
  wire \DFF_1040.Q ;
  wire \DFF_1041.CK ;
  wire \DFF_1041.D ;
  wire \DFF_1041.Q ;
  wire \DFF_1042.CK ;
  wire \DFF_1042.D ;
  wire \DFF_1042.Q ;
  wire \DFF_1043.CK ;
  wire \DFF_1043.D ;
  wire \DFF_1043.Q ;
  wire \DFF_1044.CK ;
  wire \DFF_1044.D ;
  wire \DFF_1044.Q ;
  wire \DFF_1045.CK ;
  wire \DFF_1045.D ;
  wire \DFF_1045.Q ;
  wire \DFF_1046.CK ;
  wire \DFF_1046.D ;
  wire \DFF_1046.Q ;
  wire \DFF_1047.CK ;
  wire \DFF_1047.D ;
  wire \DFF_1047.Q ;
  wire \DFF_1048.CK ;
  wire \DFF_1048.D ;
  wire \DFF_1048.Q ;
  wire \DFF_1049.CK ;
  wire \DFF_1049.D ;
  wire \DFF_1049.Q ;
  wire \DFF_105.CK ;
  wire \DFF_105.D ;
  wire \DFF_105.Q ;
  wire \DFF_1050.CK ;
  wire \DFF_1050.D ;
  wire \DFF_1050.Q ;
  wire \DFF_1051.CK ;
  wire \DFF_1051.D ;
  wire \DFF_1051.Q ;
  wire \DFF_1052.CK ;
  wire \DFF_1052.D ;
  wire \DFF_1052.Q ;
  wire \DFF_1053.CK ;
  wire \DFF_1053.D ;
  wire \DFF_1053.Q ;
  wire \DFF_1054.CK ;
  wire \DFF_1054.D ;
  wire \DFF_1054.Q ;
  wire \DFF_1055.CK ;
  wire \DFF_1055.D ;
  wire \DFF_1055.Q ;
  wire \DFF_1056.CK ;
  wire \DFF_1056.D ;
  wire \DFF_1056.Q ;
  wire \DFF_1057.CK ;
  wire \DFF_1057.D ;
  wire \DFF_1057.Q ;
  wire \DFF_1058.CK ;
  wire \DFF_1058.D ;
  wire \DFF_1058.Q ;
  wire \DFF_1059.CK ;
  wire \DFF_1059.D ;
  wire \DFF_1059.Q ;
  wire \DFF_106.CK ;
  wire \DFF_106.D ;
  wire \DFF_106.Q ;
  wire \DFF_1060.CK ;
  wire \DFF_1060.D ;
  wire \DFF_1060.Q ;
  wire \DFF_1061.CK ;
  wire \DFF_1061.D ;
  wire \DFF_1061.Q ;
  wire \DFF_1062.CK ;
  wire \DFF_1062.D ;
  wire \DFF_1062.Q ;
  wire \DFF_1063.CK ;
  wire \DFF_1063.D ;
  wire \DFF_1063.Q ;
  wire \DFF_1064.CK ;
  wire \DFF_1064.D ;
  wire \DFF_1064.Q ;
  wire \DFF_1065.CK ;
  wire \DFF_1065.D ;
  wire \DFF_1065.Q ;
  wire \DFF_1066.CK ;
  wire \DFF_1066.D ;
  wire \DFF_1066.Q ;
  wire \DFF_1067.CK ;
  wire \DFF_1067.D ;
  wire \DFF_1067.Q ;
  wire \DFF_1068.CK ;
  wire \DFF_1068.D ;
  wire \DFF_1068.Q ;
  wire \DFF_1069.CK ;
  wire \DFF_1069.D ;
  wire \DFF_1069.Q ;
  wire \DFF_107.CK ;
  wire \DFF_107.D ;
  wire \DFF_107.Q ;
  wire \DFF_1070.CK ;
  wire \DFF_1070.D ;
  wire \DFF_1070.Q ;
  wire \DFF_1071.CK ;
  wire \DFF_1071.D ;
  wire \DFF_1071.Q ;
  wire \DFF_1072.CK ;
  wire \DFF_1072.D ;
  wire \DFF_1072.Q ;
  wire \DFF_1073.CK ;
  wire \DFF_1073.D ;
  wire \DFF_1073.Q ;
  wire \DFF_1074.CK ;
  wire \DFF_1074.D ;
  wire \DFF_1074.Q ;
  wire \DFF_1075.CK ;
  wire \DFF_1075.D ;
  wire \DFF_1075.Q ;
  wire \DFF_1076.CK ;
  wire \DFF_1076.D ;
  wire \DFF_1076.Q ;
  wire \DFF_1077.CK ;
  wire \DFF_1077.D ;
  wire \DFF_1077.Q ;
  wire \DFF_1078.CK ;
  wire \DFF_1078.D ;
  wire \DFF_1078.Q ;
  wire \DFF_1079.CK ;
  wire \DFF_1079.D ;
  wire \DFF_1079.Q ;
  wire \DFF_108.CK ;
  wire \DFF_108.D ;
  wire \DFF_108.Q ;
  wire \DFF_1080.CK ;
  wire \DFF_1080.D ;
  wire \DFF_1080.Q ;
  wire \DFF_1081.CK ;
  wire \DFF_1081.D ;
  wire \DFF_1081.Q ;
  wire \DFF_1082.CK ;
  wire \DFF_1082.D ;
  wire \DFF_1082.Q ;
  wire \DFF_1083.CK ;
  wire \DFF_1083.D ;
  wire \DFF_1083.Q ;
  wire \DFF_1084.CK ;
  wire \DFF_1084.D ;
  wire \DFF_1084.Q ;
  wire \DFF_1085.CK ;
  wire \DFF_1085.D ;
  wire \DFF_1085.Q ;
  wire \DFF_1086.CK ;
  wire \DFF_1086.D ;
  wire \DFF_1086.Q ;
  wire \DFF_1087.CK ;
  wire \DFF_1087.D ;
  wire \DFF_1087.Q ;
  wire \DFF_1088.CK ;
  wire \DFF_1088.D ;
  wire \DFF_1088.Q ;
  wire \DFF_1089.CK ;
  wire \DFF_1089.D ;
  wire \DFF_1089.Q ;
  wire \DFF_109.CK ;
  wire \DFF_109.D ;
  wire \DFF_109.Q ;
  wire \DFF_1090.CK ;
  wire \DFF_1090.D ;
  wire \DFF_1090.Q ;
  wire \DFF_1091.CK ;
  wire \DFF_1091.D ;
  wire \DFF_1091.Q ;
  wire \DFF_1092.CK ;
  wire \DFF_1092.D ;
  wire \DFF_1092.Q ;
  wire \DFF_1093.CK ;
  wire \DFF_1093.D ;
  wire \DFF_1093.Q ;
  wire \DFF_1094.CK ;
  wire \DFF_1094.D ;
  wire \DFF_1094.Q ;
  wire \DFF_1095.CK ;
  wire \DFF_1095.D ;
  wire \DFF_1095.Q ;
  wire \DFF_1096.CK ;
  wire \DFF_1096.D ;
  wire \DFF_1096.Q ;
  wire \DFF_1097.CK ;
  wire \DFF_1097.D ;
  wire \DFF_1097.Q ;
  wire \DFF_1098.CK ;
  wire \DFF_1098.D ;
  wire \DFF_1098.Q ;
  wire \DFF_1099.CK ;
  wire \DFF_1099.D ;
  wire \DFF_1099.Q ;
  wire \DFF_11.CK ;
  wire \DFF_11.D ;
  wire \DFF_11.Q ;
  wire \DFF_110.CK ;
  wire \DFF_110.D ;
  wire \DFF_110.Q ;
  wire \DFF_1100.CK ;
  wire \DFF_1100.D ;
  wire \DFF_1100.Q ;
  wire \DFF_1101.CK ;
  wire \DFF_1101.D ;
  wire \DFF_1101.Q ;
  wire \DFF_1102.CK ;
  wire \DFF_1102.D ;
  wire \DFF_1102.Q ;
  wire \DFF_1103.CK ;
  wire \DFF_1103.D ;
  wire \DFF_1103.Q ;
  wire \DFF_1104.CK ;
  wire \DFF_1104.D ;
  wire \DFF_1104.Q ;
  wire \DFF_1105.CK ;
  wire \DFF_1105.D ;
  wire \DFF_1105.Q ;
  wire \DFF_1106.CK ;
  wire \DFF_1106.D ;
  wire \DFF_1106.Q ;
  wire \DFF_1107.CK ;
  wire \DFF_1107.D ;
  wire \DFF_1107.Q ;
  wire \DFF_1108.CK ;
  wire \DFF_1108.D ;
  wire \DFF_1108.Q ;
  wire \DFF_1109.CK ;
  wire \DFF_1109.D ;
  wire \DFF_1109.Q ;
  wire \DFF_111.CK ;
  wire \DFF_111.D ;
  wire \DFF_111.Q ;
  wire \DFF_1110.CK ;
  wire \DFF_1110.D ;
  wire \DFF_1110.Q ;
  wire \DFF_1111.CK ;
  wire \DFF_1111.D ;
  wire \DFF_1111.Q ;
  wire \DFF_1112.CK ;
  wire \DFF_1112.D ;
  wire \DFF_1112.Q ;
  wire \DFF_1113.CK ;
  wire \DFF_1113.D ;
  wire \DFF_1113.Q ;
  wire \DFF_1114.CK ;
  wire \DFF_1114.D ;
  wire \DFF_1114.Q ;
  wire \DFF_1115.CK ;
  wire \DFF_1115.D ;
  wire \DFF_1115.Q ;
  wire \DFF_1116.CK ;
  wire \DFF_1116.D ;
  wire \DFF_1116.Q ;
  wire \DFF_1117.CK ;
  wire \DFF_1117.D ;
  wire \DFF_1117.Q ;
  wire \DFF_1118.CK ;
  wire \DFF_1118.D ;
  wire \DFF_1118.Q ;
  wire \DFF_1119.CK ;
  wire \DFF_1119.D ;
  wire \DFF_1119.Q ;
  wire \DFF_112.CK ;
  wire \DFF_112.D ;
  wire \DFF_112.Q ;
  wire \DFF_1120.CK ;
  wire \DFF_1120.D ;
  wire \DFF_1120.Q ;
  wire \DFF_1121.CK ;
  wire \DFF_1121.D ;
  wire \DFF_1121.Q ;
  wire \DFF_1122.CK ;
  wire \DFF_1122.D ;
  wire \DFF_1122.Q ;
  wire \DFF_1123.CK ;
  wire \DFF_1123.D ;
  wire \DFF_1123.Q ;
  wire \DFF_1124.CK ;
  wire \DFF_1124.D ;
  wire \DFF_1124.Q ;
  wire \DFF_1125.CK ;
  wire \DFF_1125.D ;
  wire \DFF_1125.Q ;
  wire \DFF_1126.CK ;
  wire \DFF_1126.D ;
  wire \DFF_1126.Q ;
  wire \DFF_1127.CK ;
  wire \DFF_1127.D ;
  wire \DFF_1127.Q ;
  wire \DFF_1128.CK ;
  wire \DFF_1128.D ;
  wire \DFF_1128.Q ;
  wire \DFF_1129.CK ;
  wire \DFF_1129.D ;
  wire \DFF_1129.Q ;
  wire \DFF_113.CK ;
  wire \DFF_113.D ;
  wire \DFF_113.Q ;
  wire \DFF_1130.CK ;
  wire \DFF_1130.D ;
  wire \DFF_1130.Q ;
  wire \DFF_1131.CK ;
  wire \DFF_1131.D ;
  wire \DFF_1131.Q ;
  wire \DFF_1132.CK ;
  wire \DFF_1132.D ;
  wire \DFF_1132.Q ;
  wire \DFF_1133.CK ;
  wire \DFF_1133.D ;
  wire \DFF_1133.Q ;
  wire \DFF_1134.CK ;
  wire \DFF_1135.CK ;
  wire \DFF_1136.CK ;
  wire \DFF_1137.CK ;
  wire \DFF_1138.CK ;
  wire \DFF_1139.CK ;
  wire \DFF_114.CK ;
  wire \DFF_114.D ;
  wire \DFF_114.Q ;
  wire \DFF_1140.CK ;
  wire \DFF_1141.CK ;
  wire \DFF_1142.CK ;
  wire \DFF_1142.D ;
  wire \DFF_1142.Q ;
  wire \DFF_1143.CK ;
  wire \DFF_1143.D ;
  wire \DFF_1143.Q ;
  wire \DFF_1144.CK ;
  wire \DFF_1144.D ;
  wire \DFF_1144.Q ;
  wire \DFF_1145.CK ;
  wire \DFF_1145.D ;
  wire \DFF_1145.Q ;
  wire \DFF_1146.CK ;
  wire \DFF_1146.D ;
  wire \DFF_1146.Q ;
  wire \DFF_1147.CK ;
  wire \DFF_1147.D ;
  wire \DFF_1147.Q ;
  wire \DFF_1148.CK ;
  wire \DFF_1148.D ;
  wire \DFF_1148.Q ;
  wire \DFF_1149.CK ;
  wire \DFF_1149.D ;
  wire \DFF_1149.Q ;
  wire \DFF_115.CK ;
  wire \DFF_115.D ;
  wire \DFF_115.Q ;
  wire \DFF_1150.CK ;
  wire \DFF_1150.D ;
  wire \DFF_1150.Q ;
  wire \DFF_1151.CK ;
  wire \DFF_1151.D ;
  wire \DFF_1151.Q ;
  wire \DFF_1152.CK ;
  wire \DFF_1152.D ;
  wire \DFF_1152.Q ;
  wire \DFF_1153.CK ;
  wire \DFF_1153.D ;
  wire \DFF_1153.Q ;
  wire \DFF_1154.CK ;
  wire \DFF_1154.D ;
  wire \DFF_1154.Q ;
  wire \DFF_1155.CK ;
  wire \DFF_1155.D ;
  wire \DFF_1155.Q ;
  wire \DFF_1156.CK ;
  wire \DFF_1156.D ;
  wire \DFF_1156.Q ;
  wire \DFF_1157.CK ;
  wire \DFF_1157.D ;
  wire \DFF_1157.Q ;
  wire \DFF_1158.CK ;
  wire \DFF_1158.D ;
  wire \DFF_1158.Q ;
  wire \DFF_1159.CK ;
  wire \DFF_1159.D ;
  wire \DFF_1159.Q ;
  wire \DFF_116.CK ;
  wire \DFF_116.D ;
  wire \DFF_116.Q ;
  wire \DFF_1160.CK ;
  wire \DFF_1160.D ;
  wire \DFF_1160.Q ;
  wire \DFF_1161.CK ;
  wire \DFF_1161.D ;
  wire \DFF_1161.Q ;
  wire \DFF_1162.CK ;
  wire \DFF_1162.D ;
  wire \DFF_1162.Q ;
  wire \DFF_1163.CK ;
  wire \DFF_1163.D ;
  wire \DFF_1163.Q ;
  wire \DFF_1164.CK ;
  wire \DFF_1164.D ;
  wire \DFF_1164.Q ;
  wire \DFF_1165.CK ;
  wire \DFF_1165.D ;
  wire \DFF_1165.Q ;
  wire \DFF_1166.CK ;
  wire \DFF_1166.D ;
  wire \DFF_1166.Q ;
  wire \DFF_1167.CK ;
  wire \DFF_1167.D ;
  wire \DFF_1167.Q ;
  wire \DFF_1168.CK ;
  wire \DFF_1168.D ;
  wire \DFF_1168.Q ;
  wire \DFF_1169.CK ;
  wire \DFF_1169.D ;
  wire \DFF_1169.Q ;
  wire \DFF_117.CK ;
  wire \DFF_117.D ;
  wire \DFF_117.Q ;
  wire \DFF_1170.CK ;
  wire \DFF_1170.D ;
  wire \DFF_1170.Q ;
  wire \DFF_1171.CK ;
  wire \DFF_1171.D ;
  wire \DFF_1171.Q ;
  wire \DFF_1172.CK ;
  wire \DFF_1172.D ;
  wire \DFF_1172.Q ;
  wire \DFF_1173.CK ;
  wire \DFF_1173.D ;
  wire \DFF_1173.Q ;
  wire \DFF_1174.CK ;
  wire \DFF_1174.D ;
  wire \DFF_1174.Q ;
  wire \DFF_1175.CK ;
  wire \DFF_1175.D ;
  wire \DFF_1175.Q ;
  wire \DFF_1176.CK ;
  wire \DFF_1176.D ;
  wire \DFF_1176.Q ;
  wire \DFF_1177.CK ;
  wire \DFF_1177.D ;
  wire \DFF_1177.Q ;
  wire \DFF_1178.CK ;
  wire \DFF_1178.D ;
  wire \DFF_1178.Q ;
  wire \DFF_1179.CK ;
  wire \DFF_1179.D ;
  wire \DFF_1179.Q ;
  wire \DFF_118.CK ;
  wire \DFF_118.D ;
  wire \DFF_118.Q ;
  wire \DFF_1180.CK ;
  wire \DFF_1180.D ;
  wire \DFF_1180.Q ;
  wire \DFF_1181.CK ;
  wire \DFF_1181.D ;
  wire \DFF_1181.Q ;
  wire \DFF_1182.CK ;
  wire \DFF_1182.D ;
  wire \DFF_1182.Q ;
  wire \DFF_1183.CK ;
  wire \DFF_1183.D ;
  wire \DFF_1183.Q ;
  wire \DFF_1184.CK ;
  wire \DFF_1184.D ;
  wire \DFF_1184.Q ;
  wire \DFF_1185.CK ;
  wire \DFF_1185.D ;
  wire \DFF_1185.Q ;
  wire \DFF_1186.CK ;
  wire \DFF_1186.D ;
  wire \DFF_1186.Q ;
  wire \DFF_1187.CK ;
  wire \DFF_1187.D ;
  wire \DFF_1187.Q ;
  wire \DFF_1188.CK ;
  wire \DFF_1188.D ;
  wire \DFF_1188.Q ;
  wire \DFF_1189.CK ;
  wire \DFF_1189.D ;
  wire \DFF_1189.Q ;
  wire \DFF_119.CK ;
  wire \DFF_119.D ;
  wire \DFF_119.Q ;
  wire \DFF_1190.CK ;
  wire \DFF_1190.D ;
  wire \DFF_1190.Q ;
  wire \DFF_1191.CK ;
  wire \DFF_1191.D ;
  wire \DFF_1191.Q ;
  wire \DFF_1192.CK ;
  wire \DFF_1192.D ;
  wire \DFF_1192.Q ;
  wire \DFF_1193.CK ;
  wire \DFF_1193.D ;
  wire \DFF_1193.Q ;
  wire \DFF_1194.CK ;
  wire \DFF_1194.D ;
  wire \DFF_1194.Q ;
  wire \DFF_1195.CK ;
  wire \DFF_1195.D ;
  wire \DFF_1195.Q ;
  wire \DFF_1196.CK ;
  wire \DFF_1196.D ;
  wire \DFF_1196.Q ;
  wire \DFF_1197.CK ;
  wire \DFF_1197.D ;
  wire \DFF_1197.Q ;
  wire \DFF_1198.CK ;
  wire \DFF_1198.D ;
  wire \DFF_1198.Q ;
  wire \DFF_1199.CK ;
  wire \DFF_1199.D ;
  wire \DFF_1199.Q ;
  wire \DFF_12.CK ;
  wire \DFF_12.D ;
  wire \DFF_12.Q ;
  wire \DFF_120.CK ;
  wire \DFF_120.D ;
  wire \DFF_120.Q ;
  wire \DFF_1200.CK ;
  wire \DFF_1200.D ;
  wire \DFF_1200.Q ;
  wire \DFF_1201.CK ;
  wire \DFF_1201.D ;
  wire \DFF_1201.Q ;
  wire \DFF_1202.CK ;
  wire \DFF_1202.D ;
  wire \DFF_1202.Q ;
  wire \DFF_1203.CK ;
  wire \DFF_1203.D ;
  wire \DFF_1203.Q ;
  wire \DFF_1204.CK ;
  wire \DFF_1204.D ;
  wire \DFF_1204.Q ;
  wire \DFF_1205.CK ;
  wire \DFF_1205.D ;
  wire \DFF_1205.Q ;
  wire \DFF_1206.CK ;
  wire \DFF_1206.D ;
  wire \DFF_1206.Q ;
  wire \DFF_1207.CK ;
  wire \DFF_1207.D ;
  wire \DFF_1207.Q ;
  wire \DFF_1208.CK ;
  wire \DFF_1208.D ;
  wire \DFF_1208.Q ;
  wire \DFF_1209.CK ;
  wire \DFF_1209.D ;
  wire \DFF_1209.Q ;
  wire \DFF_121.CK ;
  wire \DFF_121.D ;
  wire \DFF_121.Q ;
  wire \DFF_1210.CK ;
  wire \DFF_1210.D ;
  wire \DFF_1210.Q ;
  wire \DFF_1211.CK ;
  wire \DFF_1211.D ;
  wire \DFF_1211.Q ;
  wire \DFF_1212.CK ;
  wire \DFF_1212.D ;
  wire \DFF_1212.Q ;
  wire \DFF_1213.CK ;
  wire \DFF_1213.D ;
  wire \DFF_1213.Q ;
  wire \DFF_1214.CK ;
  wire \DFF_1214.D ;
  wire \DFF_1214.Q ;
  wire \DFF_1215.CK ;
  wire \DFF_1215.D ;
  wire \DFF_1215.Q ;
  wire \DFF_1216.CK ;
  wire \DFF_1216.D ;
  wire \DFF_1216.Q ;
  wire \DFF_1217.CK ;
  wire \DFF_1217.D ;
  wire \DFF_1217.Q ;
  wire \DFF_1218.CK ;
  wire \DFF_1218.D ;
  wire \DFF_1218.Q ;
  wire \DFF_1219.CK ;
  wire \DFF_1219.D ;
  wire \DFF_1219.Q ;
  wire \DFF_122.CK ;
  wire \DFF_122.D ;
  wire \DFF_122.Q ;
  wire \DFF_1220.CK ;
  wire \DFF_1220.D ;
  wire \DFF_1220.Q ;
  wire \DFF_1221.CK ;
  wire \DFF_1221.D ;
  wire \DFF_1221.Q ;
  wire \DFF_1222.CK ;
  wire \DFF_1222.D ;
  wire \DFF_1222.Q ;
  wire \DFF_1223.CK ;
  wire \DFF_1223.D ;
  wire \DFF_1223.Q ;
  wire \DFF_1224.CK ;
  wire \DFF_1224.D ;
  wire \DFF_1224.Q ;
  wire \DFF_1225.CK ;
  wire \DFF_1225.D ;
  wire \DFF_1225.Q ;
  wire \DFF_1226.CK ;
  wire \DFF_1226.D ;
  wire \DFF_1226.Q ;
  wire \DFF_1227.CK ;
  wire \DFF_1227.D ;
  wire \DFF_1227.Q ;
  wire \DFF_1228.CK ;
  wire \DFF_1228.D ;
  wire \DFF_1228.Q ;
  wire \DFF_1229.CK ;
  wire \DFF_1229.D ;
  wire \DFF_1229.Q ;
  wire \DFF_123.CK ;
  wire \DFF_123.D ;
  wire \DFF_123.Q ;
  wire \DFF_1230.CK ;
  wire \DFF_1230.D ;
  wire \DFF_1230.Q ;
  wire \DFF_1231.CK ;
  wire \DFF_1231.D ;
  wire \DFF_1231.Q ;
  wire \DFF_1232.CK ;
  wire \DFF_1232.D ;
  wire \DFF_1232.Q ;
  wire \DFF_1233.CK ;
  wire \DFF_1233.D ;
  wire \DFF_1233.Q ;
  wire \DFF_1234.CK ;
  wire \DFF_1234.D ;
  wire \DFF_1234.Q ;
  wire \DFF_1235.CK ;
  wire \DFF_1235.D ;
  wire \DFF_1235.Q ;
  wire \DFF_1236.CK ;
  wire \DFF_1236.D ;
  wire \DFF_1236.Q ;
  wire \DFF_1237.CK ;
  wire \DFF_1237.D ;
  wire \DFF_1237.Q ;
  wire \DFF_1238.CK ;
  wire \DFF_1238.D ;
  wire \DFF_1238.Q ;
  wire \DFF_1239.CK ;
  wire \DFF_1239.D ;
  wire \DFF_1239.Q ;
  wire \DFF_124.CK ;
  wire \DFF_124.D ;
  wire \DFF_124.Q ;
  wire \DFF_1240.CK ;
  wire \DFF_1240.D ;
  wire \DFF_1240.Q ;
  wire \DFF_1241.CK ;
  wire \DFF_1241.D ;
  wire \DFF_1241.Q ;
  wire \DFF_1242.CK ;
  wire \DFF_1242.D ;
  wire \DFF_1242.Q ;
  wire \DFF_1243.CK ;
  wire \DFF_1243.D ;
  wire \DFF_1243.Q ;
  wire \DFF_1244.CK ;
  wire \DFF_1244.D ;
  wire \DFF_1244.Q ;
  wire \DFF_1245.CK ;
  wire \DFF_1245.D ;
  wire \DFF_1245.Q ;
  wire \DFF_1246.CK ;
  wire \DFF_1246.D ;
  wire \DFF_1246.Q ;
  wire \DFF_1247.CK ;
  wire \DFF_1247.D ;
  wire \DFF_1247.Q ;
  wire \DFF_1248.CK ;
  wire \DFF_1248.D ;
  wire \DFF_1248.Q ;
  wire \DFF_1249.CK ;
  wire \DFF_1249.D ;
  wire \DFF_1249.Q ;
  wire \DFF_125.CK ;
  wire \DFF_125.D ;
  wire \DFF_125.Q ;
  wire \DFF_1250.CK ;
  wire \DFF_1250.D ;
  wire \DFF_1250.Q ;
  wire \DFF_1251.CK ;
  wire \DFF_1251.D ;
  wire \DFF_1251.Q ;
  wire \DFF_1252.CK ;
  wire \DFF_1252.D ;
  wire \DFF_1252.Q ;
  wire \DFF_1253.CK ;
  wire \DFF_1253.D ;
  wire \DFF_1253.Q ;
  wire \DFF_1254.CK ;
  wire \DFF_1254.D ;
  wire \DFF_1254.Q ;
  wire \DFF_1255.CK ;
  wire \DFF_1255.D ;
  wire \DFF_1255.Q ;
  wire \DFF_1256.CK ;
  wire \DFF_1256.D ;
  wire \DFF_1256.Q ;
  wire \DFF_1257.CK ;
  wire \DFF_1257.D ;
  wire \DFF_1257.Q ;
  wire \DFF_1258.CK ;
  wire \DFF_1258.D ;
  wire \DFF_1258.Q ;
  wire \DFF_1259.CK ;
  wire \DFF_1259.D ;
  wire \DFF_1259.Q ;
  wire \DFF_126.CK ;
  wire \DFF_126.D ;
  wire \DFF_126.Q ;
  wire \DFF_1260.CK ;
  wire \DFF_1260.D ;
  wire \DFF_1260.Q ;
  wire \DFF_1261.CK ;
  wire \DFF_1261.D ;
  wire \DFF_1261.Q ;
  wire \DFF_1262.CK ;
  wire \DFF_1262.D ;
  wire \DFF_1262.Q ;
  wire \DFF_1263.CK ;
  wire \DFF_1263.D ;
  wire \DFF_1263.Q ;
  wire \DFF_1264.CK ;
  wire \DFF_1264.D ;
  wire \DFF_1264.Q ;
  wire \DFF_1265.CK ;
  wire \DFF_1265.D ;
  wire \DFF_1265.Q ;
  wire \DFF_1266.CK ;
  wire \DFF_1266.D ;
  wire \DFF_1266.Q ;
  wire \DFF_1267.CK ;
  wire \DFF_1267.D ;
  wire \DFF_1267.Q ;
  wire \DFF_1268.CK ;
  wire \DFF_1268.D ;
  wire \DFF_1268.Q ;
  wire \DFF_1269.CK ;
  wire \DFF_1269.D ;
  wire \DFF_1269.Q ;
  wire \DFF_127.CK ;
  wire \DFF_127.D ;
  wire \DFF_127.Q ;
  wire \DFF_1270.CK ;
  wire \DFF_1270.D ;
  wire \DFF_1270.Q ;
  wire \DFF_1271.CK ;
  wire \DFF_1271.D ;
  wire \DFF_1271.Q ;
  wire \DFF_1272.CK ;
  wire \DFF_1272.D ;
  wire \DFF_1272.Q ;
  wire \DFF_1273.CK ;
  wire \DFF_1273.D ;
  wire \DFF_1273.Q ;
  wire \DFF_1274.CK ;
  wire \DFF_1274.D ;
  wire \DFF_1274.Q ;
  wire \DFF_1275.CK ;
  wire \DFF_1275.D ;
  wire \DFF_1275.Q ;
  wire \DFF_1276.CK ;
  wire \DFF_1276.D ;
  wire \DFF_1276.Q ;
  wire \DFF_1277.CK ;
  wire \DFF_1277.D ;
  wire \DFF_1277.Q ;
  wire \DFF_1278.CK ;
  wire \DFF_1278.D ;
  wire \DFF_1278.Q ;
  wire \DFF_1279.CK ;
  wire \DFF_1279.D ;
  wire \DFF_1279.Q ;
  wire \DFF_128.CK ;
  wire \DFF_128.D ;
  wire \DFF_128.Q ;
  wire \DFF_1280.CK ;
  wire \DFF_1280.D ;
  wire \DFF_1280.Q ;
  wire \DFF_1281.CK ;
  wire \DFF_1281.D ;
  wire \DFF_1281.Q ;
  wire \DFF_1282.CK ;
  wire \DFF_1282.D ;
  wire \DFF_1282.Q ;
  wire \DFF_1283.CK ;
  wire \DFF_1283.D ;
  wire \DFF_1283.Q ;
  wire \DFF_1284.CK ;
  wire \DFF_1284.D ;
  wire \DFF_1284.Q ;
  wire \DFF_1285.CK ;
  wire \DFF_1285.D ;
  wire \DFF_1285.Q ;
  wire \DFF_1286.CK ;
  wire \DFF_1286.D ;
  wire \DFF_1286.Q ;
  wire \DFF_1287.CK ;
  wire \DFF_1287.D ;
  wire \DFF_1287.Q ;
  wire \DFF_1288.CK ;
  wire \DFF_1288.D ;
  wire \DFF_1288.Q ;
  wire \DFF_1289.CK ;
  wire \DFF_1289.D ;
  wire \DFF_1289.Q ;
  wire \DFF_129.CK ;
  wire \DFF_129.D ;
  wire \DFF_129.Q ;
  wire \DFF_1290.CK ;
  wire \DFF_1290.D ;
  wire \DFF_1290.Q ;
  wire \DFF_1291.CK ;
  wire \DFF_1291.D ;
  wire \DFF_1291.Q ;
  wire \DFF_1292.CK ;
  wire \DFF_1292.D ;
  wire \DFF_1292.Q ;
  wire \DFF_1293.CK ;
  wire \DFF_1293.D ;
  wire \DFF_1293.Q ;
  wire \DFF_1294.CK ;
  wire \DFF_1294.D ;
  wire \DFF_1294.Q ;
  wire \DFF_1295.CK ;
  wire \DFF_1295.D ;
  wire \DFF_1295.Q ;
  wire \DFF_1296.CK ;
  wire \DFF_1296.D ;
  wire \DFF_1296.Q ;
  wire \DFF_1297.CK ;
  wire \DFF_1297.D ;
  wire \DFF_1297.Q ;
  wire \DFF_1298.CK ;
  wire \DFF_1298.D ;
  wire \DFF_1298.Q ;
  wire \DFF_1299.CK ;
  wire \DFF_1299.D ;
  wire \DFF_1299.Q ;
  wire \DFF_13.CK ;
  wire \DFF_13.D ;
  wire \DFF_13.Q ;
  wire \DFF_130.CK ;
  wire \DFF_130.D ;
  wire \DFF_130.Q ;
  wire \DFF_1300.CK ;
  wire \DFF_1300.D ;
  wire \DFF_1300.Q ;
  wire \DFF_1301.CK ;
  wire \DFF_1301.D ;
  wire \DFF_1301.Q ;
  wire \DFF_1302.CK ;
  wire \DFF_1302.D ;
  wire \DFF_1302.Q ;
  wire \DFF_1303.CK ;
  wire \DFF_1303.D ;
  wire \DFF_1303.Q ;
  wire \DFF_1304.CK ;
  wire \DFF_1304.D ;
  wire \DFF_1304.Q ;
  wire \DFF_1305.CK ;
  wire \DFF_1305.D ;
  wire \DFF_1305.Q ;
  wire \DFF_1306.CK ;
  wire \DFF_1306.D ;
  wire \DFF_1306.Q ;
  wire \DFF_1307.CK ;
  wire \DFF_1307.D ;
  wire \DFF_1307.Q ;
  wire \DFF_1308.CK ;
  wire \DFF_1308.D ;
  wire \DFF_1308.Q ;
  wire \DFF_1309.CK ;
  wire \DFF_1309.D ;
  wire \DFF_1309.Q ;
  wire \DFF_131.CK ;
  wire \DFF_131.D ;
  wire \DFF_131.Q ;
  wire \DFF_1310.CK ;
  wire \DFF_1310.D ;
  wire \DFF_1310.Q ;
  wire \DFF_1311.CK ;
  wire \DFF_1311.D ;
  wire \DFF_1311.Q ;
  wire \DFF_1312.CK ;
  wire \DFF_1312.D ;
  wire \DFF_1312.Q ;
  wire \DFF_1313.CK ;
  wire \DFF_1313.D ;
  wire \DFF_1313.Q ;
  wire \DFF_1314.CK ;
  wire \DFF_1314.D ;
  wire \DFF_1314.Q ;
  wire \DFF_1315.CK ;
  wire \DFF_1315.D ;
  wire \DFF_1315.Q ;
  wire \DFF_1316.CK ;
  wire \DFF_1316.D ;
  wire \DFF_1316.Q ;
  wire \DFF_1317.CK ;
  wire \DFF_1317.D ;
  wire \DFF_1317.Q ;
  wire \DFF_1318.CK ;
  wire \DFF_1318.D ;
  wire \DFF_1318.Q ;
  wire \DFF_1319.CK ;
  wire \DFF_1319.D ;
  wire \DFF_1319.Q ;
  wire \DFF_132.CK ;
  wire \DFF_132.D ;
  wire \DFF_132.Q ;
  wire \DFF_1320.CK ;
  wire \DFF_1320.D ;
  wire \DFF_1320.Q ;
  wire \DFF_1321.CK ;
  wire \DFF_1321.D ;
  wire \DFF_1321.Q ;
  wire \DFF_1322.CK ;
  wire \DFF_1322.D ;
  wire \DFF_1322.Q ;
  wire \DFF_1323.CK ;
  wire \DFF_1323.D ;
  wire \DFF_1323.Q ;
  wire \DFF_1324.CK ;
  wire \DFF_1324.D ;
  wire \DFF_1324.Q ;
  wire \DFF_1325.CK ;
  wire \DFF_1325.D ;
  wire \DFF_1325.Q ;
  wire \DFF_1326.CK ;
  wire \DFF_1326.D ;
  wire \DFF_1326.Q ;
  wire \DFF_1327.CK ;
  wire \DFF_1327.D ;
  wire \DFF_1327.Q ;
  wire \DFF_1328.CK ;
  wire \DFF_1328.D ;
  wire \DFF_1328.Q ;
  wire \DFF_1329.CK ;
  wire \DFF_1329.D ;
  wire \DFF_1329.Q ;
  wire \DFF_133.CK ;
  wire \DFF_133.D ;
  wire \DFF_133.Q ;
  wire \DFF_1330.CK ;
  wire \DFF_1330.D ;
  wire \DFF_1330.Q ;
  wire \DFF_1331.CK ;
  wire \DFF_1331.D ;
  wire \DFF_1331.Q ;
  wire \DFF_1332.CK ;
  wire \DFF_1332.D ;
  wire \DFF_1332.Q ;
  wire \DFF_1333.CK ;
  wire \DFF_1333.D ;
  wire \DFF_1333.Q ;
  wire \DFF_1334.CK ;
  wire \DFF_1334.D ;
  wire \DFF_1334.Q ;
  wire \DFF_1335.CK ;
  wire \DFF_1335.D ;
  wire \DFF_1335.Q ;
  wire \DFF_1336.CK ;
  wire \DFF_1336.D ;
  wire \DFF_1336.Q ;
  wire \DFF_1337.CK ;
  wire \DFF_1337.D ;
  wire \DFF_1337.Q ;
  wire \DFF_1338.CK ;
  wire \DFF_1338.D ;
  wire \DFF_1338.Q ;
  wire \DFF_1339.CK ;
  wire \DFF_1339.D ;
  wire \DFF_1339.Q ;
  wire \DFF_134.CK ;
  wire \DFF_134.D ;
  wire \DFF_134.Q ;
  wire \DFF_1340.CK ;
  wire \DFF_1340.D ;
  wire \DFF_1340.Q ;
  wire \DFF_1341.CK ;
  wire \DFF_1341.D ;
  wire \DFF_1341.Q ;
  wire \DFF_1342.CK ;
  wire \DFF_1342.D ;
  wire \DFF_1342.Q ;
  wire \DFF_1343.CK ;
  wire \DFF_1343.D ;
  wire \DFF_1343.Q ;
  wire \DFF_1344.CK ;
  wire \DFF_1344.D ;
  wire \DFF_1344.Q ;
  wire \DFF_1345.CK ;
  wire \DFF_1345.D ;
  wire \DFF_1345.Q ;
  wire \DFF_1346.CK ;
  wire \DFF_1346.D ;
  wire \DFF_1346.Q ;
  wire \DFF_1347.CK ;
  wire \DFF_1347.D ;
  wire \DFF_1347.Q ;
  wire \DFF_1348.CK ;
  wire \DFF_1348.D ;
  wire \DFF_1348.Q ;
  wire \DFF_1349.CK ;
  wire \DFF_1349.D ;
  wire \DFF_1349.Q ;
  wire \DFF_135.CK ;
  wire \DFF_135.D ;
  wire \DFF_135.Q ;
  wire \DFF_1350.CK ;
  wire \DFF_1350.D ;
  wire \DFF_1350.Q ;
  wire \DFF_1351.CK ;
  wire \DFF_1351.D ;
  wire \DFF_1351.Q ;
  wire \DFF_1352.CK ;
  wire \DFF_1352.D ;
  wire \DFF_1352.Q ;
  wire \DFF_1353.CK ;
  wire \DFF_1353.D ;
  wire \DFF_1353.Q ;
  wire \DFF_1354.CK ;
  wire \DFF_1354.D ;
  wire \DFF_1354.Q ;
  wire \DFF_1355.CK ;
  wire \DFF_1355.D ;
  wire \DFF_1355.Q ;
  wire \DFF_1356.CK ;
  wire \DFF_1356.D ;
  wire \DFF_1356.Q ;
  wire \DFF_1357.CK ;
  wire \DFF_1357.D ;
  wire \DFF_1357.Q ;
  wire \DFF_1358.CK ;
  wire \DFF_1358.D ;
  wire \DFF_1358.Q ;
  wire \DFF_1359.CK ;
  wire \DFF_1359.D ;
  wire \DFF_1359.Q ;
  wire \DFF_136.CK ;
  wire \DFF_136.D ;
  wire \DFF_136.Q ;
  wire \DFF_1360.CK ;
  wire \DFF_1360.D ;
  wire \DFF_1360.Q ;
  wire \DFF_1361.CK ;
  wire \DFF_1361.D ;
  wire \DFF_1361.Q ;
  wire \DFF_1362.CK ;
  wire \DFF_1362.D ;
  wire \DFF_1362.Q ;
  wire \DFF_1363.CK ;
  wire \DFF_1363.D ;
  wire \DFF_1363.Q ;
  wire \DFF_1364.CK ;
  wire \DFF_1364.D ;
  wire \DFF_1364.Q ;
  wire \DFF_1365.CK ;
  wire \DFF_1365.D ;
  wire \DFF_1365.Q ;
  wire \DFF_1366.CK ;
  wire \DFF_1366.D ;
  wire \DFF_1366.Q ;
  wire \DFF_1367.CK ;
  wire \DFF_1367.D ;
  wire \DFF_1367.Q ;
  wire \DFF_1368.CK ;
  wire \DFF_1369.CK ;
  wire \DFF_137.CK ;
  wire \DFF_137.D ;
  wire \DFF_137.Q ;
  wire \DFF_1370.CK ;
  wire \DFF_1371.CK ;
  wire \DFF_1372.CK ;
  wire \DFF_1373.CK ;
  wire \DFF_1374.CK ;
  wire \DFF_1375.CK ;
  wire \DFF_1376.CK ;
  wire \DFF_1377.CK ;
  wire \DFF_1378.CK ;
  wire \DFF_1378.D ;
  wire \DFF_1378.Q ;
  wire \DFF_1379.CK ;
  wire \DFF_1379.D ;
  wire \DFF_1379.Q ;
  wire \DFF_138.CK ;
  wire \DFF_138.D ;
  wire \DFF_138.Q ;
  wire \DFF_1380.CK ;
  wire \DFF_1380.D ;
  wire \DFF_1380.Q ;
  wire \DFF_1381.CK ;
  wire \DFF_1381.D ;
  wire \DFF_1381.Q ;
  wire \DFF_1382.CK ;
  wire \DFF_1382.D ;
  wire \DFF_1382.Q ;
  wire \DFF_1383.CK ;
  wire \DFF_1383.D ;
  wire \DFF_1383.Q ;
  wire \DFF_1384.CK ;
  wire \DFF_1384.D ;
  wire \DFF_1384.Q ;
  wire \DFF_1385.CK ;
  wire \DFF_1385.D ;
  wire \DFF_1385.Q ;
  wire \DFF_1386.CK ;
  wire \DFF_1386.D ;
  wire \DFF_1386.Q ;
  wire \DFF_1387.CK ;
  wire \DFF_1387.D ;
  wire \DFF_1387.Q ;
  wire \DFF_1388.CK ;
  wire \DFF_1388.D ;
  wire \DFF_1388.Q ;
  wire \DFF_1389.CK ;
  wire \DFF_1389.D ;
  wire \DFF_1389.Q ;
  wire \DFF_139.CK ;
  wire \DFF_139.D ;
  wire \DFF_139.Q ;
  wire \DFF_1390.CK ;
  wire \DFF_1390.D ;
  wire \DFF_1390.Q ;
  wire \DFF_1391.CK ;
  wire \DFF_1391.D ;
  wire \DFF_1391.Q ;
  wire \DFF_1392.CK ;
  wire \DFF_1392.D ;
  wire \DFF_1392.Q ;
  wire \DFF_1393.CK ;
  wire \DFF_1393.D ;
  wire \DFF_1393.Q ;
  wire \DFF_1394.CK ;
  wire \DFF_1394.D ;
  wire \DFF_1394.Q ;
  wire \DFF_1395.CK ;
  wire \DFF_1395.D ;
  wire \DFF_1395.Q ;
  wire \DFF_1396.CK ;
  wire \DFF_1396.D ;
  wire \DFF_1396.Q ;
  wire \DFF_1397.CK ;
  wire \DFF_1397.D ;
  wire \DFF_1397.Q ;
  wire \DFF_1398.CK ;
  wire \DFF_1398.D ;
  wire \DFF_1398.Q ;
  wire \DFF_1399.CK ;
  wire \DFF_1399.D ;
  wire \DFF_1399.Q ;
  wire \DFF_14.CK ;
  wire \DFF_14.D ;
  wire \DFF_14.Q ;
  wire \DFF_140.CK ;
  wire \DFF_140.D ;
  wire \DFF_140.Q ;
  wire \DFF_1400.CK ;
  wire \DFF_1400.D ;
  wire \DFF_1400.Q ;
  wire \DFF_1401.CK ;
  wire \DFF_1401.D ;
  wire \DFF_1401.Q ;
  wire \DFF_1402.CK ;
  wire \DFF_1402.D ;
  wire \DFF_1402.Q ;
  wire \DFF_1403.CK ;
  wire \DFF_1403.D ;
  wire \DFF_1403.Q ;
  wire \DFF_1404.CK ;
  wire \DFF_1404.D ;
  wire \DFF_1404.Q ;
  wire \DFF_1405.CK ;
  wire \DFF_1405.D ;
  wire \DFF_1405.Q ;
  wire \DFF_1406.CK ;
  wire \DFF_1406.D ;
  wire \DFF_1406.Q ;
  wire \DFF_1407.CK ;
  wire \DFF_1407.D ;
  wire \DFF_1407.Q ;
  wire \DFF_1408.CK ;
  wire \DFF_1408.D ;
  wire \DFF_1408.Q ;
  wire \DFF_1409.CK ;
  wire \DFF_1409.D ;
  wire \DFF_1409.Q ;
  wire \DFF_141.CK ;
  wire \DFF_141.D ;
  wire \DFF_141.Q ;
  wire \DFF_1410.CK ;
  wire \DFF_1410.D ;
  wire \DFF_1410.Q ;
  wire \DFF_1411.CK ;
  wire \DFF_1411.D ;
  wire \DFF_1411.Q ;
  wire \DFF_1412.CK ;
  wire \DFF_1412.D ;
  wire \DFF_1412.Q ;
  wire \DFF_1413.CK ;
  wire \DFF_1413.D ;
  wire \DFF_1413.Q ;
  wire \DFF_1414.CK ;
  wire \DFF_1414.D ;
  wire \DFF_1414.Q ;
  wire \DFF_1415.CK ;
  wire \DFF_1415.D ;
  wire \DFF_1415.Q ;
  wire \DFF_1416.CK ;
  wire \DFF_1416.D ;
  wire \DFF_1416.Q ;
  wire \DFF_1417.CK ;
  wire \DFF_1417.D ;
  wire \DFF_1417.Q ;
  wire \DFF_1418.CK ;
  wire \DFF_1418.D ;
  wire \DFF_1418.Q ;
  wire \DFF_1419.CK ;
  wire \DFF_1419.D ;
  wire \DFF_1419.Q ;
  wire \DFF_142.CK ;
  wire \DFF_142.D ;
  wire \DFF_142.Q ;
  wire \DFF_1420.CK ;
  wire \DFF_1420.D ;
  wire \DFF_1420.Q ;
  wire \DFF_1421.CK ;
  wire \DFF_1421.D ;
  wire \DFF_1421.Q ;
  wire \DFF_1422.CK ;
  wire \DFF_1422.D ;
  wire \DFF_1422.Q ;
  wire \DFF_1423.CK ;
  wire \DFF_1423.D ;
  wire \DFF_1423.Q ;
  wire \DFF_1424.CK ;
  wire \DFF_1424.D ;
  wire \DFF_1424.Q ;
  wire \DFF_1425.CK ;
  wire \DFF_1425.D ;
  wire \DFF_1425.Q ;
  wire \DFF_1426.CK ;
  wire \DFF_1426.D ;
  wire \DFF_1426.Q ;
  wire \DFF_1427.CK ;
  wire \DFF_1427.D ;
  wire \DFF_1427.Q ;
  wire \DFF_1428.CK ;
  wire \DFF_1428.D ;
  wire \DFF_1428.Q ;
  wire \DFF_1429.CK ;
  wire \DFF_1429.D ;
  wire \DFF_1429.Q ;
  wire \DFF_143.CK ;
  wire \DFF_143.D ;
  wire \DFF_143.Q ;
  wire \DFF_1430.CK ;
  wire \DFF_1430.D ;
  wire \DFF_1430.Q ;
  wire \DFF_1431.CK ;
  wire \DFF_1431.D ;
  wire \DFF_1431.Q ;
  wire \DFF_1432.CK ;
  wire \DFF_1432.D ;
  wire \DFF_1432.Q ;
  wire \DFF_1433.CK ;
  wire \DFF_1433.D ;
  wire \DFF_1433.Q ;
  wire \DFF_1434.CK ;
  wire \DFF_1434.D ;
  wire \DFF_1434.Q ;
  wire \DFF_1435.CK ;
  wire \DFF_1435.D ;
  wire \DFF_1435.Q ;
  wire \DFF_1436.CK ;
  wire \DFF_1436.D ;
  wire \DFF_1436.Q ;
  wire \DFF_1437.CK ;
  wire \DFF_1437.D ;
  wire \DFF_1437.Q ;
  wire \DFF_1438.CK ;
  wire \DFF_1438.D ;
  wire \DFF_1438.Q ;
  wire \DFF_1439.CK ;
  wire \DFF_1439.D ;
  wire \DFF_1439.Q ;
  wire \DFF_144.CK ;
  wire \DFF_144.D ;
  wire \DFF_144.Q ;
  wire \DFF_1440.CK ;
  wire \DFF_1440.D ;
  wire \DFF_1440.Q ;
  wire \DFF_1441.CK ;
  wire \DFF_1441.D ;
  wire \DFF_1441.Q ;
  wire \DFF_1442.CK ;
  wire \DFF_1442.D ;
  wire \DFF_1442.Q ;
  wire \DFF_1443.CK ;
  wire \DFF_1443.D ;
  wire \DFF_1443.Q ;
  wire \DFF_1444.CK ;
  wire \DFF_1444.D ;
  wire \DFF_1444.Q ;
  wire \DFF_1445.CK ;
  wire \DFF_1445.D ;
  wire \DFF_1445.Q ;
  wire \DFF_1446.CK ;
  wire \DFF_1446.D ;
  wire \DFF_1446.Q ;
  wire \DFF_1447.CK ;
  wire \DFF_1447.D ;
  wire \DFF_1447.Q ;
  wire \DFF_1448.CK ;
  wire \DFF_1448.D ;
  wire \DFF_1448.Q ;
  wire \DFF_1449.CK ;
  wire \DFF_1449.D ;
  wire \DFF_1449.Q ;
  wire \DFF_145.CK ;
  wire \DFF_145.D ;
  wire \DFF_145.Q ;
  wire \DFF_1450.CK ;
  wire \DFF_1450.D ;
  wire \DFF_1450.Q ;
  wire \DFF_1451.CK ;
  wire \DFF_1451.D ;
  wire \DFF_1451.Q ;
  wire \DFF_1452.CK ;
  wire \DFF_1452.D ;
  wire \DFF_1452.Q ;
  wire \DFF_1453.CK ;
  wire \DFF_1453.D ;
  wire \DFF_1453.Q ;
  wire \DFF_1454.CK ;
  wire \DFF_1454.D ;
  wire \DFF_1454.Q ;
  wire \DFF_1455.CK ;
  wire \DFF_1455.D ;
  wire \DFF_1455.Q ;
  wire \DFF_1456.CK ;
  wire \DFF_1456.D ;
  wire \DFF_1456.Q ;
  wire \DFF_1457.CK ;
  wire \DFF_1457.D ;
  wire \DFF_1457.Q ;
  wire \DFF_1458.CK ;
  wire \DFF_1458.D ;
  wire \DFF_1458.Q ;
  wire \DFF_1459.CK ;
  wire \DFF_1459.D ;
  wire \DFF_1459.Q ;
  wire \DFF_146.CK ;
  wire \DFF_146.D ;
  wire \DFF_146.Q ;
  wire \DFF_1460.CK ;
  wire \DFF_1460.D ;
  wire \DFF_1460.Q ;
  wire \DFF_1461.CK ;
  wire \DFF_1461.D ;
  wire \DFF_1461.Q ;
  wire \DFF_1462.CK ;
  wire \DFF_1462.D ;
  wire \DFF_1462.Q ;
  wire \DFF_1463.CK ;
  wire \DFF_1463.D ;
  wire \DFF_1463.Q ;
  wire \DFF_1464.CK ;
  wire \DFF_1464.D ;
  wire \DFF_1464.Q ;
  wire \DFF_1465.CK ;
  wire \DFF_1465.D ;
  wire \DFF_1465.Q ;
  wire \DFF_1466.CK ;
  wire \DFF_1466.D ;
  wire \DFF_1466.Q ;
  wire \DFF_1467.CK ;
  wire \DFF_1467.D ;
  wire \DFF_1467.Q ;
  wire \DFF_1468.CK ;
  wire \DFF_1468.D ;
  wire \DFF_1468.Q ;
  wire \DFF_1469.CK ;
  wire \DFF_1469.D ;
  wire \DFF_1469.Q ;
  wire \DFF_147.CK ;
  wire \DFF_147.D ;
  wire \DFF_147.Q ;
  wire \DFF_1470.CK ;
  wire \DFF_1470.D ;
  wire \DFF_1470.Q ;
  wire \DFF_1471.CK ;
  wire \DFF_1471.D ;
  wire \DFF_1471.Q ;
  wire \DFF_1472.CK ;
  wire \DFF_1472.D ;
  wire \DFF_1472.Q ;
  wire \DFF_1473.CK ;
  wire \DFF_1473.D ;
  wire \DFF_1473.Q ;
  wire \DFF_1474.CK ;
  wire \DFF_1474.D ;
  wire \DFF_1474.Q ;
  wire \DFF_1475.CK ;
  wire \DFF_1475.D ;
  wire \DFF_1475.Q ;
  wire \DFF_1476.CK ;
  wire \DFF_1476.D ;
  wire \DFF_1476.Q ;
  wire \DFF_1477.CK ;
  wire \DFF_1477.D ;
  wire \DFF_1477.Q ;
  wire \DFF_1478.CK ;
  wire \DFF_1478.D ;
  wire \DFF_1478.Q ;
  wire \DFF_1479.CK ;
  wire \DFF_1479.D ;
  wire \DFF_1479.Q ;
  wire \DFF_148.CK ;
  wire \DFF_148.D ;
  wire \DFF_148.Q ;
  wire \DFF_1480.CK ;
  wire \DFF_1480.D ;
  wire \DFF_1480.Q ;
  wire \DFF_1481.CK ;
  wire \DFF_1481.D ;
  wire \DFF_1481.Q ;
  wire \DFF_1482.CK ;
  wire \DFF_1482.D ;
  wire \DFF_1482.Q ;
  wire \DFF_1483.CK ;
  wire \DFF_1483.D ;
  wire \DFF_1483.Q ;
  wire \DFF_1484.CK ;
  wire \DFF_1485.CK ;
  wire \DFF_1486.CK ;
  wire \DFF_1487.CK ;
  wire \DFF_1488.CK ;
  wire \DFF_1489.CK ;
  wire \DFF_149.CK ;
  wire \DFF_149.D ;
  wire \DFF_149.Q ;
  wire \DFF_1490.CK ;
  wire \DFF_1491.CK ;
  wire \DFF_1492.CK ;
  wire \DFF_1492.D ;
  wire \DFF_1492.Q ;
  wire \DFF_1493.CK ;
  wire \DFF_1493.D ;
  wire \DFF_1493.Q ;
  wire \DFF_1494.CK ;
  wire \DFF_1494.D ;
  wire \DFF_1494.Q ;
  wire \DFF_1495.CK ;
  wire \DFF_1495.D ;
  wire \DFF_1495.Q ;
  wire \DFF_1496.CK ;
  wire \DFF_1496.D ;
  wire \DFF_1496.Q ;
  wire \DFF_1497.CK ;
  wire \DFF_1497.D ;
  wire \DFF_1497.Q ;
  wire \DFF_1498.CK ;
  wire \DFF_1498.D ;
  wire \DFF_1498.Q ;
  wire \DFF_1499.CK ;
  wire \DFF_1499.D ;
  wire \DFF_1499.Q ;
  wire \DFF_15.CK ;
  wire \DFF_15.D ;
  wire \DFF_15.Q ;
  wire \DFF_150.CK ;
  wire \DFF_150.D ;
  wire \DFF_150.Q ;
  wire \DFF_1500.CK ;
  wire \DFF_1500.D ;
  wire \DFF_1500.Q ;
  wire \DFF_1501.CK ;
  wire \DFF_1501.D ;
  wire \DFF_1501.Q ;
  wire \DFF_1502.CK ;
  wire \DFF_1502.D ;
  wire \DFF_1502.Q ;
  wire \DFF_1503.CK ;
  wire \DFF_1503.D ;
  wire \DFF_1503.Q ;
  wire \DFF_1504.CK ;
  wire \DFF_1504.D ;
  wire \DFF_1504.Q ;
  wire \DFF_1505.CK ;
  wire \DFF_1505.D ;
  wire \DFF_1505.Q ;
  wire \DFF_1506.CK ;
  wire \DFF_1506.D ;
  wire \DFF_1506.Q ;
  wire \DFF_1507.CK ;
  wire \DFF_1507.D ;
  wire \DFF_1507.Q ;
  wire \DFF_1508.CK ;
  wire \DFF_1508.D ;
  wire \DFF_1508.Q ;
  wire \DFF_1509.CK ;
  wire \DFF_1509.D ;
  wire \DFF_1509.Q ;
  wire \DFF_151.CK ;
  wire \DFF_151.D ;
  wire \DFF_151.Q ;
  wire \DFF_1510.CK ;
  wire \DFF_1510.D ;
  wire \DFF_1510.Q ;
  wire \DFF_1511.CK ;
  wire \DFF_1511.D ;
  wire \DFF_1511.Q ;
  wire \DFF_1512.CK ;
  wire \DFF_1512.D ;
  wire \DFF_1512.Q ;
  wire \DFF_1513.CK ;
  wire \DFF_1513.D ;
  wire \DFF_1513.Q ;
  wire \DFF_1514.CK ;
  wire \DFF_1514.D ;
  wire \DFF_1514.Q ;
  wire \DFF_1515.CK ;
  wire \DFF_1515.D ;
  wire \DFF_1515.Q ;
  wire \DFF_1516.CK ;
  wire \DFF_1516.D ;
  wire \DFF_1516.Q ;
  wire \DFF_1517.CK ;
  wire \DFF_1517.D ;
  wire \DFF_1517.Q ;
  wire \DFF_1518.CK ;
  wire \DFF_1518.D ;
  wire \DFF_1518.Q ;
  wire \DFF_1519.CK ;
  wire \DFF_1519.D ;
  wire \DFF_1519.Q ;
  wire \DFF_152.CK ;
  wire \DFF_152.D ;
  wire \DFF_152.Q ;
  wire \DFF_1520.CK ;
  wire \DFF_1520.D ;
  wire \DFF_1520.Q ;
  wire \DFF_1521.CK ;
  wire \DFF_1521.D ;
  wire \DFF_1521.Q ;
  wire \DFF_1522.CK ;
  wire \DFF_1522.D ;
  wire \DFF_1522.Q ;
  wire \DFF_1523.CK ;
  wire \DFF_1523.D ;
  wire \DFF_1523.Q ;
  wire \DFF_1524.CK ;
  wire \DFF_1524.D ;
  wire \DFF_1524.Q ;
  wire \DFF_1525.CK ;
  wire \DFF_1525.D ;
  wire \DFF_1525.Q ;
  wire \DFF_1526.CK ;
  wire \DFF_1526.D ;
  wire \DFF_1526.Q ;
  wire \DFF_1527.CK ;
  wire \DFF_1527.D ;
  wire \DFF_1527.Q ;
  wire \DFF_1528.CK ;
  wire \DFF_1528.D ;
  wire \DFF_1528.Q ;
  wire \DFF_1529.CK ;
  wire \DFF_1529.D ;
  wire \DFF_1529.Q ;
  wire \DFF_153.CK ;
  wire \DFF_153.D ;
  wire \DFF_153.Q ;
  wire \DFF_1530.CK ;
  wire \DFF_1530.D ;
  wire \DFF_1530.Q ;
  wire \DFF_1531.CK ;
  wire \DFF_1531.D ;
  wire \DFF_1531.Q ;
  wire \DFF_1532.CK ;
  wire \DFF_1532.D ;
  wire \DFF_1532.Q ;
  wire \DFF_1533.CK ;
  wire \DFF_1533.D ;
  wire \DFF_1533.Q ;
  wire \DFF_1534.CK ;
  wire \DFF_1534.D ;
  wire \DFF_1534.Q ;
  wire \DFF_1535.CK ;
  wire \DFF_1535.D ;
  wire \DFF_1535.Q ;
  wire \DFF_1536.CK ;
  wire \DFF_1536.D ;
  wire \DFF_1536.Q ;
  wire \DFF_1537.CK ;
  wire \DFF_1537.D ;
  wire \DFF_1537.Q ;
  wire \DFF_1538.CK ;
  wire \DFF_1538.D ;
  wire \DFF_1538.Q ;
  wire \DFF_1539.CK ;
  wire \DFF_1539.D ;
  wire \DFF_1539.Q ;
  wire \DFF_154.CK ;
  wire \DFF_154.D ;
  wire \DFF_154.Q ;
  wire \DFF_1540.CK ;
  wire \DFF_1540.D ;
  wire \DFF_1540.Q ;
  wire \DFF_1541.CK ;
  wire \DFF_1541.D ;
  wire \DFF_1541.Q ;
  wire \DFF_1542.CK ;
  wire \DFF_1542.D ;
  wire \DFF_1542.Q ;
  wire \DFF_1543.CK ;
  wire \DFF_1543.D ;
  wire \DFF_1543.Q ;
  wire \DFF_1544.CK ;
  wire \DFF_1544.D ;
  wire \DFF_1544.Q ;
  wire \DFF_1545.CK ;
  wire \DFF_1545.D ;
  wire \DFF_1545.Q ;
  wire \DFF_1546.CK ;
  wire \DFF_1546.D ;
  wire \DFF_1546.Q ;
  wire \DFF_1547.CK ;
  wire \DFF_1547.D ;
  wire \DFF_1547.Q ;
  wire \DFF_1548.CK ;
  wire \DFF_1548.D ;
  wire \DFF_1548.Q ;
  wire \DFF_1549.CK ;
  wire \DFF_1549.D ;
  wire \DFF_1549.Q ;
  wire \DFF_155.CK ;
  wire \DFF_155.D ;
  wire \DFF_155.Q ;
  wire \DFF_1550.CK ;
  wire \DFF_1550.D ;
  wire \DFF_1550.Q ;
  wire \DFF_1551.CK ;
  wire \DFF_1551.D ;
  wire \DFF_1551.Q ;
  wire \DFF_1552.CK ;
  wire \DFF_1552.D ;
  wire \DFF_1552.Q ;
  wire \DFF_1553.CK ;
  wire \DFF_1553.D ;
  wire \DFF_1553.Q ;
  wire \DFF_1554.CK ;
  wire \DFF_1554.D ;
  wire \DFF_1554.Q ;
  wire \DFF_1555.CK ;
  wire \DFF_1555.D ;
  wire \DFF_1555.Q ;
  wire \DFF_1556.CK ;
  wire \DFF_1556.D ;
  wire \DFF_1556.Q ;
  wire \DFF_1557.CK ;
  wire \DFF_1557.D ;
  wire \DFF_1557.Q ;
  wire \DFF_1558.CK ;
  wire \DFF_1558.D ;
  wire \DFF_1558.Q ;
  wire \DFF_1559.CK ;
  wire \DFF_1559.D ;
  wire \DFF_1559.Q ;
  wire \DFF_156.CK ;
  wire \DFF_156.D ;
  wire \DFF_156.Q ;
  wire \DFF_1560.CK ;
  wire \DFF_1560.D ;
  wire \DFF_1560.Q ;
  wire \DFF_1561.CK ;
  wire \DFF_1561.D ;
  wire \DFF_1561.Q ;
  wire \DFF_1562.CK ;
  wire \DFF_1562.D ;
  wire \DFF_1562.Q ;
  wire \DFF_1563.CK ;
  wire \DFF_1563.D ;
  wire \DFF_1563.Q ;
  wire \DFF_1564.CK ;
  wire \DFF_1564.D ;
  wire \DFF_1564.Q ;
  wire \DFF_1565.CK ;
  wire \DFF_1565.D ;
  wire \DFF_1565.Q ;
  wire \DFF_1566.CK ;
  wire \DFF_1566.D ;
  wire \DFF_1566.Q ;
  wire \DFF_1567.CK ;
  wire \DFF_1567.D ;
  wire \DFF_1567.Q ;
  wire \DFF_1568.CK ;
  wire \DFF_1568.D ;
  wire \DFF_1568.Q ;
  wire \DFF_1569.CK ;
  wire \DFF_1569.D ;
  wire \DFF_1569.Q ;
  wire \DFF_157.CK ;
  wire \DFF_157.D ;
  wire \DFF_157.Q ;
  wire \DFF_1570.CK ;
  wire \DFF_1570.D ;
  wire \DFF_1570.Q ;
  wire \DFF_1571.CK ;
  wire \DFF_1571.D ;
  wire \DFF_1571.Q ;
  wire \DFF_1572.CK ;
  wire \DFF_1572.D ;
  wire \DFF_1572.Q ;
  wire \DFF_1573.CK ;
  wire \DFF_1573.D ;
  wire \DFF_1573.Q ;
  wire \DFF_1574.CK ;
  wire \DFF_1574.D ;
  wire \DFF_1574.Q ;
  wire \DFF_1575.CK ;
  wire \DFF_1575.D ;
  wire \DFF_1575.Q ;
  wire \DFF_1576.CK ;
  wire \DFF_1576.D ;
  wire \DFF_1576.Q ;
  wire \DFF_1577.CK ;
  wire \DFF_1577.D ;
  wire \DFF_1577.Q ;
  wire \DFF_1578.CK ;
  wire \DFF_1578.D ;
  wire \DFF_1578.Q ;
  wire \DFF_1579.CK ;
  wire \DFF_1579.D ;
  wire \DFF_1579.Q ;
  wire \DFF_158.CK ;
  wire \DFF_158.D ;
  wire \DFF_158.Q ;
  wire \DFF_1580.CK ;
  wire \DFF_1580.D ;
  wire \DFF_1580.Q ;
  wire \DFF_1581.CK ;
  wire \DFF_1581.D ;
  wire \DFF_1581.Q ;
  wire \DFF_1582.CK ;
  wire \DFF_1582.D ;
  wire \DFF_1582.Q ;
  wire \DFF_1583.CK ;
  wire \DFF_1583.D ;
  wire \DFF_1583.Q ;
  wire \DFF_1584.CK ;
  wire \DFF_1584.D ;
  wire \DFF_1584.Q ;
  wire \DFF_1585.CK ;
  wire \DFF_1585.D ;
  wire \DFF_1585.Q ;
  wire \DFF_1586.CK ;
  wire \DFF_1586.D ;
  wire \DFF_1586.Q ;
  wire \DFF_1587.CK ;
  wire \DFF_1587.D ;
  wire \DFF_1587.Q ;
  wire \DFF_1588.CK ;
  wire \DFF_1588.D ;
  wire \DFF_1588.Q ;
  wire \DFF_1589.CK ;
  wire \DFF_1589.D ;
  wire \DFF_1589.Q ;
  wire \DFF_159.CK ;
  wire \DFF_159.D ;
  wire \DFF_159.Q ;
  wire \DFF_1590.CK ;
  wire \DFF_1590.D ;
  wire \DFF_1590.Q ;
  wire \DFF_1591.CK ;
  wire \DFF_1591.D ;
  wire \DFF_1591.Q ;
  wire \DFF_1592.CK ;
  wire \DFF_1592.D ;
  wire \DFF_1592.Q ;
  wire \DFF_1593.CK ;
  wire \DFF_1593.D ;
  wire \DFF_1593.Q ;
  wire \DFF_1594.CK ;
  wire \DFF_1594.D ;
  wire \DFF_1594.Q ;
  wire \DFF_1595.CK ;
  wire \DFF_1595.D ;
  wire \DFF_1595.Q ;
  wire \DFF_1596.CK ;
  wire \DFF_1596.D ;
  wire \DFF_1596.Q ;
  wire \DFF_1597.CK ;
  wire \DFF_1597.D ;
  wire \DFF_1597.Q ;
  wire \DFF_1598.CK ;
  wire \DFF_1598.D ;
  wire \DFF_1598.Q ;
  wire \DFF_1599.CK ;
  wire \DFF_1599.D ;
  wire \DFF_1599.Q ;
  wire \DFF_16.CK ;
  wire \DFF_16.D ;
  wire \DFF_16.Q ;
  wire \DFF_160.CK ;
  wire \DFF_160.D ;
  wire \DFF_160.Q ;
  wire \DFF_1600.CK ;
  wire \DFF_1600.D ;
  wire \DFF_1600.Q ;
  wire \DFF_1601.CK ;
  wire \DFF_1601.D ;
  wire \DFF_1601.Q ;
  wire \DFF_1602.CK ;
  wire \DFF_1602.D ;
  wire \DFF_1602.Q ;
  wire \DFF_1603.CK ;
  wire \DFF_1603.D ;
  wire \DFF_1603.Q ;
  wire \DFF_1604.CK ;
  wire \DFF_1604.D ;
  wire \DFF_1604.Q ;
  wire \DFF_1605.CK ;
  wire \DFF_1605.D ;
  wire \DFF_1605.Q ;
  wire \DFF_1606.CK ;
  wire \DFF_1606.D ;
  wire \DFF_1606.Q ;
  wire \DFF_1607.CK ;
  wire \DFF_1607.D ;
  wire \DFF_1607.Q ;
  wire \DFF_1608.CK ;
  wire \DFF_1608.D ;
  wire \DFF_1608.Q ;
  wire \DFF_1609.CK ;
  wire \DFF_1609.D ;
  wire \DFF_1609.Q ;
  wire \DFF_161.CK ;
  wire \DFF_161.D ;
  wire \DFF_161.Q ;
  wire \DFF_1610.CK ;
  wire \DFF_1610.D ;
  wire \DFF_1610.Q ;
  wire \DFF_1611.CK ;
  wire \DFF_1611.D ;
  wire \DFF_1611.Q ;
  wire \DFF_1612.CK ;
  wire \DFF_1612.D ;
  wire \DFF_1612.Q ;
  wire \DFF_1613.CK ;
  wire \DFF_1613.D ;
  wire \DFF_1613.Q ;
  wire \DFF_1614.CK ;
  wire \DFF_1614.D ;
  wire \DFF_1614.Q ;
  wire \DFF_1615.CK ;
  wire \DFF_1615.D ;
  wire \DFF_1615.Q ;
  wire \DFF_1616.CK ;
  wire \DFF_1616.D ;
  wire \DFF_1616.Q ;
  wire \DFF_1617.CK ;
  wire \DFF_1617.D ;
  wire \DFF_1617.Q ;
  wire \DFF_1618.CK ;
  wire \DFF_1618.D ;
  wire \DFF_1618.Q ;
  wire \DFF_1619.CK ;
  wire \DFF_1619.D ;
  wire \DFF_1619.Q ;
  wire \DFF_162.CK ;
  wire \DFF_162.D ;
  wire \DFF_162.Q ;
  wire \DFF_1620.CK ;
  wire \DFF_1620.D ;
  wire \DFF_1620.Q ;
  wire \DFF_1621.CK ;
  wire \DFF_1621.D ;
  wire \DFF_1621.Q ;
  wire \DFF_1622.CK ;
  wire \DFF_1622.D ;
  wire \DFF_1622.Q ;
  wire \DFF_1623.CK ;
  wire \DFF_1623.D ;
  wire \DFF_1623.Q ;
  wire \DFF_1624.CK ;
  wire \DFF_1624.D ;
  wire \DFF_1624.Q ;
  wire \DFF_1625.CK ;
  wire \DFF_1625.D ;
  wire \DFF_1625.Q ;
  wire \DFF_1626.CK ;
  wire \DFF_1626.D ;
  wire \DFF_1626.Q ;
  wire \DFF_1627.CK ;
  wire \DFF_1627.D ;
  wire \DFF_1627.Q ;
  wire \DFF_1628.CK ;
  wire \DFF_1628.D ;
  wire \DFF_1628.Q ;
  wire \DFF_1629.CK ;
  wire \DFF_1629.D ;
  wire \DFF_1629.Q ;
  wire \DFF_163.CK ;
  wire \DFF_163.D ;
  wire \DFF_163.Q ;
  wire \DFF_1630.CK ;
  wire \DFF_1630.D ;
  wire \DFF_1630.Q ;
  wire \DFF_1631.CK ;
  wire \DFF_1631.D ;
  wire \DFF_1631.Q ;
  wire \DFF_1632.CK ;
  wire \DFF_1632.D ;
  wire \DFF_1632.Q ;
  wire \DFF_1633.CK ;
  wire \DFF_1633.D ;
  wire \DFF_1633.Q ;
  wire \DFF_1634.CK ;
  wire \DFF_1634.D ;
  wire \DFF_1634.Q ;
  wire \DFF_1635.CK ;
  wire \DFF_1635.D ;
  wire \DFF_1635.Q ;
  wire \DFF_164.CK ;
  wire \DFF_164.D ;
  wire \DFF_164.Q ;
  wire \DFF_165.CK ;
  wire \DFF_165.D ;
  wire \DFF_165.Q ;
  wire \DFF_166.CK ;
  wire \DFF_166.D ;
  wire \DFF_166.Q ;
  wire \DFF_167.CK ;
  wire \DFF_167.D ;
  wire \DFF_167.Q ;
  wire \DFF_168.CK ;
  wire \DFF_168.D ;
  wire \DFF_168.Q ;
  wire \DFF_169.CK ;
  wire \DFF_169.D ;
  wire \DFF_169.Q ;
  wire \DFF_17.CK ;
  wire \DFF_17.D ;
  wire \DFF_17.Q ;
  wire \DFF_170.CK ;
  wire \DFF_170.D ;
  wire \DFF_170.Q ;
  wire \DFF_171.CK ;
  wire \DFF_171.D ;
  wire \DFF_171.Q ;
  wire \DFF_172.CK ;
  wire \DFF_172.D ;
  wire \DFF_172.Q ;
  wire \DFF_173.CK ;
  wire \DFF_173.D ;
  wire \DFF_173.Q ;
  wire \DFF_174.CK ;
  wire \DFF_174.D ;
  wire \DFF_174.Q ;
  wire \DFF_175.CK ;
  wire \DFF_175.D ;
  wire \DFF_175.Q ;
  wire \DFF_176.CK ;
  wire \DFF_176.D ;
  wire \DFF_176.Q ;
  wire \DFF_177.CK ;
  wire \DFF_177.D ;
  wire \DFF_177.Q ;
  wire \DFF_178.CK ;
  wire \DFF_178.D ;
  wire \DFF_178.Q ;
  wire \DFF_179.CK ;
  wire \DFF_179.D ;
  wire \DFF_179.Q ;
  wire \DFF_18.CK ;
  wire \DFF_18.D ;
  wire \DFF_18.Q ;
  wire \DFF_180.CK ;
  wire \DFF_180.D ;
  wire \DFF_180.Q ;
  wire \DFF_181.CK ;
  wire \DFF_181.D ;
  wire \DFF_181.Q ;
  wire \DFF_182.CK ;
  wire \DFF_182.D ;
  wire \DFF_182.Q ;
  wire \DFF_183.CK ;
  wire \DFF_183.D ;
  wire \DFF_183.Q ;
  wire \DFF_184.CK ;
  wire \DFF_184.D ;
  wire \DFF_184.Q ;
  wire \DFF_185.CK ;
  wire \DFF_185.D ;
  wire \DFF_185.Q ;
  wire \DFF_186.CK ;
  wire \DFF_186.D ;
  wire \DFF_186.Q ;
  wire \DFF_187.CK ;
  wire \DFF_187.D ;
  wire \DFF_187.Q ;
  wire \DFF_188.CK ;
  wire \DFF_188.D ;
  wire \DFF_188.Q ;
  wire \DFF_189.CK ;
  wire \DFF_189.D ;
  wire \DFF_189.Q ;
  wire \DFF_19.CK ;
  wire \DFF_19.D ;
  wire \DFF_19.Q ;
  wire \DFF_190.CK ;
  wire \DFF_190.D ;
  wire \DFF_190.Q ;
  wire \DFF_191.CK ;
  wire \DFF_191.D ;
  wire \DFF_191.Q ;
  wire \DFF_192.CK ;
  wire \DFF_192.D ;
  wire \DFF_192.Q ;
  wire \DFF_193.CK ;
  wire \DFF_193.D ;
  wire \DFF_193.Q ;
  wire \DFF_194.CK ;
  wire \DFF_194.D ;
  wire \DFF_194.Q ;
  wire \DFF_195.CK ;
  wire \DFF_195.D ;
  wire \DFF_195.Q ;
  wire \DFF_196.CK ;
  wire \DFF_196.D ;
  wire \DFF_196.Q ;
  wire \DFF_197.CK ;
  wire \DFF_197.D ;
  wire \DFF_197.Q ;
  wire \DFF_198.CK ;
  wire \DFF_198.D ;
  wire \DFF_198.Q ;
  wire \DFF_199.CK ;
  wire \DFF_199.D ;
  wire \DFF_199.Q ;
  wire \DFF_2.CK ;
  wire \DFF_2.D ;
  wire \DFF_2.Q ;
  wire \DFF_20.CK ;
  wire \DFF_20.D ;
  wire \DFF_20.Q ;
  wire \DFF_200.CK ;
  wire \DFF_200.D ;
  wire \DFF_200.Q ;
  wire \DFF_201.CK ;
  wire \DFF_201.D ;
  wire \DFF_201.Q ;
  wire \DFF_202.CK ;
  wire \DFF_202.D ;
  wire \DFF_202.Q ;
  wire \DFF_203.CK ;
  wire \DFF_203.D ;
  wire \DFF_203.Q ;
  wire \DFF_204.CK ;
  wire \DFF_204.D ;
  wire \DFF_204.Q ;
  wire \DFF_205.CK ;
  wire \DFF_205.D ;
  wire \DFF_205.Q ;
  wire \DFF_206.CK ;
  wire \DFF_206.D ;
  wire \DFF_206.Q ;
  wire \DFF_207.CK ;
  wire \DFF_207.D ;
  wire \DFF_207.Q ;
  wire \DFF_208.CK ;
  wire \DFF_208.D ;
  wire \DFF_208.Q ;
  wire \DFF_209.CK ;
  wire \DFF_209.D ;
  wire \DFF_209.Q ;
  wire \DFF_21.CK ;
  wire \DFF_21.D ;
  wire \DFF_21.Q ;
  wire \DFF_210.CK ;
  wire \DFF_210.D ;
  wire \DFF_210.Q ;
  wire \DFF_211.CK ;
  wire \DFF_211.D ;
  wire \DFF_211.Q ;
  wire \DFF_212.CK ;
  wire \DFF_212.D ;
  wire \DFF_212.Q ;
  wire \DFF_213.CK ;
  wire \DFF_213.D ;
  wire \DFF_213.Q ;
  wire \DFF_214.CK ;
  wire \DFF_214.D ;
  wire \DFF_214.Q ;
  wire \DFF_215.CK ;
  wire \DFF_215.D ;
  wire \DFF_215.Q ;
  wire \DFF_216.CK ;
  wire \DFF_216.D ;
  wire \DFF_216.Q ;
  wire \DFF_217.CK ;
  wire \DFF_217.D ;
  wire \DFF_217.Q ;
  wire \DFF_218.CK ;
  wire \DFF_218.D ;
  wire \DFF_218.Q ;
  wire \DFF_219.CK ;
  wire \DFF_219.D ;
  wire \DFF_219.Q ;
  wire \DFF_22.CK ;
  wire \DFF_22.D ;
  wire \DFF_22.Q ;
  wire \DFF_220.CK ;
  wire \DFF_220.D ;
  wire \DFF_220.Q ;
  wire \DFF_221.CK ;
  wire \DFF_221.D ;
  wire \DFF_221.Q ;
  wire \DFF_222.CK ;
  wire \DFF_222.D ;
  wire \DFF_222.Q ;
  wire \DFF_223.CK ;
  wire \DFF_223.D ;
  wire \DFF_223.Q ;
  wire \DFF_224.CK ;
  wire \DFF_224.D ;
  wire \DFF_224.Q ;
  wire \DFF_225.CK ;
  wire \DFF_225.D ;
  wire \DFF_225.Q ;
  wire \DFF_226.CK ;
  wire \DFF_226.D ;
  wire \DFF_226.Q ;
  wire \DFF_227.CK ;
  wire \DFF_227.D ;
  wire \DFF_227.Q ;
  wire \DFF_228.CK ;
  wire \DFF_228.D ;
  wire \DFF_228.Q ;
  wire \DFF_229.CK ;
  wire \DFF_229.D ;
  wire \DFF_229.Q ;
  wire \DFF_23.CK ;
  wire \DFF_23.D ;
  wire \DFF_23.Q ;
  wire \DFF_230.CK ;
  wire \DFF_230.D ;
  wire \DFF_230.Q ;
  wire \DFF_231.CK ;
  wire \DFF_231.D ;
  wire \DFF_231.Q ;
  wire \DFF_232.CK ;
  wire \DFF_232.D ;
  wire \DFF_232.Q ;
  wire \DFF_233.CK ;
  wire \DFF_233.D ;
  wire \DFF_233.Q ;
  wire \DFF_234.CK ;
  wire \DFF_234.D ;
  wire \DFF_234.Q ;
  wire \DFF_235.CK ;
  wire \DFF_235.D ;
  wire \DFF_235.Q ;
  wire \DFF_236.CK ;
  wire \DFF_236.D ;
  wire \DFF_236.Q ;
  wire \DFF_237.CK ;
  wire \DFF_237.D ;
  wire \DFF_237.Q ;
  wire \DFF_238.CK ;
  wire \DFF_238.D ;
  wire \DFF_238.Q ;
  wire \DFF_239.CK ;
  wire \DFF_239.D ;
  wire \DFF_239.Q ;
  wire \DFF_24.CK ;
  wire \DFF_24.D ;
  wire \DFF_24.Q ;
  wire \DFF_240.CK ;
  wire \DFF_240.D ;
  wire \DFF_240.Q ;
  wire \DFF_241.CK ;
  wire \DFF_241.D ;
  wire \DFF_241.Q ;
  wire \DFF_242.CK ;
  wire \DFF_242.D ;
  wire \DFF_242.Q ;
  wire \DFF_243.CK ;
  wire \DFF_243.D ;
  wire \DFF_243.Q ;
  wire \DFF_244.CK ;
  wire \DFF_244.D ;
  wire \DFF_244.Q ;
  wire \DFF_245.CK ;
  wire \DFF_245.D ;
  wire \DFF_245.Q ;
  wire \DFF_246.CK ;
  wire \DFF_246.D ;
  wire \DFF_246.Q ;
  wire \DFF_247.CK ;
  wire \DFF_247.D ;
  wire \DFF_247.Q ;
  wire \DFF_248.CK ;
  wire \DFF_248.D ;
  wire \DFF_248.Q ;
  wire \DFF_249.CK ;
  wire \DFF_249.D ;
  wire \DFF_249.Q ;
  wire \DFF_25.CK ;
  wire \DFF_25.D ;
  wire \DFF_25.Q ;
  wire \DFF_250.CK ;
  wire \DFF_250.D ;
  wire \DFF_250.Q ;
  wire \DFF_251.CK ;
  wire \DFF_251.D ;
  wire \DFF_251.Q ;
  wire \DFF_252.CK ;
  wire \DFF_252.D ;
  wire \DFF_252.Q ;
  wire \DFF_253.CK ;
  wire \DFF_253.D ;
  wire \DFF_253.Q ;
  wire \DFF_254.CK ;
  wire \DFF_254.D ;
  wire \DFF_254.Q ;
  wire \DFF_255.CK ;
  wire \DFF_255.D ;
  wire \DFF_255.Q ;
  wire \DFF_256.CK ;
  wire \DFF_256.D ;
  wire \DFF_256.Q ;
  wire \DFF_257.CK ;
  wire \DFF_257.D ;
  wire \DFF_257.Q ;
  wire \DFF_258.CK ;
  wire \DFF_258.D ;
  wire \DFF_258.Q ;
  wire \DFF_259.CK ;
  wire \DFF_259.D ;
  wire \DFF_259.Q ;
  wire \DFF_26.CK ;
  wire \DFF_26.D ;
  wire \DFF_26.Q ;
  wire \DFF_260.CK ;
  wire \DFF_260.D ;
  wire \DFF_260.Q ;
  wire \DFF_261.CK ;
  wire \DFF_261.D ;
  wire \DFF_261.Q ;
  wire \DFF_262.CK ;
  wire \DFF_262.D ;
  wire \DFF_262.Q ;
  wire \DFF_263.CK ;
  wire \DFF_263.D ;
  wire \DFF_263.Q ;
  wire \DFF_264.CK ;
  wire \DFF_264.D ;
  wire \DFF_264.Q ;
  wire \DFF_265.CK ;
  wire \DFF_265.D ;
  wire \DFF_265.Q ;
  wire \DFF_266.CK ;
  wire \DFF_266.D ;
  wire \DFF_266.Q ;
  wire \DFF_267.CK ;
  wire \DFF_267.D ;
  wire \DFF_267.Q ;
  wire \DFF_268.CK ;
  wire \DFF_268.D ;
  wire \DFF_268.Q ;
  wire \DFF_269.CK ;
  wire \DFF_269.D ;
  wire \DFF_269.Q ;
  wire \DFF_27.CK ;
  wire \DFF_27.D ;
  wire \DFF_27.Q ;
  wire \DFF_270.CK ;
  wire \DFF_270.D ;
  wire \DFF_270.Q ;
  wire \DFF_271.CK ;
  wire \DFF_271.D ;
  wire \DFF_271.Q ;
  wire \DFF_272.CK ;
  wire \DFF_272.D ;
  wire \DFF_272.Q ;
  wire \DFF_273.CK ;
  wire \DFF_273.D ;
  wire \DFF_273.Q ;
  wire \DFF_274.CK ;
  wire \DFF_274.D ;
  wire \DFF_274.Q ;
  wire \DFF_275.CK ;
  wire \DFF_275.D ;
  wire \DFF_275.Q ;
  wire \DFF_276.CK ;
  wire \DFF_276.D ;
  wire \DFF_276.Q ;
  wire \DFF_277.CK ;
  wire \DFF_277.D ;
  wire \DFF_277.Q ;
  wire \DFF_278.CK ;
  wire \DFF_278.D ;
  wire \DFF_278.Q ;
  wire \DFF_279.CK ;
  wire \DFF_279.D ;
  wire \DFF_279.Q ;
  wire \DFF_28.CK ;
  wire \DFF_28.D ;
  wire \DFF_28.Q ;
  wire \DFF_280.CK ;
  wire \DFF_280.D ;
  wire \DFF_280.Q ;
  wire \DFF_281.CK ;
  wire \DFF_281.D ;
  wire \DFF_281.Q ;
  wire \DFF_282.CK ;
  wire \DFF_282.D ;
  wire \DFF_282.Q ;
  wire \DFF_283.CK ;
  wire \DFF_283.D ;
  wire \DFF_283.Q ;
  wire \DFF_284.CK ;
  wire \DFF_284.D ;
  wire \DFF_284.Q ;
  wire \DFF_285.CK ;
  wire \DFF_285.D ;
  wire \DFF_285.Q ;
  wire \DFF_286.CK ;
  wire \DFF_286.D ;
  wire \DFF_286.Q ;
  wire \DFF_287.CK ;
  wire \DFF_287.D ;
  wire \DFF_287.Q ;
  wire \DFF_288.CK ;
  wire \DFF_288.D ;
  wire \DFF_288.Q ;
  wire \DFF_289.CK ;
  wire \DFF_289.D ;
  wire \DFF_289.Q ;
  wire \DFF_29.CK ;
  wire \DFF_29.D ;
  wire \DFF_29.Q ;
  wire \DFF_290.CK ;
  wire \DFF_290.D ;
  wire \DFF_290.Q ;
  wire \DFF_291.CK ;
  wire \DFF_291.D ;
  wire \DFF_291.Q ;
  wire \DFF_292.CK ;
  wire \DFF_292.D ;
  wire \DFF_292.Q ;
  wire \DFF_293.CK ;
  wire \DFF_293.D ;
  wire \DFF_293.Q ;
  wire \DFF_294.CK ;
  wire \DFF_294.D ;
  wire \DFF_294.Q ;
  wire \DFF_295.CK ;
  wire \DFF_295.D ;
  wire \DFF_295.Q ;
  wire \DFF_296.CK ;
  wire \DFF_296.D ;
  wire \DFF_296.Q ;
  wire \DFF_297.CK ;
  wire \DFF_297.D ;
  wire \DFF_297.Q ;
  wire \DFF_298.CK ;
  wire \DFF_298.D ;
  wire \DFF_298.Q ;
  wire \DFF_299.CK ;
  wire \DFF_299.D ;
  wire \DFF_299.Q ;
  wire \DFF_3.CK ;
  wire \DFF_3.D ;
  wire \DFF_3.Q ;
  wire \DFF_30.CK ;
  wire \DFF_30.D ;
  wire \DFF_30.Q ;
  wire \DFF_300.CK ;
  wire \DFF_300.D ;
  wire \DFF_300.Q ;
  wire \DFF_301.CK ;
  wire \DFF_301.D ;
  wire \DFF_301.Q ;
  wire \DFF_302.CK ;
  wire \DFF_302.D ;
  wire \DFF_302.Q ;
  wire \DFF_303.CK ;
  wire \DFF_303.D ;
  wire \DFF_303.Q ;
  wire \DFF_304.CK ;
  wire \DFF_304.D ;
  wire \DFF_304.Q ;
  wire \DFF_305.CK ;
  wire \DFF_305.D ;
  wire \DFF_305.Q ;
  wire \DFF_306.CK ;
  wire \DFF_306.D ;
  wire \DFF_306.Q ;
  wire \DFF_307.CK ;
  wire \DFF_307.D ;
  wire \DFF_307.Q ;
  wire \DFF_308.CK ;
  wire \DFF_308.D ;
  wire \DFF_308.Q ;
  wire \DFF_309.CK ;
  wire \DFF_309.D ;
  wire \DFF_309.Q ;
  wire \DFF_31.CK ;
  wire \DFF_31.D ;
  wire \DFF_31.Q ;
  wire \DFF_310.CK ;
  wire \DFF_310.D ;
  wire \DFF_310.Q ;
  wire \DFF_311.CK ;
  wire \DFF_311.D ;
  wire \DFF_311.Q ;
  wire \DFF_312.CK ;
  wire \DFF_312.D ;
  wire \DFF_312.Q ;
  wire \DFF_313.CK ;
  wire \DFF_313.D ;
  wire \DFF_313.Q ;
  wire \DFF_314.CK ;
  wire \DFF_314.D ;
  wire \DFF_314.Q ;
  wire \DFF_315.CK ;
  wire \DFF_315.D ;
  wire \DFF_315.Q ;
  wire \DFF_316.CK ;
  wire \DFF_316.D ;
  wire \DFF_316.Q ;
  wire \DFF_317.CK ;
  wire \DFF_317.D ;
  wire \DFF_317.Q ;
  wire \DFF_318.CK ;
  wire \DFF_319.CK ;
  wire \DFF_32.CK ;
  wire \DFF_32.D ;
  wire \DFF_32.Q ;
  wire \DFF_320.CK ;
  wire \DFF_321.CK ;
  wire \DFF_322.CK ;
  wire \DFF_323.CK ;
  wire \DFF_324.CK ;
  wire \DFF_325.CK ;
  wire \DFF_326.CK ;
  wire \DFF_327.CK ;
  wire \DFF_328.CK ;
  wire \DFF_328.D ;
  wire \DFF_328.Q ;
  wire \DFF_329.CK ;
  wire \DFF_329.D ;
  wire \DFF_329.Q ;
  wire \DFF_33.CK ;
  wire \DFF_33.D ;
  wire \DFF_33.Q ;
  wire \DFF_330.CK ;
  wire \DFF_330.D ;
  wire \DFF_330.Q ;
  wire \DFF_331.CK ;
  wire \DFF_331.D ;
  wire \DFF_331.Q ;
  wire \DFF_332.CK ;
  wire \DFF_332.D ;
  wire \DFF_332.Q ;
  wire \DFF_333.CK ;
  wire \DFF_333.D ;
  wire \DFF_333.Q ;
  wire \DFF_334.CK ;
  wire \DFF_334.D ;
  wire \DFF_334.Q ;
  wire \DFF_335.CK ;
  wire \DFF_335.D ;
  wire \DFF_335.Q ;
  wire \DFF_336.CK ;
  wire \DFF_336.D ;
  wire \DFF_336.Q ;
  wire \DFF_337.CK ;
  wire \DFF_337.D ;
  wire \DFF_337.Q ;
  wire \DFF_338.CK ;
  wire \DFF_338.D ;
  wire \DFF_338.Q ;
  wire \DFF_339.CK ;
  wire \DFF_339.D ;
  wire \DFF_339.Q ;
  wire \DFF_34.CK ;
  wire \DFF_34.D ;
  wire \DFF_34.Q ;
  wire \DFF_340.CK ;
  wire \DFF_340.D ;
  wire \DFF_340.Q ;
  wire \DFF_341.CK ;
  wire \DFF_341.D ;
  wire \DFF_341.Q ;
  wire \DFF_342.CK ;
  wire \DFF_342.D ;
  wire \DFF_342.Q ;
  wire \DFF_343.CK ;
  wire \DFF_343.D ;
  wire \DFF_343.Q ;
  wire \DFF_344.CK ;
  wire \DFF_344.D ;
  wire \DFF_344.Q ;
  wire \DFF_345.CK ;
  wire \DFF_345.D ;
  wire \DFF_345.Q ;
  wire \DFF_346.CK ;
  wire \DFF_346.D ;
  wire \DFF_346.Q ;
  wire \DFF_347.CK ;
  wire \DFF_347.D ;
  wire \DFF_347.Q ;
  wire \DFF_348.CK ;
  wire \DFF_348.D ;
  wire \DFF_348.Q ;
  wire \DFF_349.CK ;
  wire \DFF_349.D ;
  wire \DFF_349.Q ;
  wire \DFF_35.CK ;
  wire \DFF_35.D ;
  wire \DFF_35.Q ;
  wire \DFF_350.CK ;
  wire \DFF_350.D ;
  wire \DFF_350.Q ;
  wire \DFF_351.CK ;
  wire \DFF_351.D ;
  wire \DFF_351.Q ;
  wire \DFF_352.CK ;
  wire \DFF_352.D ;
  wire \DFF_352.Q ;
  wire \DFF_353.CK ;
  wire \DFF_353.D ;
  wire \DFF_353.Q ;
  wire \DFF_354.CK ;
  wire \DFF_354.D ;
  wire \DFF_354.Q ;
  wire \DFF_355.CK ;
  wire \DFF_355.D ;
  wire \DFF_355.Q ;
  wire \DFF_356.CK ;
  wire \DFF_356.D ;
  wire \DFF_356.Q ;
  wire \DFF_357.CK ;
  wire \DFF_357.D ;
  wire \DFF_357.Q ;
  wire \DFF_358.CK ;
  wire \DFF_358.D ;
  wire \DFF_358.Q ;
  wire \DFF_359.CK ;
  wire \DFF_359.D ;
  wire \DFF_359.Q ;
  wire \DFF_36.CK ;
  wire \DFF_36.D ;
  wire \DFF_36.Q ;
  wire \DFF_360.CK ;
  wire \DFF_360.D ;
  wire \DFF_360.Q ;
  wire \DFF_361.CK ;
  wire \DFF_361.D ;
  wire \DFF_361.Q ;
  wire \DFF_362.CK ;
  wire \DFF_362.D ;
  wire \DFF_362.Q ;
  wire \DFF_363.CK ;
  wire \DFF_363.D ;
  wire \DFF_363.Q ;
  wire \DFF_364.CK ;
  wire \DFF_364.D ;
  wire \DFF_364.Q ;
  wire \DFF_365.CK ;
  wire \DFF_365.D ;
  wire \DFF_365.Q ;
  wire \DFF_366.CK ;
  wire \DFF_366.D ;
  wire \DFF_366.Q ;
  wire \DFF_367.CK ;
  wire \DFF_367.D ;
  wire \DFF_367.Q ;
  wire \DFF_368.CK ;
  wire \DFF_368.D ;
  wire \DFF_368.Q ;
  wire \DFF_369.CK ;
  wire \DFF_369.D ;
  wire \DFF_369.Q ;
  wire \DFF_37.CK ;
  wire \DFF_37.D ;
  wire \DFF_37.Q ;
  wire \DFF_370.CK ;
  wire \DFF_370.D ;
  wire \DFF_370.Q ;
  wire \DFF_371.CK ;
  wire \DFF_371.D ;
  wire \DFF_371.Q ;
  wire \DFF_372.CK ;
  wire \DFF_372.D ;
  wire \DFF_372.Q ;
  wire \DFF_373.CK ;
  wire \DFF_373.D ;
  wire \DFF_373.Q ;
  wire \DFF_374.CK ;
  wire \DFF_374.D ;
  wire \DFF_374.Q ;
  wire \DFF_375.CK ;
  wire \DFF_375.D ;
  wire \DFF_375.Q ;
  wire \DFF_376.CK ;
  wire \DFF_376.D ;
  wire \DFF_376.Q ;
  wire \DFF_377.CK ;
  wire \DFF_377.D ;
  wire \DFF_377.Q ;
  wire \DFF_378.CK ;
  wire \DFF_378.D ;
  wire \DFF_378.Q ;
  wire \DFF_379.CK ;
  wire \DFF_379.D ;
  wire \DFF_379.Q ;
  wire \DFF_38.CK ;
  wire \DFF_38.D ;
  wire \DFF_38.Q ;
  wire \DFF_380.CK ;
  wire \DFF_380.D ;
  wire \DFF_380.Q ;
  wire \DFF_381.CK ;
  wire \DFF_381.D ;
  wire \DFF_381.Q ;
  wire \DFF_382.CK ;
  wire \DFF_382.D ;
  wire \DFF_382.Q ;
  wire \DFF_383.CK ;
  wire \DFF_383.D ;
  wire \DFF_383.Q ;
  wire \DFF_384.CK ;
  wire \DFF_384.D ;
  wire \DFF_384.Q ;
  wire \DFF_385.CK ;
  wire \DFF_385.D ;
  wire \DFF_385.Q ;
  wire \DFF_386.CK ;
  wire \DFF_386.D ;
  wire \DFF_386.Q ;
  wire \DFF_387.CK ;
  wire \DFF_387.D ;
  wire \DFF_387.Q ;
  wire \DFF_388.CK ;
  wire \DFF_388.D ;
  wire \DFF_388.Q ;
  wire \DFF_389.CK ;
  wire \DFF_389.D ;
  wire \DFF_389.Q ;
  wire \DFF_39.CK ;
  wire \DFF_39.D ;
  wire \DFF_39.Q ;
  wire \DFF_390.CK ;
  wire \DFF_390.D ;
  wire \DFF_390.Q ;
  wire \DFF_391.CK ;
  wire \DFF_391.D ;
  wire \DFF_391.Q ;
  wire \DFF_392.CK ;
  wire \DFF_392.D ;
  wire \DFF_392.Q ;
  wire \DFF_393.CK ;
  wire \DFF_393.D ;
  wire \DFF_393.Q ;
  wire \DFF_394.CK ;
  wire \DFF_394.D ;
  wire \DFF_394.Q ;
  wire \DFF_395.CK ;
  wire \DFF_395.D ;
  wire \DFF_395.Q ;
  wire \DFF_396.CK ;
  wire \DFF_396.D ;
  wire \DFF_396.Q ;
  wire \DFF_397.CK ;
  wire \DFF_397.D ;
  wire \DFF_397.Q ;
  wire \DFF_398.CK ;
  wire \DFF_398.D ;
  wire \DFF_398.Q ;
  wire \DFF_399.CK ;
  wire \DFF_399.D ;
  wire \DFF_399.Q ;
  wire \DFF_4.CK ;
  wire \DFF_4.D ;
  wire \DFF_4.Q ;
  wire \DFF_40.CK ;
  wire \DFF_40.D ;
  wire \DFF_40.Q ;
  wire \DFF_400.CK ;
  wire \DFF_400.D ;
  wire \DFF_400.Q ;
  wire \DFF_401.CK ;
  wire \DFF_401.D ;
  wire \DFF_401.Q ;
  wire \DFF_402.CK ;
  wire \DFF_402.D ;
  wire \DFF_402.Q ;
  wire \DFF_403.CK ;
  wire \DFF_403.D ;
  wire \DFF_403.Q ;
  wire \DFF_404.CK ;
  wire \DFF_404.D ;
  wire \DFF_404.Q ;
  wire \DFF_405.CK ;
  wire \DFF_405.D ;
  wire \DFF_405.Q ;
  wire \DFF_406.CK ;
  wire \DFF_406.D ;
  wire \DFF_406.Q ;
  wire \DFF_407.CK ;
  wire \DFF_407.D ;
  wire \DFF_407.Q ;
  wire \DFF_408.CK ;
  wire \DFF_408.D ;
  wire \DFF_408.Q ;
  wire \DFF_409.CK ;
  wire \DFF_409.D ;
  wire \DFF_409.Q ;
  wire \DFF_41.CK ;
  wire \DFF_41.D ;
  wire \DFF_41.Q ;
  wire \DFF_410.CK ;
  wire \DFF_410.D ;
  wire \DFF_410.Q ;
  wire \DFF_411.CK ;
  wire \DFF_411.D ;
  wire \DFF_411.Q ;
  wire \DFF_412.CK ;
  wire \DFF_412.D ;
  wire \DFF_412.Q ;
  wire \DFF_413.CK ;
  wire \DFF_413.D ;
  wire \DFF_413.Q ;
  wire \DFF_414.CK ;
  wire \DFF_414.D ;
  wire \DFF_414.Q ;
  wire \DFF_415.CK ;
  wire \DFF_415.D ;
  wire \DFF_415.Q ;
  wire \DFF_416.CK ;
  wire \DFF_416.D ;
  wire \DFF_416.Q ;
  wire \DFF_417.CK ;
  wire \DFF_417.D ;
  wire \DFF_417.Q ;
  wire \DFF_418.CK ;
  wire \DFF_418.D ;
  wire \DFF_418.Q ;
  wire \DFF_419.CK ;
  wire \DFF_419.D ;
  wire \DFF_419.Q ;
  wire \DFF_42.CK ;
  wire \DFF_42.D ;
  wire \DFF_42.Q ;
  wire \DFF_420.CK ;
  wire \DFF_420.D ;
  wire \DFF_420.Q ;
  wire \DFF_421.CK ;
  wire \DFF_421.D ;
  wire \DFF_421.Q ;
  wire \DFF_422.CK ;
  wire \DFF_422.D ;
  wire \DFF_422.Q ;
  wire \DFF_423.CK ;
  wire \DFF_423.D ;
  wire \DFF_423.Q ;
  wire \DFF_424.CK ;
  wire \DFF_424.D ;
  wire \DFF_424.Q ;
  wire \DFF_425.CK ;
  wire \DFF_425.D ;
  wire \DFF_425.Q ;
  wire \DFF_426.CK ;
  wire \DFF_426.D ;
  wire \DFF_426.Q ;
  wire \DFF_427.CK ;
  wire \DFF_427.D ;
  wire \DFF_427.Q ;
  wire \DFF_428.CK ;
  wire \DFF_428.D ;
  wire \DFF_428.Q ;
  wire \DFF_429.CK ;
  wire \DFF_429.D ;
  wire \DFF_429.Q ;
  wire \DFF_43.CK ;
  wire \DFF_43.D ;
  wire \DFF_43.Q ;
  wire \DFF_430.CK ;
  wire \DFF_430.D ;
  wire \DFF_430.Q ;
  wire \DFF_431.CK ;
  wire \DFF_431.D ;
  wire \DFF_431.Q ;
  wire \DFF_432.CK ;
  wire \DFF_432.D ;
  wire \DFF_432.Q ;
  wire \DFF_433.CK ;
  wire \DFF_433.D ;
  wire \DFF_433.Q ;
  wire \DFF_434.CK ;
  wire \DFF_435.CK ;
  wire \DFF_436.CK ;
  wire \DFF_437.CK ;
  wire \DFF_438.CK ;
  wire \DFF_439.CK ;
  wire \DFF_44.CK ;
  wire \DFF_44.D ;
  wire \DFF_44.Q ;
  wire \DFF_440.CK ;
  wire \DFF_441.CK ;
  wire \DFF_442.CK ;
  wire \DFF_442.D ;
  wire \DFF_442.Q ;
  wire \DFF_443.CK ;
  wire \DFF_443.D ;
  wire \DFF_443.Q ;
  wire \DFF_444.CK ;
  wire \DFF_444.D ;
  wire \DFF_444.Q ;
  wire \DFF_445.CK ;
  wire \DFF_445.D ;
  wire \DFF_445.Q ;
  wire \DFF_446.CK ;
  wire \DFF_446.D ;
  wire \DFF_446.Q ;
  wire \DFF_447.CK ;
  wire \DFF_447.D ;
  wire \DFF_447.Q ;
  wire \DFF_448.CK ;
  wire \DFF_448.D ;
  wire \DFF_448.Q ;
  wire \DFF_449.CK ;
  wire \DFF_449.D ;
  wire \DFF_449.Q ;
  wire \DFF_45.CK ;
  wire \DFF_45.D ;
  wire \DFF_45.Q ;
  wire \DFF_450.CK ;
  wire \DFF_450.D ;
  wire \DFF_450.Q ;
  wire \DFF_451.CK ;
  wire \DFF_451.D ;
  wire \DFF_451.Q ;
  wire \DFF_452.CK ;
  wire \DFF_452.D ;
  wire \DFF_452.Q ;
  wire \DFF_453.CK ;
  wire \DFF_453.D ;
  wire \DFF_453.Q ;
  wire \DFF_454.CK ;
  wire \DFF_454.D ;
  wire \DFF_454.Q ;
  wire \DFF_455.CK ;
  wire \DFF_455.D ;
  wire \DFF_455.Q ;
  wire \DFF_456.CK ;
  wire \DFF_456.D ;
  wire \DFF_456.Q ;
  wire \DFF_457.CK ;
  wire \DFF_457.D ;
  wire \DFF_457.Q ;
  wire \DFF_458.CK ;
  wire \DFF_458.D ;
  wire \DFF_458.Q ;
  wire \DFF_459.CK ;
  wire \DFF_459.D ;
  wire \DFF_459.Q ;
  wire \DFF_46.CK ;
  wire \DFF_46.D ;
  wire \DFF_46.Q ;
  wire \DFF_460.CK ;
  wire \DFF_460.D ;
  wire \DFF_460.Q ;
  wire \DFF_461.CK ;
  wire \DFF_461.D ;
  wire \DFF_461.Q ;
  wire \DFF_462.CK ;
  wire \DFF_462.D ;
  wire \DFF_462.Q ;
  wire \DFF_463.CK ;
  wire \DFF_463.D ;
  wire \DFF_463.Q ;
  wire \DFF_464.CK ;
  wire \DFF_464.D ;
  wire \DFF_464.Q ;
  wire \DFF_465.CK ;
  wire \DFF_465.D ;
  wire \DFF_465.Q ;
  wire \DFF_466.CK ;
  wire \DFF_466.D ;
  wire \DFF_466.Q ;
  wire \DFF_467.CK ;
  wire \DFF_467.D ;
  wire \DFF_467.Q ;
  wire \DFF_468.CK ;
  wire \DFF_468.D ;
  wire \DFF_468.Q ;
  wire \DFF_469.CK ;
  wire \DFF_469.D ;
  wire \DFF_469.Q ;
  wire \DFF_47.CK ;
  wire \DFF_47.D ;
  wire \DFF_47.Q ;
  wire \DFF_470.CK ;
  wire \DFF_470.D ;
  wire \DFF_470.Q ;
  wire \DFF_471.CK ;
  wire \DFF_471.D ;
  wire \DFF_471.Q ;
  wire \DFF_472.CK ;
  wire \DFF_472.D ;
  wire \DFF_472.Q ;
  wire \DFF_473.CK ;
  wire \DFF_473.D ;
  wire \DFF_473.Q ;
  wire \DFF_474.CK ;
  wire \DFF_474.D ;
  wire \DFF_474.Q ;
  wire \DFF_475.CK ;
  wire \DFF_475.D ;
  wire \DFF_475.Q ;
  wire \DFF_476.CK ;
  wire \DFF_476.D ;
  wire \DFF_476.Q ;
  wire \DFF_477.CK ;
  wire \DFF_477.D ;
  wire \DFF_477.Q ;
  wire \DFF_478.CK ;
  wire \DFF_478.D ;
  wire \DFF_478.Q ;
  wire \DFF_479.CK ;
  wire \DFF_479.D ;
  wire \DFF_479.Q ;
  wire \DFF_48.CK ;
  wire \DFF_48.D ;
  wire \DFF_48.Q ;
  wire \DFF_480.CK ;
  wire \DFF_480.D ;
  wire \DFF_480.Q ;
  wire \DFF_481.CK ;
  wire \DFF_481.D ;
  wire \DFF_481.Q ;
  wire \DFF_482.CK ;
  wire \DFF_482.D ;
  wire \DFF_482.Q ;
  wire \DFF_483.CK ;
  wire \DFF_483.D ;
  wire \DFF_483.Q ;
  wire \DFF_484.CK ;
  wire \DFF_484.D ;
  wire \DFF_484.Q ;
  wire \DFF_485.CK ;
  wire \DFF_485.D ;
  wire \DFF_485.Q ;
  wire \DFF_486.CK ;
  wire \DFF_486.D ;
  wire \DFF_486.Q ;
  wire \DFF_487.CK ;
  wire \DFF_487.D ;
  wire \DFF_487.Q ;
  wire \DFF_488.CK ;
  wire \DFF_488.D ;
  wire \DFF_488.Q ;
  wire \DFF_489.CK ;
  wire \DFF_489.D ;
  wire \DFF_489.Q ;
  wire \DFF_49.CK ;
  wire \DFF_49.D ;
  wire \DFF_49.Q ;
  wire \DFF_490.CK ;
  wire \DFF_490.D ;
  wire \DFF_490.Q ;
  wire \DFF_491.CK ;
  wire \DFF_491.D ;
  wire \DFF_491.Q ;
  wire \DFF_492.CK ;
  wire \DFF_492.D ;
  wire \DFF_492.Q ;
  wire \DFF_493.CK ;
  wire \DFF_493.D ;
  wire \DFF_493.Q ;
  wire \DFF_494.CK ;
  wire \DFF_494.D ;
  wire \DFF_494.Q ;
  wire \DFF_495.CK ;
  wire \DFF_495.D ;
  wire \DFF_495.Q ;
  wire \DFF_496.CK ;
  wire \DFF_496.D ;
  wire \DFF_496.Q ;
  wire \DFF_497.CK ;
  wire \DFF_497.D ;
  wire \DFF_497.Q ;
  wire \DFF_498.CK ;
  wire \DFF_498.D ;
  wire \DFF_498.Q ;
  wire \DFF_499.CK ;
  wire \DFF_499.D ;
  wire \DFF_499.Q ;
  wire \DFF_5.CK ;
  wire \DFF_5.D ;
  wire \DFF_5.Q ;
  wire \DFF_50.CK ;
  wire \DFF_50.D ;
  wire \DFF_50.Q ;
  wire \DFF_500.CK ;
  wire \DFF_500.D ;
  wire \DFF_500.Q ;
  wire \DFF_501.CK ;
  wire \DFF_501.D ;
  wire \DFF_501.Q ;
  wire \DFF_502.CK ;
  wire \DFF_502.D ;
  wire \DFF_502.Q ;
  wire \DFF_503.CK ;
  wire \DFF_503.D ;
  wire \DFF_503.Q ;
  wire \DFF_504.CK ;
  wire \DFF_504.D ;
  wire \DFF_504.Q ;
  wire \DFF_505.CK ;
  wire \DFF_505.D ;
  wire \DFF_505.Q ;
  wire \DFF_506.CK ;
  wire \DFF_506.D ;
  wire \DFF_506.Q ;
  wire \DFF_507.CK ;
  wire \DFF_507.D ;
  wire \DFF_507.Q ;
  wire \DFF_508.CK ;
  wire \DFF_508.D ;
  wire \DFF_508.Q ;
  wire \DFF_509.CK ;
  wire \DFF_509.D ;
  wire \DFF_509.Q ;
  wire \DFF_51.CK ;
  wire \DFF_51.D ;
  wire \DFF_51.Q ;
  wire \DFF_510.CK ;
  wire \DFF_510.D ;
  wire \DFF_510.Q ;
  wire \DFF_511.CK ;
  wire \DFF_511.D ;
  wire \DFF_511.Q ;
  wire \DFF_512.CK ;
  wire \DFF_512.D ;
  wire \DFF_512.Q ;
  wire \DFF_513.CK ;
  wire \DFF_513.D ;
  wire \DFF_513.Q ;
  wire \DFF_514.CK ;
  wire \DFF_514.D ;
  wire \DFF_514.Q ;
  wire \DFF_515.CK ;
  wire \DFF_515.D ;
  wire \DFF_515.Q ;
  wire \DFF_516.CK ;
  wire \DFF_516.D ;
  wire \DFF_516.Q ;
  wire \DFF_517.CK ;
  wire \DFF_517.D ;
  wire \DFF_517.Q ;
  wire \DFF_518.CK ;
  wire \DFF_518.D ;
  wire \DFF_518.Q ;
  wire \DFF_519.CK ;
  wire \DFF_519.D ;
  wire \DFF_519.Q ;
  wire \DFF_52.CK ;
  wire \DFF_52.D ;
  wire \DFF_52.Q ;
  wire \DFF_520.CK ;
  wire \DFF_520.D ;
  wire \DFF_520.Q ;
  wire \DFF_521.CK ;
  wire \DFF_521.D ;
  wire \DFF_521.Q ;
  wire \DFF_522.CK ;
  wire \DFF_522.D ;
  wire \DFF_522.Q ;
  wire \DFF_523.CK ;
  wire \DFF_523.D ;
  wire \DFF_523.Q ;
  wire \DFF_524.CK ;
  wire \DFF_524.D ;
  wire \DFF_524.Q ;
  wire \DFF_525.CK ;
  wire \DFF_525.D ;
  wire \DFF_525.Q ;
  wire \DFF_526.CK ;
  wire \DFF_526.D ;
  wire \DFF_526.Q ;
  wire \DFF_527.CK ;
  wire \DFF_527.D ;
  wire \DFF_527.Q ;
  wire \DFF_528.CK ;
  wire \DFF_528.D ;
  wire \DFF_528.Q ;
  wire \DFF_529.CK ;
  wire \DFF_529.D ;
  wire \DFF_529.Q ;
  wire \DFF_53.CK ;
  wire \DFF_53.D ;
  wire \DFF_53.Q ;
  wire \DFF_530.CK ;
  wire \DFF_530.D ;
  wire \DFF_530.Q ;
  wire \DFF_531.CK ;
  wire \DFF_531.D ;
  wire \DFF_531.Q ;
  wire \DFF_532.CK ;
  wire \DFF_532.D ;
  wire \DFF_532.Q ;
  wire \DFF_533.CK ;
  wire \DFF_533.D ;
  wire \DFF_533.Q ;
  wire \DFF_534.CK ;
  wire \DFF_534.D ;
  wire \DFF_534.Q ;
  wire \DFF_535.CK ;
  wire \DFF_535.D ;
  wire \DFF_535.Q ;
  wire \DFF_536.CK ;
  wire \DFF_536.D ;
  wire \DFF_536.Q ;
  wire \DFF_537.CK ;
  wire \DFF_537.D ;
  wire \DFF_537.Q ;
  wire \DFF_538.CK ;
  wire \DFF_538.D ;
  wire \DFF_538.Q ;
  wire \DFF_539.CK ;
  wire \DFF_539.D ;
  wire \DFF_539.Q ;
  wire \DFF_54.CK ;
  wire \DFF_54.D ;
  wire \DFF_54.Q ;
  wire \DFF_540.CK ;
  wire \DFF_540.D ;
  wire \DFF_540.Q ;
  wire \DFF_541.CK ;
  wire \DFF_541.D ;
  wire \DFF_541.Q ;
  wire \DFF_542.CK ;
  wire \DFF_542.D ;
  wire \DFF_542.Q ;
  wire \DFF_543.CK ;
  wire \DFF_543.D ;
  wire \DFF_543.Q ;
  wire \DFF_544.CK ;
  wire \DFF_544.D ;
  wire \DFF_544.Q ;
  wire \DFF_545.CK ;
  wire \DFF_545.D ;
  wire \DFF_545.Q ;
  wire \DFF_546.CK ;
  wire \DFF_546.D ;
  wire \DFF_546.Q ;
  wire \DFF_547.CK ;
  wire \DFF_547.D ;
  wire \DFF_547.Q ;
  wire \DFF_548.CK ;
  wire \DFF_548.D ;
  wire \DFF_548.Q ;
  wire \DFF_549.CK ;
  wire \DFF_549.D ;
  wire \DFF_549.Q ;
  wire \DFF_55.CK ;
  wire \DFF_55.D ;
  wire \DFF_55.Q ;
  wire \DFF_550.CK ;
  wire \DFF_550.D ;
  wire \DFF_550.Q ;
  wire \DFF_551.CK ;
  wire \DFF_551.D ;
  wire \DFF_551.Q ;
  wire \DFF_552.CK ;
  wire \DFF_552.D ;
  wire \DFF_552.Q ;
  wire \DFF_553.CK ;
  wire \DFF_553.D ;
  wire \DFF_553.Q ;
  wire \DFF_554.CK ;
  wire \DFF_554.D ;
  wire \DFF_554.Q ;
  wire \DFF_555.CK ;
  wire \DFF_555.D ;
  wire \DFF_555.Q ;
  wire \DFF_556.CK ;
  wire \DFF_556.D ;
  wire \DFF_556.Q ;
  wire \DFF_557.CK ;
  wire \DFF_557.D ;
  wire \DFF_557.Q ;
  wire \DFF_558.CK ;
  wire \DFF_558.D ;
  wire \DFF_558.Q ;
  wire \DFF_559.CK ;
  wire \DFF_559.D ;
  wire \DFF_559.Q ;
  wire \DFF_56.CK ;
  wire \DFF_56.D ;
  wire \DFF_56.Q ;
  wire \DFF_560.CK ;
  wire \DFF_560.D ;
  wire \DFF_560.Q ;
  wire \DFF_561.CK ;
  wire \DFF_561.D ;
  wire \DFF_561.Q ;
  wire \DFF_562.CK ;
  wire \DFF_562.D ;
  wire \DFF_562.Q ;
  wire \DFF_563.CK ;
  wire \DFF_563.D ;
  wire \DFF_563.Q ;
  wire \DFF_564.CK ;
  wire \DFF_564.D ;
  wire \DFF_564.Q ;
  wire \DFF_565.CK ;
  wire \DFF_565.D ;
  wire \DFF_565.Q ;
  wire \DFF_566.CK ;
  wire \DFF_566.D ;
  wire \DFF_566.Q ;
  wire \DFF_567.CK ;
  wire \DFF_567.D ;
  wire \DFF_567.Q ;
  wire \DFF_568.CK ;
  wire \DFF_568.D ;
  wire \DFF_568.Q ;
  wire \DFF_569.CK ;
  wire \DFF_569.D ;
  wire \DFF_569.Q ;
  wire \DFF_57.CK ;
  wire \DFF_57.D ;
  wire \DFF_57.Q ;
  wire \DFF_570.CK ;
  wire \DFF_570.D ;
  wire \DFF_570.Q ;
  wire \DFF_571.CK ;
  wire \DFF_571.D ;
  wire \DFF_571.Q ;
  wire \DFF_572.CK ;
  wire \DFF_572.D ;
  wire \DFF_572.Q ;
  wire \DFF_573.CK ;
  wire \DFF_573.D ;
  wire \DFF_573.Q ;
  wire \DFF_574.CK ;
  wire \DFF_574.D ;
  wire \DFF_574.Q ;
  wire \DFF_575.CK ;
  wire \DFF_575.D ;
  wire \DFF_575.Q ;
  wire \DFF_576.CK ;
  wire \DFF_576.D ;
  wire \DFF_576.Q ;
  wire \DFF_577.CK ;
  wire \DFF_577.D ;
  wire \DFF_577.Q ;
  wire \DFF_578.CK ;
  wire \DFF_578.D ;
  wire \DFF_578.Q ;
  wire \DFF_579.CK ;
  wire \DFF_579.D ;
  wire \DFF_579.Q ;
  wire \DFF_58.CK ;
  wire \DFF_58.D ;
  wire \DFF_58.Q ;
  wire \DFF_580.CK ;
  wire \DFF_580.D ;
  wire \DFF_580.Q ;
  wire \DFF_581.CK ;
  wire \DFF_581.D ;
  wire \DFF_581.Q ;
  wire \DFF_582.CK ;
  wire \DFF_582.D ;
  wire \DFF_582.Q ;
  wire \DFF_583.CK ;
  wire \DFF_583.D ;
  wire \DFF_583.Q ;
  wire \DFF_584.CK ;
  wire \DFF_584.D ;
  wire \DFF_584.Q ;
  wire \DFF_585.CK ;
  wire \DFF_585.D ;
  wire \DFF_585.Q ;
  wire \DFF_586.CK ;
  wire \DFF_586.D ;
  wire \DFF_586.Q ;
  wire \DFF_587.CK ;
  wire \DFF_587.D ;
  wire \DFF_587.Q ;
  wire \DFF_588.CK ;
  wire \DFF_588.D ;
  wire \DFF_588.Q ;
  wire \DFF_589.CK ;
  wire \DFF_589.D ;
  wire \DFF_589.Q ;
  wire \DFF_59.CK ;
  wire \DFF_59.D ;
  wire \DFF_59.Q ;
  wire \DFF_590.CK ;
  wire \DFF_590.D ;
  wire \DFF_590.Q ;
  wire \DFF_591.CK ;
  wire \DFF_591.D ;
  wire \DFF_591.Q ;
  wire \DFF_592.CK ;
  wire \DFF_592.D ;
  wire \DFF_592.Q ;
  wire \DFF_593.CK ;
  wire \DFF_593.D ;
  wire \DFF_593.Q ;
  wire \DFF_594.CK ;
  wire \DFF_594.D ;
  wire \DFF_594.Q ;
  wire \DFF_595.CK ;
  wire \DFF_595.D ;
  wire \DFF_595.Q ;
  wire \DFF_596.CK ;
  wire \DFF_596.D ;
  wire \DFF_596.Q ;
  wire \DFF_597.CK ;
  wire \DFF_597.D ;
  wire \DFF_597.Q ;
  wire \DFF_598.CK ;
  wire \DFF_598.D ;
  wire \DFF_598.Q ;
  wire \DFF_599.CK ;
  wire \DFF_599.D ;
  wire \DFF_599.Q ;
  wire \DFF_6.CK ;
  wire \DFF_6.D ;
  wire \DFF_6.Q ;
  wire \DFF_60.CK ;
  wire \DFF_60.D ;
  wire \DFF_60.Q ;
  wire \DFF_600.CK ;
  wire \DFF_600.D ;
  wire \DFF_600.Q ;
  wire \DFF_601.CK ;
  wire \DFF_601.D ;
  wire \DFF_601.Q ;
  wire \DFF_602.CK ;
  wire \DFF_602.D ;
  wire \DFF_602.Q ;
  wire \DFF_603.CK ;
  wire \DFF_603.D ;
  wire \DFF_603.Q ;
  wire \DFF_604.CK ;
  wire \DFF_604.D ;
  wire \DFF_604.Q ;
  wire \DFF_605.CK ;
  wire \DFF_605.D ;
  wire \DFF_605.Q ;
  wire \DFF_606.CK ;
  wire \DFF_606.D ;
  wire \DFF_606.Q ;
  wire \DFF_607.CK ;
  wire \DFF_607.D ;
  wire \DFF_607.Q ;
  wire \DFF_608.CK ;
  wire \DFF_608.D ;
  wire \DFF_608.Q ;
  wire \DFF_609.CK ;
  wire \DFF_609.D ;
  wire \DFF_609.Q ;
  wire \DFF_61.CK ;
  wire \DFF_61.D ;
  wire \DFF_61.Q ;
  wire \DFF_610.CK ;
  wire \DFF_610.D ;
  wire \DFF_610.Q ;
  wire \DFF_611.CK ;
  wire \DFF_611.D ;
  wire \DFF_611.Q ;
  wire \DFF_612.CK ;
  wire \DFF_612.D ;
  wire \DFF_612.Q ;
  wire \DFF_613.CK ;
  wire \DFF_613.D ;
  wire \DFF_613.Q ;
  wire \DFF_614.CK ;
  wire \DFF_614.D ;
  wire \DFF_614.Q ;
  wire \DFF_615.CK ;
  wire \DFF_615.D ;
  wire \DFF_615.Q ;
  wire \DFF_616.CK ;
  wire \DFF_616.D ;
  wire \DFF_616.Q ;
  wire \DFF_617.CK ;
  wire \DFF_617.D ;
  wire \DFF_617.Q ;
  wire \DFF_618.CK ;
  wire \DFF_618.D ;
  wire \DFF_618.Q ;
  wire \DFF_619.CK ;
  wire \DFF_619.D ;
  wire \DFF_619.Q ;
  wire \DFF_62.CK ;
  wire \DFF_62.D ;
  wire \DFF_62.Q ;
  wire \DFF_620.CK ;
  wire \DFF_620.D ;
  wire \DFF_620.Q ;
  wire \DFF_621.CK ;
  wire \DFF_621.D ;
  wire \DFF_621.Q ;
  wire \DFF_622.CK ;
  wire \DFF_622.D ;
  wire \DFF_622.Q ;
  wire \DFF_623.CK ;
  wire \DFF_623.D ;
  wire \DFF_623.Q ;
  wire \DFF_624.CK ;
  wire \DFF_624.D ;
  wire \DFF_624.Q ;
  wire \DFF_625.CK ;
  wire \DFF_625.D ;
  wire \DFF_625.Q ;
  wire \DFF_626.CK ;
  wire \DFF_626.D ;
  wire \DFF_626.Q ;
  wire \DFF_627.CK ;
  wire \DFF_627.D ;
  wire \DFF_627.Q ;
  wire \DFF_628.CK ;
  wire \DFF_628.D ;
  wire \DFF_628.Q ;
  wire \DFF_629.CK ;
  wire \DFF_629.D ;
  wire \DFF_629.Q ;
  wire \DFF_63.CK ;
  wire \DFF_63.D ;
  wire \DFF_63.Q ;
  wire \DFF_630.CK ;
  wire \DFF_630.D ;
  wire \DFF_630.Q ;
  wire \DFF_631.CK ;
  wire \DFF_631.D ;
  wire \DFF_631.Q ;
  wire \DFF_632.CK ;
  wire \DFF_632.D ;
  wire \DFF_632.Q ;
  wire \DFF_633.CK ;
  wire \DFF_633.D ;
  wire \DFF_633.Q ;
  wire \DFF_634.CK ;
  wire \DFF_634.D ;
  wire \DFF_634.Q ;
  wire \DFF_635.CK ;
  wire \DFF_635.D ;
  wire \DFF_635.Q ;
  wire \DFF_636.CK ;
  wire \DFF_636.D ;
  wire \DFF_636.Q ;
  wire \DFF_637.CK ;
  wire \DFF_637.D ;
  wire \DFF_637.Q ;
  wire \DFF_638.CK ;
  wire \DFF_638.D ;
  wire \DFF_638.Q ;
  wire \DFF_639.CK ;
  wire \DFF_639.D ;
  wire \DFF_639.Q ;
  wire \DFF_64.CK ;
  wire \DFF_64.D ;
  wire \DFF_64.Q ;
  wire \DFF_640.CK ;
  wire \DFF_640.D ;
  wire \DFF_640.Q ;
  wire \DFF_641.CK ;
  wire \DFF_641.D ;
  wire \DFF_641.Q ;
  wire \DFF_642.CK ;
  wire \DFF_642.D ;
  wire \DFF_642.Q ;
  wire \DFF_643.CK ;
  wire \DFF_643.D ;
  wire \DFF_643.Q ;
  wire \DFF_644.CK ;
  wire \DFF_644.D ;
  wire \DFF_644.Q ;
  wire \DFF_645.CK ;
  wire \DFF_645.D ;
  wire \DFF_645.Q ;
  wire \DFF_646.CK ;
  wire \DFF_646.D ;
  wire \DFF_646.Q ;
  wire \DFF_647.CK ;
  wire \DFF_647.D ;
  wire \DFF_647.Q ;
  wire \DFF_648.CK ;
  wire \DFF_648.D ;
  wire \DFF_648.Q ;
  wire \DFF_649.CK ;
  wire \DFF_649.D ;
  wire \DFF_649.Q ;
  wire \DFF_65.CK ;
  wire \DFF_65.D ;
  wire \DFF_65.Q ;
  wire \DFF_650.CK ;
  wire \DFF_650.D ;
  wire \DFF_650.Q ;
  wire \DFF_651.CK ;
  wire \DFF_651.D ;
  wire \DFF_651.Q ;
  wire \DFF_652.CK ;
  wire \DFF_652.D ;
  wire \DFF_652.Q ;
  wire \DFF_653.CK ;
  wire \DFF_653.D ;
  wire \DFF_653.Q ;
  wire \DFF_654.CK ;
  wire \DFF_654.D ;
  wire \DFF_654.Q ;
  wire \DFF_655.CK ;
  wire \DFF_655.D ;
  wire \DFF_655.Q ;
  wire \DFF_656.CK ;
  wire \DFF_656.D ;
  wire \DFF_656.Q ;
  wire \DFF_657.CK ;
  wire \DFF_657.D ;
  wire \DFF_657.Q ;
  wire \DFF_658.CK ;
  wire \DFF_658.D ;
  wire \DFF_658.Q ;
  wire \DFF_659.CK ;
  wire \DFF_659.D ;
  wire \DFF_659.Q ;
  wire \DFF_66.CK ;
  wire \DFF_66.D ;
  wire \DFF_66.Q ;
  wire \DFF_660.CK ;
  wire \DFF_660.D ;
  wire \DFF_660.Q ;
  wire \DFF_661.CK ;
  wire \DFF_661.D ;
  wire \DFF_661.Q ;
  wire \DFF_662.CK ;
  wire \DFF_662.D ;
  wire \DFF_662.Q ;
  wire \DFF_663.CK ;
  wire \DFF_663.D ;
  wire \DFF_663.Q ;
  wire \DFF_664.CK ;
  wire \DFF_664.D ;
  wire \DFF_664.Q ;
  wire \DFF_665.CK ;
  wire \DFF_665.D ;
  wire \DFF_665.Q ;
  wire \DFF_666.CK ;
  wire \DFF_666.D ;
  wire \DFF_666.Q ;
  wire \DFF_667.CK ;
  wire \DFF_667.D ;
  wire \DFF_667.Q ;
  wire \DFF_668.CK ;
  wire \DFF_669.CK ;
  wire \DFF_67.CK ;
  wire \DFF_67.D ;
  wire \DFF_67.Q ;
  wire \DFF_670.CK ;
  wire \DFF_671.CK ;
  wire \DFF_672.CK ;
  wire \DFF_673.CK ;
  wire \DFF_674.CK ;
  wire \DFF_675.CK ;
  wire \DFF_676.CK ;
  wire \DFF_677.CK ;
  wire \DFF_678.CK ;
  wire \DFF_678.D ;
  wire \DFF_678.Q ;
  wire \DFF_679.CK ;
  wire \DFF_679.D ;
  wire \DFF_679.Q ;
  wire \DFF_68.CK ;
  wire \DFF_68.D ;
  wire \DFF_68.Q ;
  wire \DFF_680.CK ;
  wire \DFF_680.D ;
  wire \DFF_680.Q ;
  wire \DFF_681.CK ;
  wire \DFF_681.D ;
  wire \DFF_681.Q ;
  wire \DFF_682.CK ;
  wire \DFF_682.D ;
  wire \DFF_682.Q ;
  wire \DFF_683.CK ;
  wire \DFF_683.D ;
  wire \DFF_683.Q ;
  wire \DFF_684.CK ;
  wire \DFF_684.D ;
  wire \DFF_684.Q ;
  wire \DFF_685.CK ;
  wire \DFF_685.D ;
  wire \DFF_685.Q ;
  wire \DFF_686.CK ;
  wire \DFF_686.D ;
  wire \DFF_686.Q ;
  wire \DFF_687.CK ;
  wire \DFF_687.D ;
  wire \DFF_687.Q ;
  wire \DFF_688.CK ;
  wire \DFF_688.D ;
  wire \DFF_688.Q ;
  wire \DFF_689.CK ;
  wire \DFF_689.D ;
  wire \DFF_689.Q ;
  wire \DFF_69.CK ;
  wire \DFF_69.D ;
  wire \DFF_69.Q ;
  wire \DFF_690.CK ;
  wire \DFF_690.D ;
  wire \DFF_690.Q ;
  wire \DFF_691.CK ;
  wire \DFF_691.D ;
  wire \DFF_691.Q ;
  wire \DFF_692.CK ;
  wire \DFF_692.D ;
  wire \DFF_692.Q ;
  wire \DFF_693.CK ;
  wire \DFF_693.D ;
  wire \DFF_693.Q ;
  wire \DFF_694.CK ;
  wire \DFF_694.D ;
  wire \DFF_694.Q ;
  wire \DFF_695.CK ;
  wire \DFF_695.D ;
  wire \DFF_695.Q ;
  wire \DFF_696.CK ;
  wire \DFF_696.D ;
  wire \DFF_696.Q ;
  wire \DFF_697.CK ;
  wire \DFF_697.D ;
  wire \DFF_697.Q ;
  wire \DFF_698.CK ;
  wire \DFF_698.D ;
  wire \DFF_698.Q ;
  wire \DFF_699.CK ;
  wire \DFF_699.D ;
  wire \DFF_699.Q ;
  wire \DFF_7.CK ;
  wire \DFF_7.D ;
  wire \DFF_7.Q ;
  wire \DFF_70.CK ;
  wire \DFF_70.D ;
  wire \DFF_70.Q ;
  wire \DFF_700.CK ;
  wire \DFF_700.D ;
  wire \DFF_700.Q ;
  wire \DFF_701.CK ;
  wire \DFF_701.D ;
  wire \DFF_701.Q ;
  wire \DFF_702.CK ;
  wire \DFF_702.D ;
  wire \DFF_702.Q ;
  wire \DFF_703.CK ;
  wire \DFF_703.D ;
  wire \DFF_703.Q ;
  wire \DFF_704.CK ;
  wire \DFF_704.D ;
  wire \DFF_704.Q ;
  wire \DFF_705.CK ;
  wire \DFF_705.D ;
  wire \DFF_705.Q ;
  wire \DFF_706.CK ;
  wire \DFF_706.D ;
  wire \DFF_706.Q ;
  wire \DFF_707.CK ;
  wire \DFF_707.D ;
  wire \DFF_707.Q ;
  wire \DFF_708.CK ;
  wire \DFF_708.D ;
  wire \DFF_708.Q ;
  wire \DFF_709.CK ;
  wire \DFF_709.D ;
  wire \DFF_709.Q ;
  wire \DFF_71.CK ;
  wire \DFF_71.D ;
  wire \DFF_71.Q ;
  wire \DFF_710.CK ;
  wire \DFF_710.D ;
  wire \DFF_710.Q ;
  wire \DFF_711.CK ;
  wire \DFF_711.D ;
  wire \DFF_711.Q ;
  wire \DFF_712.CK ;
  wire \DFF_712.D ;
  wire \DFF_712.Q ;
  wire \DFF_713.CK ;
  wire \DFF_713.D ;
  wire \DFF_713.Q ;
  wire \DFF_714.CK ;
  wire \DFF_714.D ;
  wire \DFF_714.Q ;
  wire \DFF_715.CK ;
  wire \DFF_715.D ;
  wire \DFF_715.Q ;
  wire \DFF_716.CK ;
  wire \DFF_716.D ;
  wire \DFF_716.Q ;
  wire \DFF_717.CK ;
  wire \DFF_717.D ;
  wire \DFF_717.Q ;
  wire \DFF_718.CK ;
  wire \DFF_718.D ;
  wire \DFF_718.Q ;
  wire \DFF_719.CK ;
  wire \DFF_719.D ;
  wire \DFF_719.Q ;
  wire \DFF_72.CK ;
  wire \DFF_72.D ;
  wire \DFF_72.Q ;
  wire \DFF_720.CK ;
  wire \DFF_720.D ;
  wire \DFF_720.Q ;
  wire \DFF_721.CK ;
  wire \DFF_721.D ;
  wire \DFF_721.Q ;
  wire \DFF_722.CK ;
  wire \DFF_722.D ;
  wire \DFF_722.Q ;
  wire \DFF_723.CK ;
  wire \DFF_723.D ;
  wire \DFF_723.Q ;
  wire \DFF_724.CK ;
  wire \DFF_724.D ;
  wire \DFF_724.Q ;
  wire \DFF_725.CK ;
  wire \DFF_725.D ;
  wire \DFF_725.Q ;
  wire \DFF_726.CK ;
  wire \DFF_726.D ;
  wire \DFF_726.Q ;
  wire \DFF_727.CK ;
  wire \DFF_727.D ;
  wire \DFF_727.Q ;
  wire \DFF_728.CK ;
  wire \DFF_728.D ;
  wire \DFF_728.Q ;
  wire \DFF_729.CK ;
  wire \DFF_729.D ;
  wire \DFF_729.Q ;
  wire \DFF_73.CK ;
  wire \DFF_73.D ;
  wire \DFF_73.Q ;
  wire \DFF_730.CK ;
  wire \DFF_730.D ;
  wire \DFF_730.Q ;
  wire \DFF_731.CK ;
  wire \DFF_731.D ;
  wire \DFF_731.Q ;
  wire \DFF_732.CK ;
  wire \DFF_732.D ;
  wire \DFF_732.Q ;
  wire \DFF_733.CK ;
  wire \DFF_733.D ;
  wire \DFF_733.Q ;
  wire \DFF_734.CK ;
  wire \DFF_734.D ;
  wire \DFF_734.Q ;
  wire \DFF_735.CK ;
  wire \DFF_735.D ;
  wire \DFF_735.Q ;
  wire \DFF_736.CK ;
  wire \DFF_736.D ;
  wire \DFF_736.Q ;
  wire \DFF_737.CK ;
  wire \DFF_737.D ;
  wire \DFF_737.Q ;
  wire \DFF_738.CK ;
  wire \DFF_738.D ;
  wire \DFF_738.Q ;
  wire \DFF_739.CK ;
  wire \DFF_739.D ;
  wire \DFF_739.Q ;
  wire \DFF_74.CK ;
  wire \DFF_74.D ;
  wire \DFF_74.Q ;
  wire \DFF_740.CK ;
  wire \DFF_740.D ;
  wire \DFF_740.Q ;
  wire \DFF_741.CK ;
  wire \DFF_741.D ;
  wire \DFF_741.Q ;
  wire \DFF_742.CK ;
  wire \DFF_742.D ;
  wire \DFF_742.Q ;
  wire \DFF_743.CK ;
  wire \DFF_743.D ;
  wire \DFF_743.Q ;
  wire \DFF_744.CK ;
  wire \DFF_744.D ;
  wire \DFF_744.Q ;
  wire \DFF_745.CK ;
  wire \DFF_745.D ;
  wire \DFF_745.Q ;
  wire \DFF_746.CK ;
  wire \DFF_746.D ;
  wire \DFF_746.Q ;
  wire \DFF_747.CK ;
  wire \DFF_747.D ;
  wire \DFF_747.Q ;
  wire \DFF_748.CK ;
  wire \DFF_748.D ;
  wire \DFF_748.Q ;
  wire \DFF_749.CK ;
  wire \DFF_749.D ;
  wire \DFF_749.Q ;
  wire \DFF_75.CK ;
  wire \DFF_75.D ;
  wire \DFF_75.Q ;
  wire \DFF_750.CK ;
  wire \DFF_750.D ;
  wire \DFF_750.Q ;
  wire \DFF_751.CK ;
  wire \DFF_751.D ;
  wire \DFF_751.Q ;
  wire \DFF_752.CK ;
  wire \DFF_752.D ;
  wire \DFF_752.Q ;
  wire \DFF_753.CK ;
  wire \DFF_753.D ;
  wire \DFF_753.Q ;
  wire \DFF_754.CK ;
  wire \DFF_754.D ;
  wire \DFF_754.Q ;
  wire \DFF_755.CK ;
  wire \DFF_755.D ;
  wire \DFF_755.Q ;
  wire \DFF_756.CK ;
  wire \DFF_756.D ;
  wire \DFF_756.Q ;
  wire \DFF_757.CK ;
  wire \DFF_757.D ;
  wire \DFF_757.Q ;
  wire \DFF_758.CK ;
  wire \DFF_758.D ;
  wire \DFF_758.Q ;
  wire \DFF_759.CK ;
  wire \DFF_759.D ;
  wire \DFF_759.Q ;
  wire \DFF_76.CK ;
  wire \DFF_76.D ;
  wire \DFF_76.Q ;
  wire \DFF_760.CK ;
  wire \DFF_760.D ;
  wire \DFF_760.Q ;
  wire \DFF_761.CK ;
  wire \DFF_761.D ;
  wire \DFF_761.Q ;
  wire \DFF_762.CK ;
  wire \DFF_762.D ;
  wire \DFF_762.Q ;
  wire \DFF_763.CK ;
  wire \DFF_763.D ;
  wire \DFF_763.Q ;
  wire \DFF_764.CK ;
  wire \DFF_764.D ;
  wire \DFF_764.Q ;
  wire \DFF_765.CK ;
  wire \DFF_765.D ;
  wire \DFF_765.Q ;
  wire \DFF_766.CK ;
  wire \DFF_766.D ;
  wire \DFF_766.Q ;
  wire \DFF_767.CK ;
  wire \DFF_767.D ;
  wire \DFF_767.Q ;
  wire \DFF_768.CK ;
  wire \DFF_768.D ;
  wire \DFF_768.Q ;
  wire \DFF_769.CK ;
  wire \DFF_769.D ;
  wire \DFF_769.Q ;
  wire \DFF_77.CK ;
  wire \DFF_77.D ;
  wire \DFF_77.Q ;
  wire \DFF_770.CK ;
  wire \DFF_770.D ;
  wire \DFF_770.Q ;
  wire \DFF_771.CK ;
  wire \DFF_771.D ;
  wire \DFF_771.Q ;
  wire \DFF_772.CK ;
  wire \DFF_772.D ;
  wire \DFF_772.Q ;
  wire \DFF_773.CK ;
  wire \DFF_773.D ;
  wire \DFF_773.Q ;
  wire \DFF_774.CK ;
  wire \DFF_774.D ;
  wire \DFF_774.Q ;
  wire \DFF_775.CK ;
  wire \DFF_775.D ;
  wire \DFF_775.Q ;
  wire \DFF_776.CK ;
  wire \DFF_776.D ;
  wire \DFF_776.Q ;
  wire \DFF_777.CK ;
  wire \DFF_777.D ;
  wire \DFF_777.Q ;
  wire \DFF_778.CK ;
  wire \DFF_778.D ;
  wire \DFF_778.Q ;
  wire \DFF_779.CK ;
  wire \DFF_779.D ;
  wire \DFF_779.Q ;
  wire \DFF_78.CK ;
  wire \DFF_78.D ;
  wire \DFF_78.Q ;
  wire \DFF_780.CK ;
  wire \DFF_780.D ;
  wire \DFF_780.Q ;
  wire \DFF_781.CK ;
  wire \DFF_781.D ;
  wire \DFF_781.Q ;
  wire \DFF_782.CK ;
  wire \DFF_782.D ;
  wire \DFF_782.Q ;
  wire \DFF_783.CK ;
  wire \DFF_783.D ;
  wire \DFF_783.Q ;
  wire \DFF_784.CK ;
  wire \DFF_785.CK ;
  wire \DFF_786.CK ;
  wire \DFF_787.CK ;
  wire \DFF_788.CK ;
  wire \DFF_789.CK ;
  wire \DFF_79.CK ;
  wire \DFF_79.D ;
  wire \DFF_79.Q ;
  wire \DFF_790.CK ;
  wire \DFF_791.CK ;
  wire \DFF_792.CK ;
  wire \DFF_792.D ;
  wire \DFF_792.Q ;
  wire \DFF_793.CK ;
  wire \DFF_793.D ;
  wire \DFF_793.Q ;
  wire \DFF_794.CK ;
  wire \DFF_794.D ;
  wire \DFF_794.Q ;
  wire \DFF_795.CK ;
  wire \DFF_795.D ;
  wire \DFF_795.Q ;
  wire \DFF_796.CK ;
  wire \DFF_796.D ;
  wire \DFF_796.Q ;
  wire \DFF_797.CK ;
  wire \DFF_797.D ;
  wire \DFF_797.Q ;
  wire \DFF_798.CK ;
  wire \DFF_798.D ;
  wire \DFF_798.Q ;
  wire \DFF_799.CK ;
  wire \DFF_799.D ;
  wire \DFF_799.Q ;
  wire \DFF_8.CK ;
  wire \DFF_8.D ;
  wire \DFF_8.Q ;
  wire \DFF_80.CK ;
  wire \DFF_80.D ;
  wire \DFF_80.Q ;
  wire \DFF_800.CK ;
  wire \DFF_800.D ;
  wire \DFF_800.Q ;
  wire \DFF_801.CK ;
  wire \DFF_801.D ;
  wire \DFF_801.Q ;
  wire \DFF_802.CK ;
  wire \DFF_802.D ;
  wire \DFF_802.Q ;
  wire \DFF_803.CK ;
  wire \DFF_803.D ;
  wire \DFF_803.Q ;
  wire \DFF_804.CK ;
  wire \DFF_804.D ;
  wire \DFF_804.Q ;
  wire \DFF_805.CK ;
  wire \DFF_805.D ;
  wire \DFF_805.Q ;
  wire \DFF_806.CK ;
  wire \DFF_806.D ;
  wire \DFF_806.Q ;
  wire \DFF_807.CK ;
  wire \DFF_807.D ;
  wire \DFF_807.Q ;
  wire \DFF_808.CK ;
  wire \DFF_808.D ;
  wire \DFF_808.Q ;
  wire \DFF_809.CK ;
  wire \DFF_809.D ;
  wire \DFF_809.Q ;
  wire \DFF_81.CK ;
  wire \DFF_81.D ;
  wire \DFF_81.Q ;
  wire \DFF_810.CK ;
  wire \DFF_810.D ;
  wire \DFF_810.Q ;
  wire \DFF_811.CK ;
  wire \DFF_811.D ;
  wire \DFF_811.Q ;
  wire \DFF_812.CK ;
  wire \DFF_812.D ;
  wire \DFF_812.Q ;
  wire \DFF_813.CK ;
  wire \DFF_813.D ;
  wire \DFF_813.Q ;
  wire \DFF_814.CK ;
  wire \DFF_814.D ;
  wire \DFF_814.Q ;
  wire \DFF_815.CK ;
  wire \DFF_815.D ;
  wire \DFF_815.Q ;
  wire \DFF_816.CK ;
  wire \DFF_816.D ;
  wire \DFF_816.Q ;
  wire \DFF_817.CK ;
  wire \DFF_817.D ;
  wire \DFF_817.Q ;
  wire \DFF_818.CK ;
  wire \DFF_818.D ;
  wire \DFF_818.Q ;
  wire \DFF_819.CK ;
  wire \DFF_819.D ;
  wire \DFF_819.Q ;
  wire \DFF_82.CK ;
  wire \DFF_82.D ;
  wire \DFF_82.Q ;
  wire \DFF_820.CK ;
  wire \DFF_820.D ;
  wire \DFF_820.Q ;
  wire \DFF_821.CK ;
  wire \DFF_821.D ;
  wire \DFF_821.Q ;
  wire \DFF_822.CK ;
  wire \DFF_822.D ;
  wire \DFF_822.Q ;
  wire \DFF_823.CK ;
  wire \DFF_823.D ;
  wire \DFF_823.Q ;
  wire \DFF_824.CK ;
  wire \DFF_824.D ;
  wire \DFF_824.Q ;
  wire \DFF_825.CK ;
  wire \DFF_825.D ;
  wire \DFF_825.Q ;
  wire \DFF_826.CK ;
  wire \DFF_826.D ;
  wire \DFF_826.Q ;
  wire \DFF_827.CK ;
  wire \DFF_827.D ;
  wire \DFF_827.Q ;
  wire \DFF_828.CK ;
  wire \DFF_828.D ;
  wire \DFF_828.Q ;
  wire \DFF_829.CK ;
  wire \DFF_829.D ;
  wire \DFF_829.Q ;
  wire \DFF_83.CK ;
  wire \DFF_83.D ;
  wire \DFF_83.Q ;
  wire \DFF_830.CK ;
  wire \DFF_830.D ;
  wire \DFF_830.Q ;
  wire \DFF_831.CK ;
  wire \DFF_831.D ;
  wire \DFF_831.Q ;
  wire \DFF_832.CK ;
  wire \DFF_832.D ;
  wire \DFF_832.Q ;
  wire \DFF_833.CK ;
  wire \DFF_833.D ;
  wire \DFF_833.Q ;
  wire \DFF_834.CK ;
  wire \DFF_834.D ;
  wire \DFF_834.Q ;
  wire \DFF_835.CK ;
  wire \DFF_835.D ;
  wire \DFF_835.Q ;
  wire \DFF_836.CK ;
  wire \DFF_836.D ;
  wire \DFF_836.Q ;
  wire \DFF_837.CK ;
  wire \DFF_837.D ;
  wire \DFF_837.Q ;
  wire \DFF_838.CK ;
  wire \DFF_838.D ;
  wire \DFF_838.Q ;
  wire \DFF_839.CK ;
  wire \DFF_839.D ;
  wire \DFF_839.Q ;
  wire \DFF_84.CK ;
  wire \DFF_84.D ;
  wire \DFF_84.Q ;
  wire \DFF_840.CK ;
  wire \DFF_840.D ;
  wire \DFF_840.Q ;
  wire \DFF_841.CK ;
  wire \DFF_841.D ;
  wire \DFF_841.Q ;
  wire \DFF_842.CK ;
  wire \DFF_842.D ;
  wire \DFF_842.Q ;
  wire \DFF_843.CK ;
  wire \DFF_843.D ;
  wire \DFF_843.Q ;
  wire \DFF_844.CK ;
  wire \DFF_844.D ;
  wire \DFF_844.Q ;
  wire \DFF_845.CK ;
  wire \DFF_845.D ;
  wire \DFF_845.Q ;
  wire \DFF_846.CK ;
  wire \DFF_846.D ;
  wire \DFF_846.Q ;
  wire \DFF_847.CK ;
  wire \DFF_847.D ;
  wire \DFF_847.Q ;
  wire \DFF_848.CK ;
  wire \DFF_848.D ;
  wire \DFF_848.Q ;
  wire \DFF_849.CK ;
  wire \DFF_849.D ;
  wire \DFF_849.Q ;
  wire \DFF_85.CK ;
  wire \DFF_85.D ;
  wire \DFF_85.Q ;
  wire \DFF_850.CK ;
  wire \DFF_850.D ;
  wire \DFF_850.Q ;
  wire \DFF_851.CK ;
  wire \DFF_851.D ;
  wire \DFF_851.Q ;
  wire \DFF_852.CK ;
  wire \DFF_852.D ;
  wire \DFF_852.Q ;
  wire \DFF_853.CK ;
  wire \DFF_853.D ;
  wire \DFF_853.Q ;
  wire \DFF_854.CK ;
  wire \DFF_854.D ;
  wire \DFF_854.Q ;
  wire \DFF_855.CK ;
  wire \DFF_855.D ;
  wire \DFF_855.Q ;
  wire \DFF_856.CK ;
  wire \DFF_856.D ;
  wire \DFF_856.Q ;
  wire \DFF_857.CK ;
  wire \DFF_857.D ;
  wire \DFF_857.Q ;
  wire \DFF_858.CK ;
  wire \DFF_858.D ;
  wire \DFF_858.Q ;
  wire \DFF_859.CK ;
  wire \DFF_859.D ;
  wire \DFF_859.Q ;
  wire \DFF_86.CK ;
  wire \DFF_86.D ;
  wire \DFF_86.Q ;
  wire \DFF_860.CK ;
  wire \DFF_860.D ;
  wire \DFF_860.Q ;
  wire \DFF_861.CK ;
  wire \DFF_861.D ;
  wire \DFF_861.Q ;
  wire \DFF_862.CK ;
  wire \DFF_862.D ;
  wire \DFF_862.Q ;
  wire \DFF_863.CK ;
  wire \DFF_863.D ;
  wire \DFF_863.Q ;
  wire \DFF_864.CK ;
  wire \DFF_864.D ;
  wire \DFF_864.Q ;
  wire \DFF_865.CK ;
  wire \DFF_865.D ;
  wire \DFF_865.Q ;
  wire \DFF_866.CK ;
  wire \DFF_866.D ;
  wire \DFF_866.Q ;
  wire \DFF_867.CK ;
  wire \DFF_867.D ;
  wire \DFF_867.Q ;
  wire \DFF_868.CK ;
  wire \DFF_868.D ;
  wire \DFF_868.Q ;
  wire \DFF_869.CK ;
  wire \DFF_869.D ;
  wire \DFF_869.Q ;
  wire \DFF_87.CK ;
  wire \DFF_87.D ;
  wire \DFF_87.Q ;
  wire \DFF_870.CK ;
  wire \DFF_870.D ;
  wire \DFF_870.Q ;
  wire \DFF_871.CK ;
  wire \DFF_871.D ;
  wire \DFF_871.Q ;
  wire \DFF_872.CK ;
  wire \DFF_872.D ;
  wire \DFF_872.Q ;
  wire \DFF_873.CK ;
  wire \DFF_873.D ;
  wire \DFF_873.Q ;
  wire \DFF_874.CK ;
  wire \DFF_874.D ;
  wire \DFF_874.Q ;
  wire \DFF_875.CK ;
  wire \DFF_875.D ;
  wire \DFF_875.Q ;
  wire \DFF_876.CK ;
  wire \DFF_876.D ;
  wire \DFF_876.Q ;
  wire \DFF_877.CK ;
  wire \DFF_877.D ;
  wire \DFF_877.Q ;
  wire \DFF_878.CK ;
  wire \DFF_878.D ;
  wire \DFF_878.Q ;
  wire \DFF_879.CK ;
  wire \DFF_879.D ;
  wire \DFF_879.Q ;
  wire \DFF_88.CK ;
  wire \DFF_88.D ;
  wire \DFF_88.Q ;
  wire \DFF_880.CK ;
  wire \DFF_880.D ;
  wire \DFF_880.Q ;
  wire \DFF_881.CK ;
  wire \DFF_881.D ;
  wire \DFF_881.Q ;
  wire \DFF_882.CK ;
  wire \DFF_882.D ;
  wire \DFF_882.Q ;
  wire \DFF_883.CK ;
  wire \DFF_883.D ;
  wire \DFF_883.Q ;
  wire \DFF_884.CK ;
  wire \DFF_884.D ;
  wire \DFF_884.Q ;
  wire \DFF_885.CK ;
  wire \DFF_885.D ;
  wire \DFF_885.Q ;
  wire \DFF_886.CK ;
  wire \DFF_886.D ;
  wire \DFF_886.Q ;
  wire \DFF_887.CK ;
  wire \DFF_887.D ;
  wire \DFF_887.Q ;
  wire \DFF_888.CK ;
  wire \DFF_888.D ;
  wire \DFF_888.Q ;
  wire \DFF_889.CK ;
  wire \DFF_889.D ;
  wire \DFF_889.Q ;
  wire \DFF_89.CK ;
  wire \DFF_89.D ;
  wire \DFF_89.Q ;
  wire \DFF_890.CK ;
  wire \DFF_890.D ;
  wire \DFF_890.Q ;
  wire \DFF_891.CK ;
  wire \DFF_891.D ;
  wire \DFF_891.Q ;
  wire \DFF_892.CK ;
  wire \DFF_892.D ;
  wire \DFF_892.Q ;
  wire \DFF_893.CK ;
  wire \DFF_893.D ;
  wire \DFF_893.Q ;
  wire \DFF_894.CK ;
  wire \DFF_894.D ;
  wire \DFF_894.Q ;
  wire \DFF_895.CK ;
  wire \DFF_895.D ;
  wire \DFF_895.Q ;
  wire \DFF_896.CK ;
  wire \DFF_896.D ;
  wire \DFF_896.Q ;
  wire \DFF_897.CK ;
  wire \DFF_897.D ;
  wire \DFF_897.Q ;
  wire \DFF_898.CK ;
  wire \DFF_898.D ;
  wire \DFF_898.Q ;
  wire \DFF_899.CK ;
  wire \DFF_899.D ;
  wire \DFF_899.Q ;
  wire \DFF_9.CK ;
  wire \DFF_9.D ;
  wire \DFF_9.Q ;
  wire \DFF_90.CK ;
  wire \DFF_90.D ;
  wire \DFF_90.Q ;
  wire \DFF_900.CK ;
  wire \DFF_900.D ;
  wire \DFF_900.Q ;
  wire \DFF_901.CK ;
  wire \DFF_901.D ;
  wire \DFF_901.Q ;
  wire \DFF_902.CK ;
  wire \DFF_902.D ;
  wire \DFF_902.Q ;
  wire \DFF_903.CK ;
  wire \DFF_903.D ;
  wire \DFF_903.Q ;
  wire \DFF_904.CK ;
  wire \DFF_904.D ;
  wire \DFF_904.Q ;
  wire \DFF_905.CK ;
  wire \DFF_905.D ;
  wire \DFF_905.Q ;
  wire \DFF_906.CK ;
  wire \DFF_906.D ;
  wire \DFF_906.Q ;
  wire \DFF_907.CK ;
  wire \DFF_907.D ;
  wire \DFF_907.Q ;
  wire \DFF_908.CK ;
  wire \DFF_908.D ;
  wire \DFF_908.Q ;
  wire \DFF_909.CK ;
  wire \DFF_909.D ;
  wire \DFF_909.Q ;
  wire \DFF_91.CK ;
  wire \DFF_91.D ;
  wire \DFF_91.Q ;
  wire \DFF_910.CK ;
  wire \DFF_910.D ;
  wire \DFF_910.Q ;
  wire \DFF_911.CK ;
  wire \DFF_911.D ;
  wire \DFF_911.Q ;
  wire \DFF_912.CK ;
  wire \DFF_912.D ;
  wire \DFF_912.Q ;
  wire \DFF_913.CK ;
  wire \DFF_913.D ;
  wire \DFF_913.Q ;
  wire \DFF_914.CK ;
  wire \DFF_914.D ;
  wire \DFF_914.Q ;
  wire \DFF_915.CK ;
  wire \DFF_915.D ;
  wire \DFF_915.Q ;
  wire \DFF_916.CK ;
  wire \DFF_916.D ;
  wire \DFF_916.Q ;
  wire \DFF_917.CK ;
  wire \DFF_917.D ;
  wire \DFF_917.Q ;
  wire \DFF_918.CK ;
  wire \DFF_918.D ;
  wire \DFF_918.Q ;
  wire \DFF_919.CK ;
  wire \DFF_919.D ;
  wire \DFF_919.Q ;
  wire \DFF_92.CK ;
  wire \DFF_92.D ;
  wire \DFF_92.Q ;
  wire \DFF_920.CK ;
  wire \DFF_920.D ;
  wire \DFF_920.Q ;
  wire \DFF_921.CK ;
  wire \DFF_921.D ;
  wire \DFF_921.Q ;
  wire \DFF_922.CK ;
  wire \DFF_922.D ;
  wire \DFF_922.Q ;
  wire \DFF_923.CK ;
  wire \DFF_923.D ;
  wire \DFF_923.Q ;
  wire \DFF_924.CK ;
  wire \DFF_924.D ;
  wire \DFF_924.Q ;
  wire \DFF_925.CK ;
  wire \DFF_925.D ;
  wire \DFF_925.Q ;
  wire \DFF_926.CK ;
  wire \DFF_926.D ;
  wire \DFF_926.Q ;
  wire \DFF_927.CK ;
  wire \DFF_927.D ;
  wire \DFF_927.Q ;
  wire \DFF_928.CK ;
  wire \DFF_928.D ;
  wire \DFF_928.Q ;
  wire \DFF_929.CK ;
  wire \DFF_929.D ;
  wire \DFF_929.Q ;
  wire \DFF_93.CK ;
  wire \DFF_93.D ;
  wire \DFF_93.Q ;
  wire \DFF_930.CK ;
  wire \DFF_930.D ;
  wire \DFF_930.Q ;
  wire \DFF_931.CK ;
  wire \DFF_931.D ;
  wire \DFF_931.Q ;
  wire \DFF_932.CK ;
  wire \DFF_932.D ;
  wire \DFF_932.Q ;
  wire \DFF_933.CK ;
  wire \DFF_933.D ;
  wire \DFF_933.Q ;
  wire \DFF_934.CK ;
  wire \DFF_934.D ;
  wire \DFF_934.Q ;
  wire \DFF_935.CK ;
  wire \DFF_935.D ;
  wire \DFF_935.Q ;
  wire \DFF_936.CK ;
  wire \DFF_936.D ;
  wire \DFF_936.Q ;
  wire \DFF_937.CK ;
  wire \DFF_937.D ;
  wire \DFF_937.Q ;
  wire \DFF_938.CK ;
  wire \DFF_938.D ;
  wire \DFF_938.Q ;
  wire \DFF_939.CK ;
  wire \DFF_939.D ;
  wire \DFF_939.Q ;
  wire \DFF_94.CK ;
  wire \DFF_94.D ;
  wire \DFF_94.Q ;
  wire \DFF_940.CK ;
  wire \DFF_940.D ;
  wire \DFF_940.Q ;
  wire \DFF_941.CK ;
  wire \DFF_941.D ;
  wire \DFF_941.Q ;
  wire \DFF_942.CK ;
  wire \DFF_942.D ;
  wire \DFF_942.Q ;
  wire \DFF_943.CK ;
  wire \DFF_943.D ;
  wire \DFF_943.Q ;
  wire \DFF_944.CK ;
  wire \DFF_944.D ;
  wire \DFF_944.Q ;
  wire \DFF_945.CK ;
  wire \DFF_945.D ;
  wire \DFF_945.Q ;
  wire \DFF_946.CK ;
  wire \DFF_946.D ;
  wire \DFF_946.Q ;
  wire \DFF_947.CK ;
  wire \DFF_947.D ;
  wire \DFF_947.Q ;
  wire \DFF_948.CK ;
  wire \DFF_948.D ;
  wire \DFF_948.Q ;
  wire \DFF_949.CK ;
  wire \DFF_949.D ;
  wire \DFF_949.Q ;
  wire \DFF_95.CK ;
  wire \DFF_95.D ;
  wire \DFF_95.Q ;
  wire \DFF_950.CK ;
  wire \DFF_950.D ;
  wire \DFF_950.Q ;
  wire \DFF_951.CK ;
  wire \DFF_951.D ;
  wire \DFF_951.Q ;
  wire \DFF_952.CK ;
  wire \DFF_952.D ;
  wire \DFF_952.Q ;
  wire \DFF_953.CK ;
  wire \DFF_953.D ;
  wire \DFF_953.Q ;
  wire \DFF_954.CK ;
  wire \DFF_954.D ;
  wire \DFF_954.Q ;
  wire \DFF_955.CK ;
  wire \DFF_955.D ;
  wire \DFF_955.Q ;
  wire \DFF_956.CK ;
  wire \DFF_956.D ;
  wire \DFF_956.Q ;
  wire \DFF_957.CK ;
  wire \DFF_957.D ;
  wire \DFF_957.Q ;
  wire \DFF_958.CK ;
  wire \DFF_958.D ;
  wire \DFF_958.Q ;
  wire \DFF_959.CK ;
  wire \DFF_959.D ;
  wire \DFF_959.Q ;
  wire \DFF_96.CK ;
  wire \DFF_96.D ;
  wire \DFF_96.Q ;
  wire \DFF_960.CK ;
  wire \DFF_960.D ;
  wire \DFF_960.Q ;
  wire \DFF_961.CK ;
  wire \DFF_961.D ;
  wire \DFF_961.Q ;
  wire \DFF_962.CK ;
  wire \DFF_962.D ;
  wire \DFF_962.Q ;
  wire \DFF_963.CK ;
  wire \DFF_963.D ;
  wire \DFF_963.Q ;
  wire \DFF_964.CK ;
  wire \DFF_964.D ;
  wire \DFF_964.Q ;
  wire \DFF_965.CK ;
  wire \DFF_965.D ;
  wire \DFF_965.Q ;
  wire \DFF_966.CK ;
  wire \DFF_966.D ;
  wire \DFF_966.Q ;
  wire \DFF_967.CK ;
  wire \DFF_967.D ;
  wire \DFF_967.Q ;
  wire \DFF_968.CK ;
  wire \DFF_968.D ;
  wire \DFF_968.Q ;
  wire \DFF_969.CK ;
  wire \DFF_969.D ;
  wire \DFF_969.Q ;
  wire \DFF_97.CK ;
  wire \DFF_97.D ;
  wire \DFF_97.Q ;
  wire \DFF_970.CK ;
  wire \DFF_970.D ;
  wire \DFF_970.Q ;
  wire \DFF_971.CK ;
  wire \DFF_971.D ;
  wire \DFF_971.Q ;
  wire \DFF_972.CK ;
  wire \DFF_972.D ;
  wire \DFF_972.Q ;
  wire \DFF_973.CK ;
  wire \DFF_973.D ;
  wire \DFF_973.Q ;
  wire \DFF_974.CK ;
  wire \DFF_974.D ;
  wire \DFF_974.Q ;
  wire \DFF_975.CK ;
  wire \DFF_975.D ;
  wire \DFF_975.Q ;
  wire \DFF_976.CK ;
  wire \DFF_976.D ;
  wire \DFF_976.Q ;
  wire \DFF_977.CK ;
  wire \DFF_977.D ;
  wire \DFF_977.Q ;
  wire \DFF_978.CK ;
  wire \DFF_978.D ;
  wire \DFF_978.Q ;
  wire \DFF_979.CK ;
  wire \DFF_979.D ;
  wire \DFF_979.Q ;
  wire \DFF_98.CK ;
  wire \DFF_98.D ;
  wire \DFF_98.Q ;
  wire \DFF_980.CK ;
  wire \DFF_980.D ;
  wire \DFF_980.Q ;
  wire \DFF_981.CK ;
  wire \DFF_981.D ;
  wire \DFF_981.Q ;
  wire \DFF_982.CK ;
  wire \DFF_982.D ;
  wire \DFF_982.Q ;
  wire \DFF_983.CK ;
  wire \DFF_983.D ;
  wire \DFF_983.Q ;
  wire \DFF_984.CK ;
  wire \DFF_984.D ;
  wire \DFF_984.Q ;
  wire \DFF_985.CK ;
  wire \DFF_985.D ;
  wire \DFF_985.Q ;
  wire \DFF_986.CK ;
  wire \DFF_986.D ;
  wire \DFF_986.Q ;
  wire \DFF_987.CK ;
  wire \DFF_987.D ;
  wire \DFF_987.Q ;
  wire \DFF_988.CK ;
  wire \DFF_988.D ;
  wire \DFF_988.Q ;
  wire \DFF_989.CK ;
  wire \DFF_989.D ;
  wire \DFF_989.Q ;
  wire \DFF_99.CK ;
  wire \DFF_99.D ;
  wire \DFF_99.Q ;
  wire \DFF_990.CK ;
  wire \DFF_990.D ;
  wire \DFF_990.Q ;
  wire \DFF_991.CK ;
  wire \DFF_991.D ;
  wire \DFF_991.Q ;
  wire \DFF_992.CK ;
  wire \DFF_992.D ;
  wire \DFF_992.Q ;
  wire \DFF_993.CK ;
  wire \DFF_993.D ;
  wire \DFF_993.Q ;
  wire \DFF_994.CK ;
  wire \DFF_994.D ;
  wire \DFF_994.Q ;
  wire \DFF_995.CK ;
  wire \DFF_995.D ;
  wire \DFF_995.Q ;
  wire \DFF_996.CK ;
  wire \DFF_996.D ;
  wire \DFF_996.Q ;
  wire \DFF_997.CK ;
  wire \DFF_997.D ;
  wire \DFF_997.Q ;
  wire \DFF_998.CK ;
  wire \DFF_998.D ;
  wire \DFF_998.Q ;
  wire \DFF_999.CK ;
  wire \DFF_999.D ;
  wire \DFF_999.Q ;
  input GND;
  wire II13430;
  wire II13433;
  wire II13501;
  wire II13504;
  wire II13575;
  wire II13578;
  wire II13601;
  wire II13604;
  wire II13652;
  wire II13655;
  wire II13677;
  wire II13680;
  wire II13742;
  wire II13745;
  wire II13775;
  wire II13801;
  wire II13804;
  wire II13820;
  wire II13849;
  wire II13868;
  wire II14163;
  wire II14219;
  wire II14280;
  wire II14306;
  wire II14338;
  wire II14357;
  wire II14402;
  wire II14424;
  wire II14442;
  wire II14459;
  wire II14489;
  wire II14513;
  wire II15562;
  wire II15580;
  wire II15629;
  wire II15850;
  wire II15873;
  wire II15887;
  wire II15899;
  wire II15909;
  wire II15922;
  wire II15932;
  wire II15946;
  wire II15964;
  wire II15975;
  wire II15995;
  wire II16024;
  wire II16056;
  wire II17632;
  wire II17637;
  wire II17641;
  wire II17645;
  wire II17649;
  wire II17653;
  wire II17658;
  wire II17662;
  wire II17666;
  wire II17670;
  wire II17677;
  wire II17681;
  wire II17685;
  wire II17689;
  wire II17698;
  wire II17701;
  wire II17705;
  wire II17709;
  wire II17721;
  wire II17724;
  wire II17727;
  wire II17730;
  wire II17734;
  wire II17750;
  wire II17753;
  wire II17756;
  wire II17759;
  wire II17762;
  wire II17780;
  wire II17783;
  wire II17786;
  wire II17789;
  wire II17792;
  wire II17813;
  wire II17816;
  wire II17822;
  wire II17825;
  wire II17828;
  wire II17831;
  wire II17849;
  wire II17860;
  wire II17863;
  wire II17869;
  wire II17872;
  wire II17907;
  wire II17910;
  wire II17916;
  wire II17942;
  wire II17945;
  wire II17969;
  wire II17972;
  wire II17998;
  wire II18013;
  wire II18016;
  wire II18055;
  wire II18070;
  wire II18085;
  wire II18088;
  wire II18130;
  wire II18136;
  wire II18151;
  wire II18166;
  wire II18181;
  wire II18184;
  wire II18226;
  wire II18238;
  wire II18244;
  wire II18259;
  wire II18274;
  wire II18311;
  wire II18329;
  wire II18341;
  wire II18347;
  wire II18362;
  wire II18405;
  wire II18423;
  wire II18435;
  wire II18441;
  wire II18449;
  wire II18452;
  wire II18455;
  wire II18458;
  wire II18461;
  wire II18503;
  wire II18506;
  wire II18509;
  wire II18530;
  wire II18533;
  wire II18536;
  wire II18539;
  wire II18542;
  wire II18584;
  wire II18587;
  wire II18590;
  wire II18611;
  wire II18614;
  wire II18617;
  wire II18620;
  wire II18623;
  wire II18665;
  wire II18668;
  wire II18671;
  wire II18692;
  wire II18695;
  wire II18698;
  wire II18701;
  wire II18704;
  wire II18746;
  wire II18749;
  wire II18752;
  wire II18773;
  wire II18780;
  wire II18787;
  wire II18794;
  wire II18810;
  wire II18813;
  wire II18820;
  wire II18827;
  wire II18835;
  wire II18838;
  wire II18845;
  wire II18854;
  wire II18857;
  wire II18866;
  wire II18969;
  wire II19030;
  wire II19105;
  wire II19195;
  wire II19307;
  wire II19718;
  wire II19727;
  wire II19733;
  wire II19747;
  wire II19750;
  wire II19767;
  wire II19784;
  wire II19787;
  wire II19808;
  wire II19833;
  wire II19836;
  wire II19869;
  wire II19905;
  wire II20299;
  wire II20320;
  wire II20328;
  wire II20347;
  wire II20351;
  wire II20359;
  wire II20382;
  wire II20386;
  wire II20390;
  wire II20398;
  wire II20410;
  wire II20417;
  wire II20421;
  wire II20425;
  wire II20444;
  wire II20451;
  wire II20458;
  wire II20462;
  wire II20479;
  wire II20486;
  wire II20493;
  wire II20500;
  wire II20529;
  wire II20532;
  wire II20535;
  wire II20538;
  wire II20541;
  wire II20544;
  wire II20547;
  wire II20550;
  wire II20553;
  wire II20577;
  wire II20580;
  wire II20583;
  wire II20586;
  wire II20589;
  wire II20592;
  wire II20595;
  wire II20598;
  wire II20601;
  wire II20625;
  wire II20628;
  wire II20631;
  wire II20634;
  wire II20637;
  wire II20640;
  wire II20643;
  wire II20646;
  wire II20649;
  wire II20673;
  wire II20676;
  wire II20679;
  wire II20682;
  wire II20685;
  wire II20688;
  wire II20691;
  wire II20694;
  wire II20697;
  wire II21381;
  wire II21420;
  wire II24913;
  wire II25258;
  wire II25308;
  wire II25315;
  wire II25320;
  wire II25325;
  wire II26960;
  wire II26972;
  wire II26985;
  wire II32248;
  wire II32251;
  wire II33257;
  wire II33260;
  wire II34029;
  wire II34032;
  wire II35373;
  wire II35708;
  wire II35711;
  wire II35723;
  wire II36046;
  wire II36162;
  wire II36224;
  wire II36234;
  wire II36362;
  wire II36864;
  wire II37182;
  wire II37188;
  wire II37200;
  wire II37232;
  wire II37252;
  wire II37266;
  wire II37319;
  wire II37400;
  wire II37629;
  wire II37635;
  wire II37647;
  wire II37653;
  wire II37662;
  wire II37793;
  wire II38128;
  wire II38241;
  wire II38330;
  wire II38339;
  wire II38462;
  wire II38764;
  wire II38767;
  wire II38770;
  wire II38801;
  wire II38807;
  wire II39086;
  wire II39089;
  input VDD;
  wire g1;
  wire g1000;
  wire g10004;
  wire g1001;
  wire g10015;
  wire g10016;
  wire g10017;
  wire g10018;
  wire g1002;
  wire g10021;
  wire g1003;
  wire g1004;
  wire g10049;
  wire g1005;
  wire g10052;
  wire g1006;
  wire g10067;
  wire g1007;
  wire g10070;
  wire g1008;
  wire g10086;
  wire g10087;
  wire g1009;
  wire g10090;
  wire g10096;
  wire g10099;
  wire g101;
  wire g1010;
  wire g10109;
  wire g1011;
  wire g1012;
  wire g10124;
  wire g10125;
  wire g10126;
  wire g10127;
  wire g10130;
  wire g10158;
  wire g10161;
  wire g10176;
  wire g10179;
  wire g1018;
  wire g10189;
  wire g10214;
  wire g10229;
  wire g10230;
  wire g10231;
  wire g10232;
  wire g10235;
  wire g1024;
  wire g10263;
  wire g10266;
  wire g10273;
  wire g10276;
  wire g1029;
  wire g1030;
  wire g10316;
  wire g1033;
  wire g10331;
  wire g10332;
  wire g10333;
  wire g10334;
  wire g10337;
  wire g10357;
  wire g1036;
  wire g1037;
  wire g1038;
  wire g1039;
  wire g1040;
  wire g10409;
  wire g1041;
  wire g10416;
  wire g10419;
  wire g10424;
  wire g1044;
  wire g1045;
  wire g1048;
  wire g10481;
  wire g10482;
  wire g10486;
  wire g105;
  wire g10500;
  wire g1051;
  wire g1052;
  wire g1053;
  wire g1054;
  wire g10542;
  wire g10545;
  wire g10549;
  wire g1055;
  wire g1056;
  wire g10560;
  wire g10574;
  wire g1059;
  wire g1060;
  wire g10601;
  wire g10606;
  wire g10617;
  wire g1063;
  wire g10631;
  wire g10646;
  wire g10653;
  wire g1066;
  wire g10664;
  wire g1067;
  wire g1068;
  wire g10683;
  wire g1069;
  wire g10694;
  wire g1070;
  wire g1071;
  wire g10714;
  wire g10730;
  wire g10735;
  wire g1074;
  wire g10749;
  wire g1075;
  wire g10754;
  wire g10766;
  wire g10767;
  wire g10772;
  wire g10773;
  wire g1078;
  wire g10783;
  wire g10787;
  wire g10788;
  wire g10792;
  wire g10796;
  wire g10800;
  wire g10804;
  wire g10808;
  wire g1081;
  wire g10813;
  wire g10817;
  wire g1082;
  wire g10821;
  wire g10825;
  wire g10826;
  wire g1083;
  wire g10830;
  wire g10834;
  wire g10838;
  wire g1084;
  wire g10842;
  wire g10843;
  wire g10849;
  wire g1085;
  wire g10850;
  wire g10854;
  wire g10858;
  wire g10859;
  wire g10862;
  wire g10868;
  wire g10869;
  wire g10870;
  wire g10871;
  wire g10875;
  wire g10876;
  wire g10877;
  wire g1088;
  wire g10880;
  wire g10883;
  wire g10887;
  wire g10888;
  wire g10889;
  wire g1089;
  wire g10890;
  wire g10891;
  wire g10892;
  wire g10895;
  wire g10898;
  wire g109;
  wire g1090;
  wire g10901;
  wire g10907;
  wire g10908;
  wire g10909;
  wire g1091;
  wire g10910;
  wire g10911;
  wire g10912;
  wire g10915;
  wire g10918;
  wire g1092;
  wire g10921;
  wire g10924;
  wire g10930;
  wire g10931;
  wire g10932;
  wire g10933;
  wire g10934;
  wire g10935;
  wire g10936;
  wire g10937;
  wire g10940;
  wire g10943;
  wire g10946;
  wire g10949;
  wire g1095;
  wire g10963;
  wire g10966;
  wire g10967;
  wire g10968;
  wire g10969;
  wire g10972;
  wire g10973;
  wire g10974;
  wire g10977;
  wire g1098;
  wire g10980;
  wire g10983;
  wire g10988;
  wire g10991;
  wire g10994;
  wire g10995;
  wire g10996;
  wire g10999;
  wire g11;
  wire g11002;
  wire g11003;
  wire g11004;
  wire g11007;
  wire g11008;
  wire g1101;
  wire g11011;
  wire g11014;
  wire g11017;
  wire g11022;
  wire g11025;
  wire g11028;
  wire g11031;
  wire g11035;
  wire g11036;
  wire g11039;
  wire g1104;
  wire g11042;
  wire g11045;
  wire g11048;
  wire g11051;
  wire g11054;
  wire g11055;
  wire g11056;
  wire g11063;
  wire g11066;
  wire g11069;
  wire g1107;
  wire g11079;
  wire g11082;
  wire g11085;
  wire g11091;
  wire g11092;
  wire g11095;
  wire g11098;
  wire g1110;
  wire g11101;
  wire g11105;
  wire g11108;
  wire g11111;
  wire g11114;
  wire g11117;
  wire g11120;
  wire g11123;
  wire g11126;
  wire g11129;
  wire g1113;
  wire g11132;
  wire g11135;
  wire g11138;
  wire g1114;
  wire g11144;
  wire g11145;
  wire g11148;
  wire g1115;
  wire g11151;
  wire g11157;
  wire g1116;
  wire g11160;
  wire g11163;
  wire g11166;
  wire g11169;
  wire g11173;
  wire g11176;
  wire g11179;
  wire g11182;
  wire g11185;
  wire g1119;
  wire g11190;
  wire g11199;
  wire g11202;
  wire g11205;
  wire g11208;
  wire g11209;
  wire g11213;
  wire g11216;
  wire g11219;
  wire g1122;
  wire g11222;
  wire g11228;
  wire g11231;
  wire g11234;
  wire g11237;
  wire g11243;
  wire g11246;
  wire g11249;
  wire g1125;
  wire g11252;
  wire g11255;
  wire g11259;
  wire g11265;
  wire g11268;
  wire g11271;
  wire g11274;
  wire g11277;
  wire g1128;
  wire g11281;
  wire g11284;
  wire g11287;
  wire g11290;
  wire g11291;
  wire g11297;
  wire g113;
  wire g11300;
  wire g11303;
  wire g11306;
  wire g1131;
  wire g11312;
  wire g11315;
  wire g11318;
  wire g11321;
  wire g11327;
  wire g11332;
  wire g1134;
  wire g11341;
  wire g11344;
  wire g11348;
  wire g1135;
  wire g11351;
  wire g11354;
  wire g11358;
  wire g1136;
  wire g11361;
  wire g11364;
  wire g11367;
  wire g1137;
  wire g11370;
  wire g11376;
  wire g11379;
  wire g1138;
  wire g11382;
  wire g11385;
  wire g11386;
  wire g1139;
  wire g11392;
  wire g11395;
  wire g11398;
  wire g1140;
  wire g11401;
  wire g11407;
  wire g1141;
  wire g11411;
  wire g11414;
  wire g11417;
  wire g1142;
  wire g11422;
  wire g11425;
  wire g11428;
  wire g11432;
  wire g11435;
  wire g11438;
  wire g11444;
  wire g11447;
  wire g1145;
  wire g11450;
  wire g11453;
  wire g11456;
  wire g11462;
  wire g11465;
  wire g11468;
  wire g11471;
  wire g11472;
  wire g11478;
  wire g1148;
  wire g11481;
  wire g11490;
  wire g11491;
  wire g11492;
  wire g11493;
  wire g11494;
  wire g11495;
  wire g11496;
  wire g11497;
  wire g11498;
  wire g11499;
  wire g11500;
  wire g11501;
  wire g11502;
  wire g11503;
  wire g11504;
  wire g11505;
  wire g11506;
  wire g11507;
  wire g11508;
  wire g11509;
  wire g1151;
  wire g11510;
  wire g11511;
  wire g11512;
  wire g11513;
  wire g11514;
  wire g11515;
  wire g11516;
  wire g11517;
  wire g11518;
  wire g11519;
  wire g1152;
  wire g11520;
  wire g11521;
  wire g11522;
  wire g11523;
  wire g11524;
  wire g11525;
  wire g11526;
  wire g11527;
  wire g11528;
  wire g11529;
  wire g11530;
  wire g11531;
  wire g11532;
  wire g11533;
  wire g11534;
  wire g11535;
  wire g11536;
  wire g11537;
  wire g11538;
  wire g11539;
  wire g11540;
  wire g11541;
  wire g11542;
  wire g11543;
  wire g11544;
  wire g11545;
  wire g11546;
  wire g11547;
  wire g11548;
  wire g11549;
  wire g1155;
  wire g11550;
  wire g11551;
  wire g11552;
  wire g11553;
  wire g11554;
  wire g11555;
  wire g11556;
  wire g11557;
  wire g11558;
  wire g11559;
  wire g11560;
  wire g11561;
  wire g11562;
  wire g11563;
  wire g11564;
  wire g11565;
  wire g11566;
  wire g11567;
  wire g11568;
  wire g11569;
  wire g11570;
  wire g11571;
  wire g11572;
  wire g11573;
  wire g11574;
  wire g11575;
  wire g11576;
  wire g11577;
  wire g11578;
  wire g11579;
  wire g1158;
  wire g11580;
  wire g11581;
  wire g11582;
  wire g11583;
  wire g11584;
  wire g11585;
  wire g11586;
  wire g11587;
  wire g11588;
  wire g11589;
  wire g11590;
  wire g11591;
  wire g11592;
  wire g11593;
  wire g11594;
  wire g11595;
  wire g11596;
  wire g11597;
  wire g11598;
  wire g11599;
  wire g11603;
  wire g11606;
  wire g11608;
  wire g1161;
  wire g11611;
  wire g11613;
  wire g11616;
  wire g11623;
  wire g11628;
  wire g11629;
  wire g11633;
  wire g11636;
  wire g11638;
  wire g1164;
  wire g11641;
  wire g1165;
  wire g11651;
  wire g11652;
  wire g11656;
  wire g11659;
  wire g1166;
  wire g1167;
  wire g11670;
  wire g11671;
  wire g1168;
  wire g11682;
  wire g117;
  wire g11706;
  wire g1171;
  wire g11713;
  wire g1172;
  wire g1173;
  wire g11737;
  wire g1174;
  wire g11743;
  wire g1175;
  wire g11758;
  wire g1176;
  wire g11766;
  wire g11769;
  wire g1177;
  wire g11779;
  wire g11786;
  wire g11798;
  wire g1180;
  wire g11812;
  wire g11821;
  wire g11827;
  wire g1183;
  wire g11845;
  wire g11854;
  wire g11859;
  wire g1186;
  wire g11869;
  wire g11888;
  wire g11894;
  wire g11901;
  wire g11911;
  wire g1192;
  wire g11927;
  wire g1193;
  wire g11933;
  wire g11937;
  wire g11944;
  wire g11951;
  wire g1196;
  wire g11961;
  wire g11973;
  wire g11976;
  wire g11986;
  wire g1199;
  wire g11990;
  wire g11997;
  wire g12004;
  wire g12025;
  wire g12027;
  wire g12030;
  wire g12042;
  wire g12045;
  wire g12055;
  wire g12059;
  wire g1206;
  wire g12066;
  wire g12089;
  wire g1209;
  wire g12091;
  wire g12094;
  wire g121;
  wire g1210;
  wire g12106;
  wire g12109;
  wire g1211;
  wire g12119;
  wire g12123;
  wire g12136;
  wire g12139;
  wire g1214;
  wire g12142;
  wire g1215;
  wire g1216;
  wire g12161;
  wire g12163;
  wire g12166;
  wire g1217;
  wire g12178;
  wire g1218;
  wire g12181;
  wire g1219;
  wire g12198;
  wire g1220;
  wire g12201;
  wire g12204;
  wire g1221;
  wire g1222;
  wire g12223;
  wire g12225;
  wire g12228;
  wire g1223;
  wire g12239;
  wire g1224;
  wire g12242;
  wire g12253;
  wire g12256;
  wire g12259;
  wire g1227;
  wire g12279;
  wire g1228;
  wire g12282;
  wire g12285;
  wire g1229;
  wire g12296;
  wire g12299;
  wire g1230;
  wire g12302;
  wire g1231;
  wire g12312;
  wire g12315;
  wire g12318;
  wire g12321;
  wire g12332;
  wire g12333;
  wire g12336;
  wire g1234;
  wire g12340;
  wire g12343;
  wire g12346;
  wire g12349;
  wire g1235;
  wire g1236;
  wire g12362;
  wire g12363;
  wire g12366;
  wire g1237;
  wire g12370;
  wire g12373;
  wire g12378;
  wire g12379;
  wire g12382;
  wire g12385;
  wire g12389;
  wire g1240;
  wire g12408;
  wire g12409;
  wire g12412;
  wire g12415;
  wire g12420;
  wire g12421;
  wire g12424;
  wire g12425;
  wire g12426;
  wire g1243;
  wire g12430;
  wire g12432;
  wire g12433;
  wire g12434;
  wire g12435;
  wire g12437;
  wire g12438;
  wire g1244;
  wire g12440;
  wire g12442;
  wire g12445;
  wire g1245;
  wire g12450;
  wire g12457;
  wire g12467;
  wire g1248;
  wire g12482;
  wire g12487;
  input g1249;
  wire g12499;
  wire g125;
  wire g1250;
  wire g12507;
  wire g1251;
  wire g12519;
  wire g1252;
  wire g12524;
  wire g1253;
  wire g12534;
  wire g12539;
  wire g1254;
  wire g12543;
  wire g1255;
  wire g12552;
  wire g1256;
  wire g12564;
  wire g12565;
  wire g1257;
  wire g1258;
  wire g1259;
  wire g1260;
  wire g12607;
  wire g12608;
  wire g1261;
  wire g12611;
  wire g1262;
  wire g1263;
  wire g1264;
  wire g1265;
  wire g12654;
  wire g12657;
  wire g1266;
  wire g1267;
  wire g1268;
  wire g1269;
  wire g12699;
  wire g1270;
  wire g12708;
  wire g1271;
  wire g12711;
  wire g1272;
  wire g1273;
  wire g12756;
  wire g1276;
  wire g12765;
  wire g1279;
  wire g12798;
  wire g12811;
  wire g1282;
  wire g12837;
  wire g1285;
  wire g1288;
  wire g129;
  wire g12909;
  wire g1291;
  wire g1294;
  wire g12962;
  wire g1297;
  wire g130;
  wire g1300;
  wire g1303;
  wire g1306;
  wire g13070;
  wire g1309;
  wire g131;
  wire g13110;
  wire g13111;
  wire g1312;
  wire g13124;
  wire g13135;
  wire g13143;
  wire g13149;
  wire g1315;
  wire g13155;
  wire g1316;
  wire g13160;
  wire g13164;
  wire g13171;
  wire g13175;
  wire g13182;
  wire g1319;
  wire g13194;
  wire g132;
  wire g13215;
  wire g13229;
  wire g13234;
  wire g13246;
  wire g13248;
  wire g13252;
  wire g13257;
  wire g1326;
  wire g13265;
  wire g13267;
  wire g13269;
  wire g13271;
  wire g13275;
  wire g13280;
  wire g13290;
  wire g13292;
  wire g13294;
  wire g13296;
  wire g133;
  wire g13300;
  wire g13317;
  wire g13318;
  wire g13319;
  wire g1332;
  wire g13321;
  wire g13323;
  wire g13325;
  wire g13327;
  wire g13336;
  wire g13339;
  wire g13341;
  wire g13342;
  wire g13344;
  wire g13346;
  wire g13356;
  wire g13359;
  wire g13361;
  wire g13364;
  wire g13366;
  wire g13367;
  wire g13369;
  wire g13381;
  wire g13384;
  wire g13386;
  wire g13389;
  wire g1339;
  wire g13391;
  wire g13394;
  wire g13396;
  wire g13397;
  wire g134;
  wire g13405;
  wire g13406;
  wire g13407;
  wire g13408;
  wire g13409;
  wire g13410;
  wire g13411;
  wire g13412;
  wire g13413;
  wire g13414;
  wire g13415;
  wire g13416;
  wire g13417;
  wire g13418;
  wire g13419;
  wire g13420;
  wire g13421;
  wire g13422;
  wire g13423;
  wire g13424;
  wire g13425;
  wire g13426;
  wire g13427;
  wire g13428;
  wire g13429;
  wire g13430;
  wire g13431;
  wire g13432;
  wire g13433;
  wire g13434;
  wire g13435;
  wire g13436;
  wire g13437;
  wire g13438;
  wire g13439;
  wire g13440;
  wire g13441;
  wire g13442;
  wire g13443;
  wire g13444;
  wire g13445;
  wire g13446;
  wire g13447;
  wire g13448;
  wire g13449;
  wire g1345;
  wire g13450;
  wire g13451;
  wire g13452;
  wire g13453;
  wire g13454;
  wire g13455;
  wire g13456;
  wire g13457;
  wire g13458;
  wire g13459;
  wire g1346;
  wire g13460;
  wire g13461;
  wire g13462;
  wire g13463;
  wire g13464;
  wire g13465;
  wire g13466;
  wire g13467;
  wire g13468;
  wire g13469;
  wire g13475;
  wire g135;
  wire g1352;
  wire g13571;
  wire g13572;
  wire g13579;
  wire g1358;
  wire g13580;
  wire g13581;
  wire g13588;
  wire g13589;
  wire g13598;
  wire g13600;
  wire g13601;
  wire g13608;
  wire g13610;
  wire g13612;
  wire g13613;
  wire g13620;
  wire g13622;
  wire g13624;
  wire g13632;
  wire g13635;
  wire g13647;
  wire g1365;
  wire g13673;
  wire g1372;
  wire g1378;
  wire g138;
  wire g1384;
  wire g1385;
  wire g1386;
  wire g13863;
  wire g1387;
  wire g1388;
  wire g1389;
  wire g1390;
  wire g1391;
  wire g1392;
  wire g1393;
  wire g1394;
  wire g1395;
  wire g1396;
  wire g1397;
  wire g1398;
  wire g1399;
  wire g14;
  wire g1400;
  wire g1401;
  wire g1402;
  wire g1403;
  wire g1404;
  wire g1405;
  wire g1406;
  wire g1407;
  wire g1408;
  wire g1409;
  wire g141;
  wire g1410;
  wire g1411;
  wire g1412;
  wire g1413;
  wire g1414;
  wire g1415;
  wire g1416;
  wire g1417;
  wire g1418;
  wire g1419;
  wire g142;
  wire g1420;
  wire g1421;
  wire g1422;
  wire g1423;
  wire g1424;
  wire g1425;
  wire g1426;
  wire g143;
  wire g1430;
  wire g14337;
  wire g1435;
  wire g1439;
  wire g144;
  wire g1444;
  wire g1448;
  wire g145;
  wire g1453;
  wire g1457;
  wire g146;
  wire g1462;
  wire g1466;
  wire g14684;
  wire g147;
  wire g1471;
  wire g14718;
  wire g14745;
  wire g14746;
  wire g1476;
  wire g14764;
  wire g14765;
  wire g14766;
  wire g14774;
  wire g14775;
  wire g14794;
  wire g14795;
  wire g14796;
  wire g148;
  wire g1481;
  wire g14829;
  wire g14830;
  wire g1486;
  wire g14881;
  wire g14882;
  wire g14883;
  wire g14885;
  wire g149;
  wire g1491;
  wire g14954;
  wire g14955;
  wire g1496;
  wire g14966;
  wire g150;
  wire g1501;
  wire g15017;
  wire g15018;
  wire g15019;
  wire g15055;
  wire g1506;
  wire g15092;
  wire g151;
  wire g1511;
  wire g1512;
  wire g1513;
  wire g1514;
  wire g1515;
  wire g15151;
  wire g1516;
  wire g1517;
  wire g15170;
  wire g152;
  wire g1520;
  wire g1523;
  wire g1524;
  wire g1525;
  wire g1526;
  wire g1527;
  wire g1528;
  wire g1529;
  wire g153;
  wire g1530;
  wire g1531;
  wire g1532;
  wire g1533;
  wire g1534;
  wire g1535;
  wire g1536;
  wire g1537;
  wire g1538;
  wire g1539;
  wire g154;
  wire g1540;
  wire g1541;
  wire g1542;
  wire g1543;
  wire g1544;
  wire g1545;
  wire g1546;
  wire g1547;
  wire g155;
  wire g1550;
  wire g1551;
  wire g1552;
  wire g1553;
  wire g1554;
  wire g1555;
  wire g1556;
  wire g1557;
  wire g1558;
  wire g1559;
  wire g156;
  wire g1560;
  wire g1561;
  wire g1562;
  wire g1563;
  wire g1564;
  wire g1567;
  wire g157;
  wire g1570;
  wire g1573;
  wire g1576;
  wire g1579;
  wire g158;
  wire g1582;
  wire g1585;
  wire g15876;
  wire g1588;
  wire g159;
  wire g1591;
  wire g1594;
  wire g1597;
  wire g15989;
  wire g15991;
  wire g15994;
  wire g15997;
  wire g160;
  wire g1600;
  wire g16001;
  wire g16002;
  wire g16007;
  wire g16013;
  wire g16014;
  wire g16027;
  wire g1603;
  wire g16043;
  wire g16044;
  wire g1606;
  wire g16064;
  wire g1609;
  wire g16099;
  wire g161;
  wire g1612;
  wire g16132;
  wire g1615;
  wire g1618;
  wire g16181;
  wire g162;
  wire g1621;
  wire g1624;
  wire g1627;
  output g16297;
  wire g163;
  wire g1630;
  wire g1633;
  output g16355;
  wire g1636;
  wire g1639;
  output g16399;
  wire g164;
  wire g1642;
  output g16437;
  wire g1645;
  wire g16467;
  wire g16468;
  wire g16469;
  wire g16470;
  wire g16471;
  wire g16472;
  wire g16473;
  wire g16474;
  wire g16475;
  wire g16476;
  wire g16477;
  wire g16478;
  wire g16479;
  wire g1648;
  wire g16480;
  wire g16481;
  wire g16482;
  wire g16483;
  wire g16484;
  wire g16485;
  wire g16486;
  wire g16487;
  wire g16488;
  wire g16489;
  wire g16490;
  wire g16491;
  wire g16492;
  wire g16493;
  wire g16494;
  wire g16495;
  output g16496;
  wire g16497;
  wire g165;
  wire g16506;
  wire g1651;
  wire g16528;
  wire g1654;
  wire g16559;
  wire g16566;
  wire g1657;
  wire g1660;
  wire g1661;
  wire g1662;
  wire g1663;
  wire g1664;
  wire g1665;
  wire g16654;
  wire g1666;
  wire g1667;
  wire g16671;
  wire g1668;
  wire g1669;
  wire g16692;
  wire g1670;
  wire g1671;
  wire g16718;
  wire g1672;
  wire g1679;
  wire g168;
  wire g1680;
  wire g16802;
  wire g16803;
  wire g16813;
  wire g16823;
  wire g16824;
  wire g16831;
  wire g16835;
  wire g16843;
  wire g16844;
  wire g16845;
  wire g16849;
  wire g16851;
  wire g16853;
  wire g16854;
  wire g16857;
  wire g16858;
  wire g1686;
  wire g16860;
  wire g16861;
  wire g16862;
  wire g16863;
  wire g16866;
  wire g16877;
  wire g16878;
  wire g16880;
  wire g16881;
  wire g169;
  wire g1690;
  wire g16905;
  wire g16906;
  wire g16910;
  wire g1693;
  wire g16934;
  wire g1694;
  wire g16940;
  wire g1695;
  wire g1696;
  wire g1697;
  wire g16971;
  wire g1698;
  wire g1699;
  wire g17;
  wire g170;
  wire g1700;
  wire g1701;
  wire g1702;
  wire g1703;
  wire g1704;
  wire g1705;
  wire g1706;
  wire g171;
  wire g1712;
  wire g1718;
  wire g172;
  wire g17222;
  wire g17224;
  wire g17225;
  wire g17226;
  wire g17227;
  wire g17228;
  wire g17229;
  wire g1723;
  wire g17233;
  wire g17234;
  wire g17235;
  wire g17236;
  wire g1724;
  wire g17246;
  wire g17247;
  wire g17248;
  wire g17269;
  wire g1727;
  wire g17270;
  wire g17271;
  wire g173;
  wire g1730;
  wire g17300;
  wire g17302;
  wire g17303;
  wire g1731;
  wire g1732;
  wire g1733;
  wire g1734;
  wire g17340;
  wire g17341;
  wire g1735;
  wire g1738;
  wire g17383;
  wire g1739;
  wire g174;
  wire g1742;
  wire g17429;
  wire g17442;
  wire g1745;
  wire g1746;
  wire g1747;
  wire g1748;
  wire g1749;
  wire g175;
  wire g1750;
  wire g17500;
  wire g17503;
  wire g17523;
  wire g1753;
  wire g1754;
  wire g1757;
  wire g17570;
  wire g17591;
  wire g17594;
  wire g176;
  wire g1760;
  wire g1761;
  wire g17613;
  wire g1762;
  wire g1763;
  wire g1764;
  wire g17645;
  wire g1765;
  wire g17667;
  wire g1768;
  wire g17688;
  wire g1769;
  wire g17691;
  wire g177;
  wire g17710;
  wire g1772;
  wire g17746;
  wire g1775;
  wire g1776;
  wire g17767;
  wire g1777;
  wire g1778;
  wire g17788;
  wire g1779;
  wire g17791;
  wire g178;
  wire g1782;
  wire g1783;
  wire g1784;
  wire g17847;
  wire g1785;
  wire g1786;
  wire g17868;
  wire g1789;
  wire g179;
  wire g1792;
  wire g1795;
  wire g17959;
  wire g1798;
  wire g180;
  wire g1801;
  wire g1804;
  wire g1807;
  wire g1808;
  wire g1809;
  wire g181;
  wire g1810;
  wire g1813;
  wire g1816;
  wire g1819;
  wire g182;
  wire g1822;
  wire g1825;
  wire g1828;
  wire g1829;
  wire g1830;
  wire g1831;
  wire g1832;
  wire g1833;
  wire g1834;
  wire g1835;
  wire g1836;
  wire g1839;
  wire g1842;
  wire g1845;
  wire g1846;
  wire g1849;
  wire g185;
  wire g1852;
  wire g18542;
  wire g1855;
  wire g1858;
  wire g1859;
  wire g186;
  wire g1860;
  wire g1861;
  wire g1862;
  wire g1865;
  wire g1866;
  wire g18669;
  wire g1867;
  wire g18678;
  wire g1868;
  wire g1869;
  wire g1870;
  wire g18707;
  wire g1871;
  wire g18719;
  wire g18726;
  wire g1874;
  wire g18743;
  wire g18754;
  wire g18755;
  wire g18763;
  wire g1877;
  wire g18780;
  wire g18781;
  wire g18782;
  wire g18794;
  wire g1880;
  wire g18803;
  wire g18804;
  wire g18820;
  wire g18821;
  wire g18835;
  wire g18836;
  wire g18837;
  wire g18852;
  wire g1886;
  wire g18866;
  wire g18867;
  wire g18868;
  wire g1887;
  wire g18883;
  wire g18885;
  wire g189;
  wire g1890;
  wire g18906;
  wire g18907;
  wire g1893;
  wire g18942;
  wire g18957;
  wire g18968;
  wire g18975;
  wire g1900;
  wire g19000;
  wire g19012;
  wire g19021;
  wire g19022;
  wire g19023;
  wire g19024;
  wire g1903;
  wire g19033;
  wire g19034;
  wire g19035;
  wire g19036;
  wire g1904;
  wire g19045;
  wire g19046;
  wire g19047;
  wire g19048;
  wire g1905;
  wire g19057;
  wire g19058;
  wire g19059;
  wire g19060;
  wire g19061;
  wire g19062;
  wire g1908;
  wire g1909;
  wire g19096;
  wire g1910;
  wire g1911;
  wire g1912;
  wire g1913;
  wire g1914;
  wire g19144;
  wire g19145;
  wire g19147;
  wire g19149;
  wire g1915;
  wire g19151;
  wire g19152;
  wire g19153;
  wire g19154;
  wire g19156;
  wire g19157;
  wire g19158;
  wire g19159;
  wire g1916;
  wire g19162;
  wire g19163;
  wire g19164;
  wire g19167;
  wire g19168;
  wire g19169;
  wire g1917;
  wire g19170;
  wire g19172;
  wire g19173;
  wire g19174;
  wire g19175;
  wire g19176;
  wire g19178;
  wire g1918;
  wire g19180;
  wire g19182;
  wire g19183;
  wire g19184;
  wire g19185;
  wire g19189;
  wire g19190;
  wire g19196;
  wire g19197;
  wire g19198;
  wire g19199;
  wire g192;
  wire g19207;
  wire g19208;
  wire g1921;
  wire g19217;
  wire g19218;
  wire g1922;
  wire g19220;
  wire g19229;
  wire g1923;
  wire g19237;
  wire g19238;
  wire g19239;
  wire g1924;
  wire g19247;
  wire g19249;
  wire g1925;
  wire g19258;
  wire g19259;
  wire g19270;
  wire g1928;
  wire g1929;
  wire g1930;
  wire g1931;
  wire g1934;
  wire g1937;
  wire g1938;
  wire g1939;
  wire g1942;
  input g1943;
  wire g1944;
  wire g1945;
  wire g1946;
  wire g1947;
  wire g1948;
  wire g19484;
  wire g1949;
  wire g195;
  wire g1950;
  wire g19505;
  wire g1951;
  wire g1952;
  wire g19524;
  wire g1953;
  wire g19534;
  wire g1954;
  wire g19543;
  wire g19546;
  wire g1955;
  wire g19550;
  wire g19556;
  wire g1956;
  wire g19563;
  wire g1957;
  wire g19573;
  wire g19578;
  wire g1958;
  wire g1959;
  wire g19595;
  wire g19596;
  wire g1960;
  wire g19608;
  wire g1961;
  wire g1962;
  wire g19622;
  wire g1963;
  wire g1964;
  wire g19641;
  wire g1965;
  wire g19652;
  wire g1966;
  wire g1967;
  wire g19681;
  wire g19689;
  wire g19690;
  wire g19696;
  wire g1970;
  wire g19725;
  wire g1973;
  wire g19740;
  wire g1976;
  wire g19762;
  wire g19763;
  wire g19783;
  wire g1979;
  wire g19798;
  wire g198;
  wire g1982;
  wire g19825;
  wire g19830;
  wire g19838;
  wire g1985;
  wire g1988;
  wire g19893;
  wire g1991;
  wire g1994;
  wire g1997;
  wire g2;
  wire g20;
  wire g2000;
  wire g2003;
  wire g2006;
  wire g20082;
  wire g20083;
  wire g2009;
  wire g201;
  wire g2010;
  wire g20105;
  wire g2013;
  wire g20164;
  wire g20193;
  wire g20198;
  wire g2020;
  wire g20223;
  wire g20228;
  wire g20250;
  wire g20255;
  wire g2026;
  wire g20273;
  wire g20310;
  wire g20314;
  wire g2033;
  wire g20333;
  wire g20343;
  wire g20353;
  wire g20360;
  wire g20375;
  wire g20376;
  wire g20377;
  wire g2039;
  wire g20395;
  wire g20396;
  wire g204;
  wire g2040;
  wire g20417;
  wire g20418;
  wire g20419;
  wire g20439;
  wire g20440;
  wire g20441;
  wire g20457;
  wire g20458;
  wire g20459;
  wire g2046;
  wire g20469;
  wire g20470;
  wire g20471;
  wire g20478;
  wire g20479;
  wire g20484;
  wire g20485;
  wire g20491;
  wire g20497;
  wire g20498;
  wire g2052;
  wire g20555;
  wire g20556;
  wire g20557;
  wire g20558;
  wire g20559;
  wire g20560;
  wire g20561;
  wire g20562;
  wire g20563;
  wire g20564;
  wire g20565;
  wire g20566;
  wire g20567;
  wire g20568;
  wire g20569;
  wire g20570;
  wire g20571;
  wire g20572;
  wire g20573;
  wire g20574;
  wire g20575;
  wire g20576;
  wire g20577;
  wire g20578;
  wire g20579;
  wire g20580;
  wire g20581;
  wire g20582;
  wire g20583;
  wire g20584;
  wire g20585;
  wire g20586;
  wire g20587;
  wire g20588;
  wire g20589;
  wire g2059;
  wire g20590;
  wire g20591;
  wire g20592;
  wire g20593;
  wire g20594;
  wire g20595;
  wire g20596;
  wire g20597;
  wire g20598;
  wire g20599;
  wire g20600;
  wire g20601;
  wire g20602;
  wire g20603;
  wire g20604;
  wire g20605;
  wire g20606;
  wire g20607;
  wire g20608;
  wire g20609;
  wire g20610;
  wire g20611;
  wire g20612;
  wire g20613;
  wire g20614;
  wire g20615;
  wire g20616;
  wire g20617;
  wire g20618;
  wire g20619;
  wire g20620;
  wire g20621;
  wire g20622;
  wire g20623;
  wire g20624;
  wire g20625;
  wire g20626;
  wire g20627;
  wire g20628;
  wire g20629;
  wire g20630;
  wire g20631;
  wire g20632;
  wire g2066;
  wire g20682;
  wire g207;
  wire g20717;
  wire g2072;
  wire g20752;
  wire g2078;
  wire g20789;
  wire g2079;
  wire g2080;
  wire g2081;
  wire g2082;
  wire g20825;
  wire g2083;
  wire g2084;
  wire g2085;
  wire g2086;
  wire g2087;
  wire g20874;
  wire g20875;
  wire g20876;
  wire g20877;
  wire g20879;
  wire g2088;
  wire g20880;
  wire g20881;
  wire g20882;
  wire g20883;
  wire g20884;
  wire g2089;
  wire g20891;
  wire g20892;
  wire g20893;
  wire g20894;
  wire g20896;
  wire g20897;
  wire g20898;
  wire g20899;
  wire g2090;
  wire g20900;
  wire g20901;
  wire g20902;
  wire g20903;
  wire g2091;
  wire g20910;
  wire g20911;
  wire g20912;
  wire g20913;
  wire g20915;
  wire g20916;
  wire g20917;
  wire g20918;
  wire g20919;
  wire g2092;
  wire g20921;
  wire g20922;
  wire g20923;
  wire g20924;
  wire g20925;
  wire g20926;
  wire g20927;
  wire g2093;
  wire g20934;
  wire g20935;
  wire g20936;
  wire g20937;
  wire g20939;
  wire g2094;
  wire g20940;
  wire g20941;
  wire g20942;
  wire g20943;
  wire g20944;
  wire g20945;
  wire g20946;
  wire g20947;
  wire g20948;
  wire g20949;
  wire g2095;
  wire g20950;
  wire g20951;
  wire g20952;
  wire g20953;
  wire g20954;
  wire g20955;
  wire g2096;
  wire g20962;
  wire g20963;
  wire g20964;
  wire g20965;
  wire g20966;
  wire g20967;
  wire g20968;
  wire g20969;
  wire g2097;
  wire g20970;
  wire g20971;
  wire g20972;
  wire g20973;
  wire g20974;
  wire g20975;
  wire g20976;
  wire g20977;
  wire g20978;
  wire g20979;
  wire g2098;
  wire g20980;
  wire g20981;
  wire g20982;
  wire g20983;
  wire g20984;
  wire g20985;
  wire g20989;
  wire g2099;
  wire g20990;
  wire g20991;
  wire g20992;
  wire g20993;
  wire g20994;
  wire g20995;
  wire g20996;
  wire g20997;
  wire g20998;
  wire g20999;
  wire g210;
  wire g2100;
  wire g21000;
  wire g21001;
  wire g21002;
  wire g21003;
  wire g21004;
  wire g21005;
  wire g21006;
  wire g21007;
  wire g21009;
  wire g2101;
  wire g21010;
  wire g21011;
  wire g21015;
  wire g21016;
  wire g21017;
  wire g21018;
  wire g21019;
  wire g2102;
  wire g21020;
  wire g21021;
  wire g21022;
  wire g21023;
  wire g21024;
  wire g21025;
  wire g21026;
  wire g21027;
  wire g21028;
  wire g21029;
  wire g2103;
  wire g21030;
  wire g21031;
  wire g21032;
  wire g21033;
  wire g21034;
  wire g21035;
  wire g21039;
  wire g2104;
  wire g21040;
  wire g21041;
  wire g21042;
  wire g21043;
  wire g21044;
  wire g21045;
  wire g21046;
  wire g21047;
  wire g2105;
  wire g21050;
  wire g21051;
  wire g21052;
  wire g21053;
  wire g21054;
  wire g21055;
  wire g21056;
  wire g2106;
  wire g21060;
  wire g21061;
  wire g21062;
  wire g21063;
  wire g21064;
  wire g21069;
  wire g2107;
  wire g21070;
  wire g21071;
  wire g21072;
  wire g21073;
  wire g21074;
  wire g21075;
  wire g21079;
  wire g2108;
  wire g21080;
  wire g21081;
  wire g21082;
  wire g2109;
  wire g21093;
  wire g21094;
  wire g2110;
  wire g2111;
  wire g2112;
  wire g2113;
  wire g2114;
  wire g2115;
  wire g2116;
  wire g2117;
  wire g2118;
  wire g21187;
  wire g2119;
  wire g2120;
  wire g21202;
  wire g21217;
  wire g21225;
  wire g2124;
  wire g2129;
  wire g213;
  wire g21327;
  wire g2133;
  wire g21346;
  wire g21358;
  wire g21359;
  wire g21376;
  wire g21377;
  wire g2138;
  wire g21399;
  wire g2142;
  wire g21426;
  wire g21427;
  wire g21435;
  wire g21457;
  wire g2147;
  wire g21495;
  wire g21496;
  wire g2151;
  wire g21528;
  wire g21557;
  wire g2156;
  wire g216;
  wire g2160;
  wire g2165;
  wire g2170;
  wire g2175;
  wire g21795;
  wire g2180;
  wire g21824;
  wire g21842;
  wire g21843;
  wire g21845;
  wire g21847;
  wire g2185;
  wire g21851;
  wire g21878;
  wire g21880;
  wire g21882;
  wire g219;
  wire g2190;
  wire g21943;
  wire g21944;
  wire g21945;
  wire g21946;
  wire g21947;
  wire g21948;
  wire g21949;
  wire g2195;
  wire g21950;
  wire g21951;
  wire g21952;
  wire g21953;
  wire g21954;
  wire g21955;
  wire g21956;
  wire g21957;
  wire g21958;
  wire g21959;
  wire g21960;
  wire g21961;
  wire g21962;
  wire g21963;
  wire g21964;
  wire g21965;
  wire g21966;
  wire g21969;
  wire g21970;
  wire g21972;
  wire g21974;
  wire g21989;
  wire g2200;
  wire g22002;
  wire g22025;
  wire g22026;
  wire g22027;
  wire g22028;
  wire g22029;
  wire g22030;
  wire g22031;
  wire g22032;
  wire g22033;
  wire g22034;
  wire g22035;
  wire g22037;
  wire g22038;
  wire g22039;
  wire g22040;
  wire g22041;
  wire g22042;
  wire g22043;
  wire g22044;
  wire g22045;
  wire g22047;
  wire g22048;
  wire g22049;
  wire g2205;
  wire g22054;
  wire g22055;
  wire g22056;
  wire g22057;
  wire g22058;
  wire g22059;
  wire g2206;
  wire g22060;
  wire g22061;
  wire g22063;
  wire g22064;
  wire g22065;
  wire g22066;
  wire g22067;
  wire g22068;
  wire g2207;
  wire g22073;
  wire g22074;
  wire g22075;
  wire g22076;
  wire g22077;
  wire g22078;
  wire g22079;
  wire g2208;
  wire g22080;
  wire g22081;
  wire g22082;
  wire g22087;
  wire g22088;
  wire g22089;
  wire g2209;
  wire g22090;
  wire g22091;
  wire g22092;
  wire g22097;
  wire g22098;
  wire g22099;
  wire g2210;
  wire g22100;
  wire g22101;
  wire g22102;
  wire g22103;
  wire g22104;
  wire g22105;
  wire g22106;
  wire g22107;
  wire g2211;
  wire g22112;
  wire g22113;
  wire g22114;
  wire g22115;
  wire g22116;
  wire g22117;
  wire g22122;
  wire g22123;
  wire g22124;
  wire g22125;
  wire g22126;
  wire g22127;
  wire g22128;
  wire g22129;
  wire g22130;
  wire g22131;
  wire g22132;
  wire g22133;
  wire g22138;
  wire g22139;
  wire g2214;
  wire g22140;
  wire g22141;
  wire g22142;
  wire g22143;
  wire g22145;
  wire g22146;
  wire g22147;
  wire g22148;
  wire g22149;
  wire g22150;
  wire g22151;
  wire g22152;
  wire g22153;
  wire g22154;
  wire g22155;
  wire g22156;
  wire g22161;
  wire g22162;
  wire g22163;
  wire g22164;
  wire g22166;
  wire g22167;
  wire g22168;
  wire g22169;
  wire g2217;
  wire g22170;
  wire g22171;
  wire g22172;
  wire g22173;
  wire g22176;
  wire g22177;
  wire g22178;
  wire g22179;
  wire g2218;
  wire g22180;
  wire g22182;
  wire g22183;
  wire g22184;
  wire g22185;
  wire g2219;
  wire g22191;
  wire g22192;
  wire g22193;
  wire g22194;
  wire g222;
  wire g2220;
  wire g22200;
  wire g2221;
  wire g22218;
  wire g2222;
  wire g22225;
  wire g22226;
  wire g2223;
  wire g22231;
  wire g22234;
  wire g2224;
  wire g22242;
  wire g22247;
  wire g22249;
  wire g2225;
  wire g22253;
  wire g2226;
  wire g22263;
  wire g22267;
  wire g22269;
  wire g2227;
  wire g2228;
  wire g22280;
  wire g22284;
  wire g2229;
  wire g22299;
  wire g2230;
  wire g2231;
  wire g2232;
  wire g2233;
  wire g2234;
  wire g2235;
  wire g2236;
  wire g2237;
  wire g2238;
  wire g2239;
  wire g2240;
  wire g2241;
  wire g2244;
  wire g22444;
  wire g2245;
  wire g2246;
  wire g2247;
  wire g2248;
  wire g2249;
  wire g225;
  wire g2250;
  wire g2251;
  wire g22518;
  wire g22519;
  wire g2252;
  wire g2253;
  wire g2254;
  wire g22548;
  wire g22549;
  wire g2255;
  wire g22550;
  wire g22551;
  wire g22558;
  wire g22559;
  wire g2256;
  wire g2257;
  wire g22578;
  wire g2258;
  wire g22582;
  wire g22583;
  wire g22584;
  wire g22585;
  wire g22586;
  wire g22589;
  wire g22590;
  wire g22591;
  wire g22598;
  wire g22599;
  wire g2261;
  wire g22611;
  wire g22612;
  wire g22613;
  wire g22615;
  wire g22619;
  wire g22620;
  wire g22621;
  wire g22622;
  wire g22623;
  wire g22626;
  wire g22627;
  wire g22628;
  wire g22635;
  wire g22636;
  wire g22639;
  wire g2264;
  wire g22640;
  wire g22641;
  wire g22642;
  wire g22647;
  wire g22648;
  wire g22649;
  wire g22651;
  wire g22655;
  wire g22656;
  wire g22657;
  wire g22658;
  wire g22659;
  wire g22662;
  wire g22663;
  wire g22664;
  wire g22669;
  wire g2267;
  wire g22670;
  wire g22671;
  wire g22672;
  wire g22673;
  wire g22675;
  wire g22676;
  wire g22677;
  wire g22678;
  wire g22683;
  wire g22684;
  wire g22685;
  wire g22687;
  wire g22691;
  wire g22692;
  wire g22693;
  wire g22694;
  wire g22695;
  wire g2270;
  wire g22702;
  wire g22703;
  wire g22704;
  wire g22705;
  wire g22706;
  wire g22709;
  wire g22710;
  wire g22711;
  wire g22712;
  wire g22713;
  wire g22715;
  wire g22716;
  wire g22717;
  wire g22718;
  wire g22723;
  wire g22724;
  wire g22725;
  wire g22728;
  wire g22729;
  wire g2273;
  wire g22730;
  wire g22731;
  wire g22733;
  wire g22734;
  wire g22735;
  wire g22736;
  wire g22737;
  wire g22740;
  wire g22741;
  wire g22742;
  wire g22743;
  wire g22744;
  wire g22746;
  wire g22747;
  wire g22748;
  wire g22749;
  wire g22756;
  wire g22757;
  wire g22758;
  wire g2276;
  wire g22760;
  wire g22761;
  wire g22762;
  wire g22763;
  wire g22765;
  wire g22766;
  wire g22767;
  wire g22768;
  wire g22769;
  wire g22772;
  wire g22773;
  wire g22774;
  wire g22775;
  wire g22776;
  wire g22785;
  wire g22786;
  wire g2279;
  wire g22790;
  wire g22791;
  wire g22792;
  wire g22794;
  wire g22795;
  wire g22796;
  wire g22797;
  wire g22799;
  wire g228;
  wire g22800;
  wire g22801;
  wire g22802;
  wire g22803;
  wire g2282;
  wire g22824;
  wire g22827;
  wire g22828;
  wire g22832;
  wire g22833;
  wire g22834;
  wire g22836;
  wire g22837;
  wire g22838;
  wire g22839;
  wire g22840;
  wire g2285;
  wire g22864;
  wire g22866;
  wire g22867;
  wire g22871;
  wire g22872;
  wire g22873;
  wire g2288;
  wire g22899;
  wire g22901;
  wire g22902;
  wire g2291;
  wire g22934;
  wire g2294;
  wire g22945;
  wire g22948;
  wire g2297;
  wire g22970;
  wire g22979;
  wire g23;
  wire g2300;
  wire g23000;
  wire g23014;
  wire g23022;
  wire g2303;
  wire g23030;
  wire g23039;
  wire g23047;
  wire g23055;
  wire g23058;
  wire g2306;
  wire g23067;
  wire g23076;
  wire g23081;
  wire g2309;
  wire g23092;
  wire g23093;
  wire g23097;
  wire g231;
  wire g23110;
  wire g23111;
  wire g23114;
  wire g23116;
  wire g23117;
  wire g2312;
  wire g23123;
  wire g23124;
  wire g23126;
  wire g23132;
  wire g23133;
  wire g23136;
  wire g23137;
  wire g23148;
  wire g2315;
  wire g23154;
  wire g23159;
  wire g23160;
  wire g23161;
  wire g23162;
  wire g23163;
  wire g23164;
  wire g23165;
  wire g23166;
  wire g23167;
  wire g23168;
  wire g23169;
  wire g23170;
  wire g23171;
  wire g23172;
  wire g23173;
  wire g23174;
  wire g23175;
  wire g23176;
  wire g23177;
  wire g23178;
  wire g23179;
  wire g2318;
  wire g23180;
  wire g23181;
  wire g23182;
  wire g23183;
  wire g23184;
  wire g23185;
  wire g23186;
  wire g23187;
  wire g23188;
  wire g23189;
  wire g23190;
  wire g23191;
  wire g23192;
  wire g23193;
  wire g23194;
  wire g23195;
  wire g23196;
  wire g23197;
  wire g23198;
  wire g23199;
  wire g23200;
  wire g23201;
  wire g23202;
  wire g23203;
  wire g23204;
  wire g23205;
  wire g23206;
  wire g23207;
  wire g23208;
  wire g23209;
  wire g2321;
  wire g23210;
  wire g23211;
  wire g23212;
  wire g23213;
  wire g23214;
  wire g23215;
  wire g23216;
  wire g23217;
  wire g23218;
  wire g23219;
  wire g23220;
  wire g23221;
  wire g23222;
  wire g23223;
  wire g23224;
  wire g23225;
  wire g23226;
  wire g23227;
  wire g23228;
  wire g23229;
  wire g23230;
  wire g23231;
  wire g23232;
  wire g23233;
  wire g23234;
  wire g23235;
  wire g23236;
  wire g23237;
  wire g23238;
  wire g23239;
  wire g2324;
  wire g23240;
  wire g23241;
  wire g23242;
  wire g23243;
  wire g23244;
  wire g23245;
  wire g23246;
  wire g23247;
  wire g23248;
  wire g23249;
  wire g23250;
  wire g23251;
  wire g23252;
  wire g23253;
  wire g23254;
  wire g23255;
  wire g23256;
  wire g23257;
  wire g23258;
  wire g23259;
  wire g23260;
  wire g23261;
  wire g23262;
  wire g23263;
  wire g23264;
  wire g23265;
  wire g23266;
  wire g23267;
  wire g23268;
  wire g23269;
  wire g2327;
  wire g23270;
  wire g23271;
  wire g23272;
  wire g23273;
  wire g23274;
  wire g23275;
  wire g23276;
  wire g23277;
  wire g23278;
  wire g23279;
  wire g23280;
  wire g23281;
  wire g23282;
  wire g23283;
  wire g23284;
  wire g23285;
  wire g23286;
  wire g23287;
  wire g23288;
  wire g23289;
  wire g23290;
  wire g23291;
  wire g23292;
  wire g23293;
  wire g23294;
  wire g23295;
  wire g23296;
  wire g23297;
  wire g23298;
  wire g23299;
  wire g2330;
  wire g23300;
  wire g23301;
  wire g23302;
  wire g23303;
  wire g23304;
  wire g23305;
  wire g23306;
  wire g23307;
  wire g23308;
  wire g23309;
  wire g23310;
  wire g23311;
  wire g23312;
  wire g23313;
  wire g23314;
  wire g23315;
  wire g23316;
  wire g23317;
  wire g23318;
  wire g23324;
  wire g23329;
  wire g2333;
  wire g23330;
  wire g23339;
  wire g23348;
  wire g23357;
  wire g23358;
  wire g23359;
  wire g2336;
  wire g23385;
  wire g2339;
  wire g23392;
  wire g23399;
  wire g234;
  wire g23400;
  wire g23406;
  wire g23407;
  wire g23413;
  wire g23418;
  wire g2342;
  wire g23438;
  wire g23439;
  wire g2345;
  wire g23452;
  wire g23453;
  wire g23454;
  wire g23459;
  wire g23460;
  wire g23463;
  wire g23468;
  wire g23469;
  wire g23472;
  wire g2348;
  wire g23481;
  wire g23485;
  wire g23492;
  wire g23500;
  wire g23501;
  wire g23508;
  wire g2351;
  wire g23516;
  wire g23517;
  wire g23524;
  wire g23531;
  wire g23532;
  wire g2354;
  wire g23542;
  wire g23543;
  wire g23546;
  wire g23548;
  wire g23549;
  wire g2355;
  wire g23553;
  wire g23555;
  wire g23556;
  wire g23557;
  wire g2356;
  wire g23561;
  wire g23562;
  wire g23566;
  wire g23568;
  wire g23569;
  wire g2357;
  wire g23570;
  wire g23574;
  wire g23575;
  wire g23576;
  wire g2358;
  wire g23580;
  wire g23581;
  wire g23585;
  wire g23587;
  wire g23588;
  wire g23589;
  wire g2359;
  wire g23594;
  wire g23595;
  wire g23596;
  wire g23597;
  wire g2360;
  wire g23601;
  wire g23602;
  wire g23603;
  wire g23607;
  wire g23608;
  wire g2361;
  wire g23612;
  wire g23613;
  wire g23614;
  wire g23619;
  wire g2362;
  wire g23620;
  wire g23621;
  wire g23626;
  wire g23627;
  wire g23628;
  wire g23629;
  wire g2363;
  wire g23633;
  wire g23634;
  wire g23635;
  wire g2364;
  wire g23640;
  wire g23641;
  wire g23642;
  wire g2365;
  wire g2366;
  wire g23661;
  wire g23662;
  wire g23663;
  wire g23668;
  wire g23669;
  wire g23670;
  wire g23675;
  wire g23676;
  wire g23677;
  wire g23678;
  wire g23682;
  wire g23683;
  wire g23684;
  wire g23685;
  wire g23690;
  wire g23691;
  wire g23692;
  wire g237;
  wire g23711;
  wire g23712;
  wire g23713;
  wire g23718;
  wire g23719;
  wire g23720;
  wire g23725;
  wire g23727;
  wire g23728;
  wire g23729;
  wire g2373;
  wire g23730;
  wire g23736;
  wire g23737;
  wire g23738;
  wire g23739;
  wire g2374;
  wire g23744;
  wire g23745;
  wire g23746;
  wire g23765;
  wire g23766;
  wire g23767;
  wire g23773;
  wire g23774;
  wire g23775;
  wire g23782;
  wire g23783;
  wire g23784;
  wire g23785;
  wire g23791;
  wire g23792;
  wire g23793;
  wire g23794;
  wire g23799;
  wire g2380;
  wire g23800;
  wire g23801;
  wire g23821;
  wire g23826;
  wire g23827;
  wire g23828;
  wire g23835;
  wire g23836;
  wire g23837;
  wire g23838;
  wire g2384;
  wire g23844;
  wire g23845;
  wire g23846;
  wire g23847;
  wire g23856;
  wire g23861;
  wire g23862;
  wire g23863;
  wire g2387;
  wire g23870;
  wire g23871;
  wire g23872;
  wire g23873;
  wire g2388;
  wire g2389;
  wire g23890;
  wire g23895;
  wire g23896;
  wire g23897;
  wire g2390;
  wire g2391;
  wire g23911;
  wire g23916;
  wire g23919;
  wire g2392;
  wire g23923;
  wire g2393;
  wire g2394;
  wire g23943;
  wire g2395;
  wire g23955;
  wire g2396;
  wire g2397;
  wire g2398;
  wire g23984;
  wire g2399;
  wire g240;
  wire g2400;
  wire g24000;
  wire g24001;
  wire g24014;
  wire g24033;
  wire g24035;
  wire g24051;
  wire g24053;
  wire g24055;
  wire g24059;
  wire g2406;
  wire g24064;
  wire g24066;
  wire g24068;
  wire g24072;
  wire g24077;
  wire g24079;
  wire g24083;
  wire g24088;
  wire g24092;
  wire g2412;
  wire g2417;
  wire g24174;
  wire g24178;
  wire g24179;
  wire g2418;
  wire g24181;
  wire g24182;
  wire g24206;
  wire g24207;
  wire g24208;
  wire g24209;
  wire g2421;
  wire g24212;
  wire g24213;
  wire g24214;
  wire g24215;
  wire g24216;
  wire g24218;
  wire g24219;
  wire g24222;
  wire g24223;
  wire g24225;
  wire g24226;
  wire g24228;
  wire g24230;
  wire g24231;
  wire g24233;
  wire g24235;
  wire g24237;
  wire g24238;
  wire g2424;
  wire g24240;
  wire g24243;
  wire g24248;
  wire g2425;
  wire g24250;
  wire g24255;
  wire g24259;
  wire g2426;
  wire g24260;
  wire g24261;
  wire g24262;
  wire g24263;
  wire g24264;
  wire g24265;
  wire g24266;
  wire g24267;
  wire g24268;
  wire g24269;
  wire g2427;
  wire g24270;
  wire g24271;
  wire g24272;
  wire g24273;
  wire g24274;
  wire g24275;
  wire g24276;
  wire g24277;
  wire g24278;
  wire g24279;
  wire g2428;
  wire g24280;
  wire g24281;
  wire g24282;
  wire g24283;
  wire g24284;
  wire g24285;
  wire g24286;
  wire g24287;
  wire g24288;
  wire g24289;
  wire g2429;
  wire g24290;
  wire g24291;
  wire g24292;
  wire g24293;
  wire g24294;
  wire g24295;
  wire g24296;
  wire g24297;
  wire g24298;
  wire g24299;
  wire g243;
  wire g24300;
  wire g24301;
  wire g24302;
  wire g24303;
  wire g24304;
  wire g24305;
  wire g24306;
  wire g24307;
  wire g24308;
  wire g24309;
  wire g24310;
  wire g24311;
  wire g24312;
  wire g24313;
  wire g24314;
  wire g24315;
  wire g24316;
  wire g24317;
  wire g24318;
  wire g24319;
  wire g2432;
  wire g24320;
  wire g24321;
  wire g24322;
  wire g24323;
  wire g24324;
  wire g24325;
  wire g24326;
  wire g24327;
  wire g24328;
  wire g24329;
  wire g2433;
  wire g24330;
  wire g24331;
  wire g24332;
  wire g24333;
  wire g24334;
  wire g24335;
  wire g24336;
  wire g24337;
  wire g24338;
  wire g24339;
  wire g24340;
  wire g24341;
  wire g24342;
  wire g24343;
  wire g24344;
  wire g24345;
  wire g24346;
  wire g24347;
  wire g24348;
  wire g24349;
  wire g24350;
  wire g24351;
  wire g24352;
  wire g24353;
  wire g24354;
  wire g24355;
  wire g24356;
  wire g24357;
  wire g24358;
  wire g24359;
  wire g2436;
  wire g24360;
  wire g24361;
  wire g24362;
  wire g24363;
  wire g24364;
  wire g24365;
  wire g24366;
  wire g24367;
  wire g24368;
  wire g24369;
  wire g24370;
  wire g24371;
  wire g24372;
  wire g24373;
  wire g24374;
  wire g24375;
  wire g24376;
  wire g24377;
  wire g24378;
  wire g24379;
  wire g24380;
  wire g24381;
  wire g24382;
  wire g24383;
  wire g24384;
  wire g24385;
  wire g24386;
  wire g24387;
  wire g24388;
  wire g24389;
  wire g2439;
  wire g24390;
  wire g24391;
  wire g24392;
  wire g24393;
  wire g24394;
  wire g24395;
  wire g24396;
  wire g24397;
  wire g24398;
  wire g24399;
  wire g2440;
  wire g24400;
  wire g24401;
  wire g24402;
  wire g24403;
  wire g24404;
  wire g24405;
  wire g24406;
  wire g24407;
  wire g24408;
  wire g24409;
  wire g2441;
  wire g24410;
  wire g24411;
  wire g24412;
  wire g24413;
  wire g24414;
  wire g24415;
  wire g24416;
  wire g24417;
  wire g24418;
  wire g24419;
  wire g2442;
  wire g24420;
  wire g24421;
  wire g24422;
  wire g24423;
  wire g24424;
  wire g24425;
  wire g24426;
  wire g2443;
  wire g24430;
  wire g24434;
  wire g24438;
  wire g2444;
  wire g24445;
  wire g24446;
  wire g2447;
  wire g24473;
  wire g24476;
  wire g2448;
  wire g24491;
  wire g24498;
  wire g24499;
  wire g24501;
  wire g24507;
  wire g24508;
  wire g2451;
  wire g24510;
  wire g24511;
  wire g24513;
  wire g24518;
  wire g24519;
  wire g24521;
  wire g24522;
  wire g24524;
  wire g24525;
  wire g24527;
  wire g24531;
  wire g24532;
  wire g24534;
  wire g24535;
  wire g24537;
  wire g24538;
  wire g24539;
  wire g2454;
  wire g24544;
  wire g24545;
  wire g24547;
  wire g24548;
  wire g24549;
  wire g2455;
  wire g24551;
  wire g24556;
  wire g24557;
  wire g2456;
  wire g24560;
  wire g24562;
  wire g24567;
  wire g24568;
  wire g2457;
  wire g24570;
  wire g24572;
  wire g24576;
  wire g24577;
  wire g24579;
  wire g2458;
  wire g24581;
  wire g24582;
  wire g24583;
  wire g24584;
  wire g24586;
  wire g24587;
  wire g24588;
  wire g24589;
  wire g2459;
  wire g24592;
  wire g24593;
  wire g24594;
  wire g24597;
  wire g24598;
  wire g24599;
  wire g246;
  wire g24605;
  wire g24612;
  wire g2462;
  wire g2463;
  wire g2466;
  wire g2469;
  wire g2470;
  wire g2471;
  wire g2472;
  wire g2473;
  output g24734;
  wire g24735;
  wire g2476;
  wire g2477;
  wire g2478;
  wire g2479;
  wire g2480;
  wire g24816;
  wire g2483;
  wire g24835;
  wire g24851;
  wire g24856;
  wire g2486;
  wire g24865;
  wire g24872;
  wire g24879;
  wire g24886;
  wire g2489;
  wire g24890;
  wire g249;
  wire g24903;
  wire g24909;
  wire g2492;
  wire g24925;
  wire g24949;
  wire g2495;
  wire g24956;
  wire g24957;
  wire g2498;
  wire g2501;
  wire g2502;
  wire g25027;
  wire g2503;
  wire g2504;
  wire g25042;
  wire g25056;
  wire g25067;
  wire g2507;
  wire g2510;
  wire g25103;
  wire g25109;
  wire g25119;
  wire g25122;
  wire g2513;
  wire g25131;
  wire g25132;
  wire g25133;
  wire g25134;
  wire g25135;
  wire g25136;
  wire g25137;
  wire g25138;
  wire g25139;
  wire g25140;
  wire g25142;
  wire g25143;
  wire g25144;
  wire g25145;
  wire g25146;
  wire g25147;
  wire g25148;
  wire g25149;
  wire g25150;
  wire g25151;
  wire g25153;
  wire g25154;
  wire g25155;
  wire g25156;
  wire g25157;
  wire g25158;
  wire g25159;
  wire g2516;
  wire g25160;
  wire g25161;
  wire g25162;
  wire g25164;
  wire g25165;
  wire g25166;
  wire g25167;
  wire g25168;
  wire g25169;
  wire g25170;
  wire g25171;
  wire g25172;
  wire g25173;
  wire g25174;
  wire g25175;
  wire g25176;
  wire g25177;
  wire g25179;
  wire g25180;
  wire g25185;
  wire g25189;
  wire g2519;
  wire g25191;
  wire g25194;
  wire g25197;
  wire g25199;
  wire g252;
  wire g25201;
  wire g25202;
  wire g25204;
  wire g25206;
  wire g25207;
  wire g25209;
  wire g25211;
  wire g25212;
  wire g25213;
  wire g25214;
  wire g25215;
  wire g25217;
  wire g25218;
  wire g25219;
  wire g2522;
  wire g25220;
  wire g25221;
  wire g25222;
  wire g25223;
  wire g25224;
  wire g25225;
  wire g25227;
  wire g25228;
  wire g25229;
  wire g2523;
  wire g25230;
  wire g25231;
  wire g25232;
  wire g25233;
  wire g25234;
  wire g25235;
  wire g25236;
  wire g25237;
  wire g25239;
  wire g2524;
  wire g25240;
  wire g25241;
  wire g25242;
  wire g25243;
  wire g25244;
  wire g25245;
  wire g25246;
  wire g25247;
  wire g25248;
  wire g25249;
  wire g2525;
  wire g25250;
  wire g25251;
  wire g25252;
  wire g25253;
  wire g25255;
  wire g25256;
  wire g25257;
  wire g25259;
  wire g2526;
  wire g25260;
  wire g25262;
  wire g25263;
  wire g25265;
  wire g25266;
  wire g25267;
  wire g25268;
  wire g2527;
  wire g25270;
  wire g25271;
  wire g25272;
  wire g25279;
  wire g2528;
  wire g25280;
  wire g25288;
  wire g2529;
  wire g2530;
  wire g25327;
  wire g2533;
  wire g25336;
  wire g25350;
  wire g2536;
  wire g25364;
  wire g2539;
  wire g2540;
  output g25420;
  wire g25421;
  wire g2543;
  output g25435;
  wire g25436;
  output g25442;
  wire g25443;
  wire g25450;
  wire g25451;
  wire g25452;
  wire g2546;
  wire g25462;
  wire g25471;
  wire g25488;
  output g25489;
  wire g2549;
  wire g25490;
  wire g255;
  wire g25519;
  wire g2552;
  wire g25520;
  wire g2553;
  wire g2554;
  wire g2555;
  wire g2556;
  wire g25566;
  wire g25588;
  wire g2559;
  wire g2560;
  wire g2561;
  wire g2562;
  wire g2563;
  wire g2564;
  wire g25646;
  wire g25647;
  wire g2565;
  wire g25667;
  wire g2568;
  wire g25706;
  wire g25707;
  wire g2571;
  wire g25723;
  wire g25724;
  wire g2574;
  wire g25744;
  wire g25762;
  wire g25763;
  wire g25770;
  wire g25779;
  wire g25780;
  wire g25796;
  wire g25797;
  wire g258;
  wire g2580;
  wire g2581;
  wire g25817;
  wire g25824;
  wire g25833;
  wire g25834;
  wire g2584;
  wire g25850;
  wire g25851;
  wire g25859;
  wire g25868;
  wire g25869;
  wire g2587;
  wire g25880;
  wire g25886;
  wire g25891;
  wire g25932;
  wire g25935;
  wire g25938;
  wire g2594;
  wire g25940;
  wire g25952;
  wire g2597;
  wire g25976;
  wire g2598;
  wire g25982;
  wire g25983;
  wire g25984;
  wire g25985;
  wire g25986;
  wire g25987;
  wire g25988;
  wire g25989;
  wire g2599;
  wire g25990;
  wire g25991;
  wire g25992;
  wire g25993;
  wire g25994;
  wire g25995;
  wire g25996;
  wire g25997;
  wire g25998;
  wire g25999;
  wire g26;
  wire g26000;
  wire g26001;
  wire g26002;
  wire g26003;
  wire g26004;
  wire g26005;
  wire g26006;
  wire g26007;
  wire g26008;
  wire g26009;
  wire g26010;
  wire g26011;
  wire g26012;
  wire g26013;
  wire g26014;
  wire g26015;
  wire g26016;
  wire g26017;
  wire g26018;
  wire g26019;
  wire g2602;
  wire g26020;
  wire g26021;
  wire g26022;
  wire g26025;
  wire g2603;
  wire g26031;
  wire g26037;
  wire g2604;
  wire g26048;
  wire g2605;
  wire g2606;
  wire g2607;
  wire g2608;
  wire g26086;
  wire g2609;
  wire g261;
  wire g2610;
  wire g26102;
  output g26104;
  wire g26105;
  wire g26106;
  wire g2611;
  wire g26118;
  wire g2612;
  wire g26120;
  wire g26125;
  wire g26130;
  output g26135;
  wire g26136;
  wire g26144;
  output g26149;
  wire g2615;
  wire g26150;
  wire g26159;
  wire g2616;
  wire g26164;
  wire g26165;
  wire g26167;
  wire g2617;
  wire g26172;
  wire g26173;
  wire g26174;
  wire g2618;
  wire g26181;
  wire g26182;
  wire g26183;
  wire g26187;
  wire g26189;
  wire g2619;
  wire g26190;
  wire g26191;
  wire g26192;
  wire g26193;
  wire g26194;
  wire g26195;
  wire g26205;
  wire g26206;
  wire g26208;
  wire g26210;
  wire g26211;
  wire g26214;
  wire g26215;
  wire g26216;
  wire g2622;
  wire g26220;
  wire g26221;
  wire g26222;
  wire g26229;
  wire g2623;
  wire g26230;
  wire g26232;
  wire g26238;
  wire g26239;
  wire g2624;
  wire g26245;
  wire g26246;
  wire g26247;
  wire g26248;
  wire g26249;
  wire g2625;
  wire g26250;
  wire g26264;
  wire g26272;
  wire g26276;
  wire g26277;
  wire g2628;
  wire g26280;
  wire g26281;
  wire g26282;
  wire g26294;
  wire g26308;
  wire g2631;
  wire g26314;
  wire g26315;
  wire g2632;
  wire g2633;
  wire g26341;
  wire g26349;
  wire g26354;
  wire g26355;
  wire g2636;
  wire g26364;
  input g2637;
  wire g2638;
  wire g26385;
  wire g2639;
  wire g26398;
  wire g264;
  wire g2640;
  wire g26407;
  wire g2641;
  wire g2642;
  wire g26428;
  wire g2643;
  wire g26433;
  wire g26439;
  wire g2644;
  wire g26448;
  wire g2645;
  wire g2646;
  wire g26465;
  wire g2647;
  wire g26471;
  wire g2648;
  wire g26480;
  wire g26489;
  wire g2649;
  wire g26495;
  wire g26496;
  wire g2650;
  wire g26505;
  wire g26506;
  wire g26507;
  wire g2651;
  wire g2652;
  wire g26529;
  wire g2653;
  wire g26530;
  wire g26531;
  wire g26532;
  wire g26534;
  wire g2654;
  wire g26541;
  wire g26545;
  wire g26547;
  wire g26548;
  wire g2655;
  wire g26553;
  wire g26557;
  wire g26559;
  wire g2656;
  wire g26569;
  wire g2657;
  wire g26573;
  wire g26575;
  wire g26576;
  wire g26577;
  wire g2658;
  wire g2659;
  wire g26592;
  wire g26596;
  wire g2660;
  wire g2661;
  wire g26616;
  wire g26618;
  wire g2664;
  wire g26655;
  wire g26659;
  wire g26660;
  wire g26661;
  wire g26664;
  wire g26665;
  wire g26666;
  wire g26667;
  wire g26669;
  wire g2667;
  wire g26670;
  wire g26671;
  wire g26672;
  wire g26675;
  wire g26676;
  wire g26677;
  wire g26678;
  wire g26679;
  wire g26680;
  wire g26681;
  wire g26682;
  wire g26683;
  wire g26684;
  wire g26685;
  wire g26686;
  wire g26687;
  wire g26688;
  wire g26689;
  wire g26690;
  wire g26691;
  wire g26692;
  wire g26693;
  wire g26694;
  wire g26695;
  wire g26696;
  wire g26697;
  wire g26698;
  wire g26699;
  wire g267;
  wire g2670;
  wire g26700;
  wire g26701;
  wire g26702;
  wire g26703;
  wire g26704;
  wire g26705;
  wire g26706;
  wire g26707;
  wire g26708;
  wire g26709;
  wire g26710;
  wire g26711;
  wire g26712;
  wire g26713;
  wire g26714;
  wire g26715;
  wire g26716;
  wire g26717;
  wire g26718;
  wire g26719;
  wire g26720;
  wire g26721;
  wire g26722;
  wire g26723;
  wire g26724;
  wire g26725;
  wire g26726;
  wire g26727;
  wire g26728;
  wire g26729;
  wire g2673;
  wire g26730;
  wire g26731;
  wire g26732;
  wire g26733;
  wire g26734;
  wire g26735;
  wire g26736;
  wire g26737;
  wire g26738;
  wire g26739;
  wire g26740;
  wire g26741;
  wire g26742;
  wire g26743;
  wire g26744;
  wire g26745;
  wire g26746;
  wire g26747;
  wire g26748;
  wire g26749;
  wire g26750;
  wire g26751;
  wire g26752;
  wire g26753;
  wire g2676;
  wire g26776;
  wire g26781;
  wire g26786;
  wire g26789;
  wire g2679;
  wire g26795;
  wire g26798;
  wire g26803;
  wire g26804;
  wire g26805;
  wire g26806;
  wire g26807;
  wire g26808;
  wire g26809;
  wire g26810;
  wire g26811;
  wire g26812;
  wire g26813;
  wire g26814;
  wire g26815;
  wire g26816;
  wire g26817;
  wire g26818;
  wire g26819;
  wire g2682;
  wire g26820;
  wire g26821;
  wire g26822;
  wire g26823;
  wire g26824;
  wire g26825;
  wire g26826;
  wire g26827;
  wire g26828;
  wire g26830;
  wire g26831;
  wire g26832;
  wire g26834;
  wire g26836;
  wire g26840;
  wire g26843;
  wire g26844;
  wire g2685;
  wire g26850;
  wire g26852;
  wire g26858;
  wire g26864;
  wire g26868;
  wire g26872;
  wire g26875;
  wire g26876;
  wire g2688;
  wire g26881;
  wire g26883;
  wire g26884;
  wire g26886;
  wire g26890;
  wire g26895;
  wire g26896;
  wire g26900;
  wire g26909;
  wire g2691;
  wire g26910;
  wire g26921;
  wire g2694;
  wire g26953;
  wire g26954;
  wire g26956;
  wire g26957;
  wire g26959;
  wire g26960;
  wire g26964;
  wire g2697;
  wire g26974;
  wire g26983;
  wire g27;
  wire g270;
  wire g2700;
  wire g2703;
  wire g2704;
  wire g2707;
  wire g27075;
  wire g27102;
  wire g27116;
  wire g27120;
  wire g27123;
  wire g27126;
  wire g27129;
  wire g27131;
  wire g27132;
  wire g2714;
  wire g27140;
  wire g27145;
  wire g27150;
  wire g27156;
  wire g27158;
  wire g27166;
  wire g27168;
  wire g27183;
  wire g27189;
  wire g27190;
  wire g27191;
  wire g27192;
  wire g27193;
  wire g27194;
  wire g27195;
  wire g27196;
  wire g27197;
  wire g27198;
  wire g27199;
  wire g2720;
  wire g27200;
  wire g27206;
  wire g27207;
  wire g27208;
  wire g27209;
  wire g27210;
  wire g27211;
  wire g27212;
  wire g27217;
  wire g27218;
  wire g27219;
  wire g27220;
  wire g27221;
  wire g27222;
  wire g27223;
  wire g27224;
  wire g27225;
  wire g27226;
  wire g27227;
  wire g27228;
  wire g27229;
  wire g27230;
  wire g27231;
  wire g27232;
  wire g27233;
  wire g27234;
  wire g27235;
  wire g27236;
  wire g27237;
  wire g27238;
  wire g27239;
  wire g27243;
  wire g27253;
  wire g27255;
  wire g27256;
  wire g27257;
  wire g27258;
  wire g27259;
  wire g27260;
  wire g27261;
  wire g27262;
  wire g27263;
  wire g27264;
  wire g27265;
  wire g27266;
  wire g27267;
  wire g27268;
  wire g27269;
  wire g2727;
  wire g27270;
  wire g27271;
  wire g27272;
  wire g27273;
  wire g27274;
  wire g27275;
  wire g27276;
  wire g27277;
  wire g27278;
  wire g27279;
  wire g27280;
  wire g27281;
  wire g27282;
  wire g27283;
  wire g27284;
  wire g27285;
  wire g27286;
  wire g27287;
  wire g27288;
  wire g27289;
  wire g27290;
  wire g27291;
  wire g27292;
  wire g27293;
  wire g27294;
  wire g27295;
  wire g27296;
  wire g27297;
  wire g27298;
  wire g27299;
  wire g273;
  wire g27300;
  wire g27301;
  wire g27302;
  wire g27303;
  wire g27304;
  wire g27305;
  wire g27306;
  wire g27307;
  wire g27308;
  wire g27309;
  wire g27310;
  wire g27311;
  wire g27312;
  wire g27313;
  wire g27314;
  wire g27315;
  wire g27316;
  wire g27317;
  wire g27318;
  wire g27319;
  wire g27320;
  wire g27321;
  wire g27322;
  wire g27323;
  wire g27324;
  wire g27325;
  wire g27326;
  wire g27327;
  wire g27328;
  wire g27329;
  wire g2733;
  wire g27330;
  wire g27331;
  wire g27332;
  wire g27333;
  wire g27334;
  wire g27335;
  wire g27336;
  wire g27337;
  wire g27338;
  wire g27339;
  wire g2734;
  wire g27340;
  wire g27341;
  wire g27342;
  wire g27343;
  wire g27344;
  wire g27345;
  wire g27346;
  wire g27347;
  wire g27348;
  wire g27353;
  wire g27354;
  wire g27357;
  wire g27360;
  wire g27366;
  output g27380;
  wire g27381;
  wire g27383;
  wire g27384;
  wire g27385;
  wire g27386;
  wire g2740;
  wire g2746;
  wire g27463;
  wire g27479;
  wire g27480;
  wire g27483;
  wire g27493;
  wire g27494;
  wire g27497;
  wire g27502;
  wire g27503;
  wire g27505;
  wire g27508;
  wire g27514;
  wire g27515;
  wire g27517;
  wire g27522;
  wire g27523;
  wire g27525;
  wire g27526;
  wire g2753;
  wire g27533;
  wire g27539;
  wire g27540;
  wire g27542;
  wire g27547;
  wire g27548;
  wire g27553;
  wire g27559;
  wire g27560;
  wire g27562;
  wire g27569;
  wire g27586;
  wire g27589;
  wire g27594;
  wire g276;
  wire g2760;
  wire g27603;
  wire g27612;
  wire g27621;
  wire g2766;
  wire g27662;
  wire g27667;
  wire g27672;
  wire g27674;
  wire g27678;
  wire g27682;
  wire g27683;
  wire g27684;
  wire g27685;
  wire g27686;
  wire g27687;
  wire g27688;
  wire g27689;
  wire g27690;
  wire g27691;
  wire g27692;
  wire g27693;
  wire g27694;
  wire g27695;
  wire g27696;
  wire g27697;
  wire g27698;
  wire g27699;
  wire g27700;
  wire g27701;
  wire g27702;
  wire g27703;
  wire g27704;
  wire g27705;
  wire g27706;
  wire g27707;
  wire g27708;
  wire g27709;
  wire g27710;
  wire g27711;
  wire g27712;
  wire g27713;
  wire g27714;
  wire g27715;
  wire g27716;
  wire g27717;
  wire g27718;
  wire g2772;
  wire g27722;
  wire g27724;
  wire g2773;
  wire g2774;
  wire g2775;
  wire g27759;
  wire g2776;
  wire g27760;
  wire g27761;
  wire g27762;
  wire g27763;
  wire g27764;
  wire g27765;
  wire g27766;
  wire g27767;
  wire g27768;
  wire g27769;
  wire g2777;
  wire g27771;
  wire g2778;
  wire g27784;
  wire g27785;
  wire g27786;
  wire g2779;
  wire g27791;
  wire g27792;
  wire g27793;
  wire g27797;
  wire g27799;
  wire g2780;
  wire g27800;
  wire g27805;
  wire g2781;
  wire g2782;
  wire g2783;
  wire g2784;
  wire g2785;
  wire g2786;
  wire g2787;
  wire g2788;
  wire g2789;
  wire g279;
  wire g2790;
  wire g27903;
  wire g27905;
  wire g27907;
  wire g2791;
  wire g27910;
  wire g27912;
  wire g27918;
  wire g2792;
  wire g27927;
  wire g2793;
  wire g2794;
  wire g2795;
  wire g27955;
  wire g2796;
  wire g2797;
  wire g27971;
  wire g27972;
  wire g27976;
  wire g2798;
  wire g27986;
  wire g27987;
  wire g27988;
  wire g27989;
  wire g2799;
  wire g27992;
  wire g27993;
  wire g27998;
  wire g280;
  wire g2800;
  wire g28003;
  wire g28004;
  wire g28005;
  wire g28006;
  wire g28007;
  wire g2801;
  wire g28010;
  wire g28011;
  wire g28012;
  wire g28013;
  wire g28016;
  wire g28017;
  wire g2802;
  wire g28021;
  wire g28022;
  wire g28023;
  wire g28024;
  wire g28025;
  wire g28026;
  wire g2803;
  wire g28030;
  wire g28031;
  wire g28032;
  wire g28033;
  wire g28034;
  wire g28037;
  wire g28038;
  wire g28039;
  wire g2804;
  wire g28040;
  wire g28043;
  wire g28044;
  wire g28045;
  wire g28047;
  wire g28048;
  wire g28049;
  wire g2805;
  wire g28052;
  wire g28053;
  wire g28054;
  wire g28055;
  wire g28056;
  wire g2806;
  wire g28060;
  wire g28061;
  wire g28062;
  wire g28063;
  wire g28064;
  wire g28067;
  wire g28068;
  wire g28069;
  wire g2807;
  wire g28070;
  wire g28071;
  wire g28072;
  wire g28074;
  wire g28076;
  wire g28077;
  wire g28078;
  wire g2808;
  wire g28081;
  wire g28082;
  wire g28083;
  wire g28084;
  wire g28085;
  wire g28089;
  wire g2809;
  wire g28090;
  wire g28091;
  wire g28092;
  wire g28093;
  wire g28095;
  wire g28096;
  wire g28097;
  wire g28099;
  wire g281;
  wire g2810;
  wire g28101;
  wire g28102;
  wire g28103;
  wire g28106;
  wire g28107;
  wire g28108;
  wire g28109;
  wire g2811;
  wire g28110;
  wire g28113;
  wire g28114;
  wire g28115;
  wire g28117;
  wire g28119;
  wire g2812;
  wire g28120;
  wire g28121;
  wire g28124;
  wire g28125;
  wire g28126;
  wire g2813;
  wire g28132;
  wire g2814;
  wire g28145;
  wire g28146;
  wire g28147;
  wire g28148;
  wire g28149;
  wire g28151;
  wire g2817;
  wire g28179;
  wire g2818;
  wire g28194;
  wire g28199;
  wire g282;
  wire g28200;
  wire g28206;
  wire g28207;
  wire g28208;
  wire g28209;
  wire g2821;
  wire g28210;
  wire g28211;
  wire g28212;
  wire g28213;
  wire g28214;
  wire g28215;
  wire g28216;
  wire g28217;
  wire g28218;
  wire g28219;
  wire g28220;
  wire g28221;
  wire g28222;
  wire g28223;
  wire g28224;
  wire g28225;
  wire g28226;
  wire g28227;
  wire g28228;
  wire g28229;
  wire g28230;
  wire g28231;
  wire g28232;
  wire g28233;
  wire g28234;
  wire g28235;
  wire g28236;
  wire g28237;
  wire g28238;
  wire g28239;
  wire g2824;
  wire g28240;
  wire g28241;
  wire g28242;
  wire g28243;
  wire g28244;
  wire g28245;
  wire g28246;
  wire g28247;
  wire g28248;
  wire g28249;
  wire g28250;
  wire g28251;
  wire g28252;
  wire g28253;
  wire g28254;
  wire g28255;
  wire g28256;
  wire g28257;
  wire g28258;
  wire g28259;
  wire g28260;
  wire g28261;
  wire g28262;
  wire g28263;
  wire g28264;
  wire g28265;
  wire g28266;
  wire g28267;
  wire g28268;
  wire g28269;
  wire g2827;
  wire g28270;
  wire g28271;
  wire g28272;
  wire g28273;
  wire g28274;
  wire g28275;
  wire g28276;
  wire g28277;
  wire g28278;
  wire g28279;
  wire g28280;
  wire g28281;
  wire g28282;
  wire g28283;
  wire g28284;
  wire g28285;
  wire g28286;
  wire g28287;
  wire g28288;
  wire g28289;
  wire g28290;
  wire g28291;
  wire g28292;
  wire g28293;
  wire g28294;
  wire g28295;
  wire g28296;
  wire g28297;
  wire g28298;
  wire g28299;
  wire g283;
  wire g2830;
  wire g28300;
  wire g28301;
  wire g28302;
  wire g28303;
  wire g28304;
  wire g28305;
  wire g28306;
  wire g28307;
  wire g28308;
  wire g28309;
  wire g28310;
  wire g28311;
  wire g28312;
  wire g28313;
  wire g28314;
  wire g28315;
  wire g28316;
  wire g28317;
  wire g28318;
  wire g28321;
  wire g28325;
  wire g28328;
  wire g2833;
  wire g28341;
  wire g28342;
  wire g28343;
  wire g28344;
  wire g28345;
  wire g28346;
  wire g28347;
  wire g28348;
  wire g28349;
  wire g28350;
  wire g28351;
  wire g28352;
  wire g28353;
  wire g28354;
  wire g28355;
  wire g28356;
  wire g28357;
  wire g28358;
  wire g28359;
  wire g2836;
  wire g28360;
  wire g28361;
  wire g28362;
  wire g28363;
  wire g28364;
  wire g28365;
  wire g28366;
  wire g28367;
  wire g28368;
  wire g28369;
  wire g28370;
  wire g28371;
  wire g28372;
  wire g28374;
  wire g28375;
  wire g28377;
  wire g28382;
  wire g2839;
  wire g28390;
  wire g28393;
  wire g28395;
  wire g284;
  wire g28419;
  wire g2842;
  wire g28420;
  wire g28421;
  wire g28425;
  wire g28432;
  wire g28437;
  wire g28443;
  wire g28447;
  wire g2845;
  wire g28455;
  wire g28458;
  wire g28467;
  wire g2848;
  wire g28498;
  wire g285;
  wire g2851;
  wire g28524;
  wire g28526;
  wire g28527;
  wire g2854;
  wire g28552;
  wire g28553;
  wire g28555;
  wire g2857;
  wire g28579;
  wire g2858;
  wire g28580;
  wire g28583;
  wire g286;
  wire g28607;
  wire g2861;
  wire g28611;
  wire g28634;
  wire g28635;
  wire g28636;
  wire g28637;
  wire g28638;
  wire g2864;
  wire g28668;
  wire g2867;
  wire g28673;
  wire g28674;
  wire g28675;
  wire g28676;
  wire g28677;
  wire g28678;
  wire g28679;
  wire g28680;
  wire g28681;
  wire g28682;
  wire g28683;
  wire g28684;
  wire g28685;
  wire g28686;
  wire g28687;
  wire g28688;
  wire g28689;
  wire g28690;
  wire g28691;
  wire g28692;
  wire g28693;
  wire g28694;
  wire g28695;
  wire g28696;
  wire g28697;
  wire g28698;
  wire g28699;
  wire g287;
  wire g2870;
  wire g28700;
  wire g28701;
  wire g28702;
  wire g28703;
  wire g28704;
  wire g28705;
  wire g28706;
  wire g28720;
  wire g28721;
  wire g28723;
  wire g28725;
  wire g28727;
  wire g2873;
  wire g28730;
  wire g28732;
  wire g28734;
  wire g28735;
  wire g28736;
  wire g28738;
  wire g2874;
  wire g28740;
  wire g28744;
  wire g28745;
  wire g28746;
  wire g28747;
  wire g28749;
  wire g28754;
  wire g28758;
  wire g28759;
  wire g28760;
  wire g28761;
  wire g28763;
  wire g28767;
  wire g2877;
  wire g28771;
  wire g28772;
  wire g28773;
  wire g28774;
  wire g28778;
  wire g2878;
  wire g28782;
  wire g28783;
  wire g28788;
  wire g2879;
  wire g288;
  wire g2883;
  wire g28832;
  wire g28833;
  wire g28835;
  wire g28837;
  wire g28839;
  wire g2888;
  wire g28882;
  wire g28899;
  wire g289;
  wire g28903;
  wire g2892;
  wire g28924;
  wire g28950;
  wire g2896;
  wire g28990;
  wire g290;
  wire g2900;
  wire g2903;
  wire g29061;
  wire g29073;
  wire g29074;
  wire g29075;
  wire g2908;
  wire g29081;
  wire g29082;
  wire g29084;
  wire g29085;
  wire g29086;
  wire g29089;
  wire g29091;
  wire g29092;
  wire g29093;
  wire g29094;
  wire g29095;
  wire g29098;
  wire g29099;
  wire g291;
  wire g29100;
  wire g29101;
  wire g29102;
  wire g29104;
  wire g29105;
  wire g29106;
  wire g29108;
  wire g29109;
  wire g29110;
  wire g29111;
  wire g29112;
  wire g29113;
  wire g29117;
  wire g29118;
  wire g29119;
  wire g2912;
  wire g29120;
  wire g29131;
  wire g29132;
  wire g29133;
  wire g29134;
  wire g29135;
  wire g29136;
  wire g29137;
  wire g29138;
  wire g29139;
  wire g29140;
  wire g29141;
  wire g29142;
  wire g29143;
  wire g29144;
  wire g29145;
  wire g29146;
  wire g29147;
  wire g29148;
  wire g29149;
  wire g29150;
  wire g29151;
  wire g29152;
  wire g29153;
  wire g29154;
  wire g29155;
  wire g29156;
  wire g29157;
  wire g29158;
  wire g29159;
  wire g29160;
  wire g29161;
  wire g29162;
  wire g29163;
  wire g29164;
  wire g29165;
  wire g29166;
  wire g29167;
  wire g29169;
  wire g2917;
  wire g29170;
  wire g29172;
  wire g29173;
  wire g29178;
  wire g29179;
  wire g29181;
  wire g29182;
  wire g29184;
  wire g29185;
  wire g29187;
  wire g29192;
  wire g29194;
  wire g29197;
  wire g29198;
  wire g2920;
  wire g29201;
  wire g29204;
  wire g29205;
  wire g29209;
  wire g29212;
  wire g29213;
  wire g29218;
  wire g29221;
  wire g29226;
  wire g29230;
  wire g29237;
  wire g2924;
  wire g29244;
  wire g29246;
  wire g29249;
  wire g29253;
  wire g29258;
  wire g29267;
  wire g29270;
  wire g29273;
  wire g29276;
  wire g29278;
  wire g29279;
  wire g29281;
  wire g29288;
  wire g2929;
  wire g29293;
  wire g29297;
  wire g29298;
  wire g29299;
  wire g2930;
  wire g29304;
  wire g29305;
  wire g29306;
  wire g29307;
  wire g29308;
  wire g29309;
  wire g29311;
  wire g29314;
  wire g29315;
  wire g29316;
  wire g29317;
  wire g29318;
  wire g29319;
  wire g29322;
  wire g29325;
  wire g29326;
  wire g29327;
  wire g29328;
  wire g2933;
  wire g29331;
  wire g29334;
  wire g29335;
  wire g29339;
  wire g2934;
  wire g2935;
  wire g29350;
  wire g29353;
  wire g29354;
  wire g29355;
  wire g29356;
  wire g29357;
  wire g29358;
  wire g29359;
  wire g2938;
  wire g29401;
  wire g2941;
  wire g29412;
  wire g29413;
  wire g29414;
  wire g29415;
  wire g29416;
  wire g29417;
  wire g29418;
  wire g29419;
  wire g29420;
  wire g29421;
  wire g29422;
  wire g29423;
  wire g29424;
  wire g29425;
  wire g29426;
  wire g29427;
  wire g29428;
  wire g29434;
  wire g29435;
  wire g29436;
  wire g29437;
  wire g29438;
  wire g29439;
  wire g2944;
  wire g29440;
  wire g29445;
  wire g29446;
  wire g29447;
  wire g29448;
  wire g29449;
  wire g29450;
  wire g29451;
  wire g29452;
  wire g29453;
  wire g29454;
  wire g29455;
  wire g29456;
  wire g29457;
  wire g29458;
  wire g29459;
  wire g29460;
  wire g29461;
  wire g29462;
  wire g29463;
  wire g2947;
  wire g29495;
  wire g29496;
  wire g29497;
  wire g29499;
  wire g2950;
  wire g29501;
  wire g29504;
  wire g29506;
  wire g29507;
  wire g29508;
  wire g29509;
  wire g29510;
  wire g29511;
  wire g29512;
  wire g29513;
  wire g29514;
  wire g29515;
  wire g29516;
  wire g29517;
  wire g29519;
  wire g2953;
  wire g29530;
  wire g29535;
  wire g29537;
  wire g29542;
  wire g29544;
  wire g29546;
  wire g29551;
  wire g29554;
  wire g29556;
  wire g2956;
  wire g29561;
  wire g29563;
  wire g29568;
  wire g29579;
  wire g29580;
  wire g29581;
  wire g29582;
  wire g2959;
  wire g29606;
  wire g29608;
  wire g29609;
  wire g29611;
  wire g29612;
  wire g29613;
  wire g29616;
  wire g29617;
  wire g29618;
  wire g2962;
  wire g29620;
  wire g29621;
  wire g29623;
  wire g29627;
  wire g29628;
  wire g29629;
  wire g2963;
  wire g29630;
  wire g29631;
  wire g29632;
  wire g29633;
  wire g29634;
  wire g29635;
  wire g29636;
  wire g29637;
  wire g29638;
  wire g29639;
  wire g29640;
  wire g29641;
  wire g29642;
  wire g29643;
  wire g29644;
  wire g29645;
  wire g29646;
  wire g29647;
  wire g29648;
  wire g29649;
  wire g29650;
  wire g29651;
  wire g29652;
  wire g29653;
  wire g29654;
  wire g29655;
  wire g29656;
  wire g29657;
  wire g29658;
  wire g29659;
  wire g2966;
  wire g29660;
  wire g29661;
  wire g29662;
  wire g29664;
  wire g29666;
  wire g29668;
  wire g29689;
  wire g2969;
  wire g29690;
  wire g29691;
  wire g29692;
  wire g29693;
  wire g29694;
  wire g29695;
  wire g29696;
  wire g29697;
  wire g29698;
  wire g29699;
  wire g29700;
  wire g29701;
  wire g29702;
  wire g29704;
  wire g29708;
  wire g2972;
  wire g2975;
  wire g2978;
  wire g29794;
  wire g29795;
  wire g29796;
  wire g29797;
  wire g29798;
  wire g29799;
  wire g298;
  wire g29800;
  wire g29801;
  wire g29802;
  wire g29803;
  wire g29804;
  wire g29805;
  wire g29806;
  wire g29807;
  wire g29808;
  wire g29809;
  wire g2981;
  wire g2984;
  wire g29848;
  wire g2985;
  wire g2986;
  wire g2987;
  wire g299;
  wire g2990;
  wire g2991;
  wire g2992;
  wire g2993;
  wire g29932;
  wire g29933;
  wire g29934;
  wire g29935;
  wire g29936;
  wire g29937;
  wire g29938;
  wire g29939;
  wire g29940;
  wire g29941;
  wire g29943;
  wire g2997;
  wire g29972;
  wire g29973;
  wire g29974;
  wire g29975;
  wire g29976;
  wire g29977;
  wire g29978;
  wire g29979;
  wire g2998;
  wire g30;
  wire g3002;
  wire g30052;
  wire g30055;
  wire g3006;
  wire g30061;
  wire g30072;
  wire g30076;
  wire g30078;
  wire g30084;
  wire g3010;
  wire g30119;
  wire g30120;
  wire g30121;
  wire g30122;
  wire g30124;
  wire g3013;
  wire g3018;
  wire g30215;
  wire g3024;
  wire g30245;
  wire g30246;
  wire g30247;
  wire g30248;
  wire g30249;
  wire g30250;
  wire g30251;
  wire g30252;
  wire g30253;
  wire g30254;
  wire g30255;
  wire g30256;
  wire g30257;
  wire g30258;
  wire g30259;
  wire g30260;
  wire g30261;
  wire g30262;
  wire g30263;
  wire g30264;
  wire g30265;
  wire g30266;
  wire g30267;
  wire g30268;
  wire g30269;
  wire g30270;
  wire g30271;
  wire g30272;
  wire g30273;
  wire g30274;
  wire g30275;
  wire g30276;
  wire g30277;
  wire g30278;
  wire g30279;
  wire g3028;
  wire g30280;
  wire g30281;
  wire g30282;
  wire g30283;
  wire g30284;
  wire g30285;
  wire g30286;
  wire g30287;
  wire g30288;
  wire g30289;
  wire g30290;
  wire g30291;
  wire g30292;
  wire g30293;
  wire g30294;
  wire g30295;
  wire g30296;
  wire g30297;
  wire g30298;
  wire g30299;
  wire g30300;
  wire g30301;
  wire g30302;
  wire g30303;
  wire g30304;
  wire g30306;
  wire g30308;
  wire g30314;
  wire g3032;
  wire g30320;
  wire g30325;
  wire g30326;
  wire g30328;
  wire g30329;
  wire g30331;
  wire g30332;
  wire g30335;
  wire g30336;
  wire g30338;
  wire g30339;
  wire g30341;
  wire g30342;
  wire g30343;
  wire g30344;
  wire g30346;
  wire g30347;
  wire g30349;
  wire g30350;
  wire g30353;
  wire g30354;
  wire g30356;
  wire g30357;
  wire g30358;
  wire g30359;
  wire g3036;
  wire g30360;
  wire g30362;
  wire g30363;
  wire g30365;
  wire g30366;
  wire g30368;
  wire g30369;
  wire g30370;
  wire g30371;
  wire g30373;
  wire g30375;
  wire g30376;
  wire g30377;
  wire g30378;
  wire g30379;
  wire g30380;
  wire g30381;
  wire g30382;
  wire g3040;
  wire g30408;
  wire g3043;
  wire g30435;
  wire g30439;
  wire g3044;
  wire g30443;
  wire g30446;
  wire g3045;
  wire g30450;
  wire g30455;
  wire g30456;
  wire g30459;
  wire g3046;
  wire g30463;
  wire g30466;
  wire g30468;
  wire g3047;
  wire g30470;
  wire g30471;
  wire g30474;
  wire g30479;
  wire g3048;
  wire g30480;
  wire g30482;
  wire g30483;
  wire g30485;
  wire g30487;
  wire g30488;
  wire g3049;
  wire g30491;
  wire g30493;
  wire g30494;
  wire g30497;
  wire g30498;
  wire g305;
  wire g3050;
  wire g30500;
  wire g30501;
  wire g30503;
  wire g30505;
  wire g30506;
  wire g30507;
  wire g30508;
  wire g30509;
  wire g3051;
  wire g30510;
  wire g30511;
  wire g30512;
  wire g30513;
  wire g30514;
  wire g30515;
  wire g30516;
  wire g30517;
  wire g30518;
  wire g30519;
  wire g3052;
  wire g30520;
  wire g30521;
  wire g30522;
  wire g30523;
  wire g30524;
  wire g30525;
  wire g30526;
  wire g30527;
  wire g30528;
  wire g30529;
  wire g3053;
  wire g30530;
  wire g30531;
  wire g30532;
  wire g30533;
  wire g30534;
  wire g30535;
  wire g30536;
  wire g30537;
  wire g30538;
  wire g30539;
  wire g3054;
  wire g30540;
  wire g30541;
  wire g30542;
  wire g30543;
  wire g30544;
  wire g30545;
  wire g30546;
  wire g30547;
  wire g30548;
  wire g30549;
  wire g3055;
  wire g30550;
  wire g30551;
  wire g30552;
  wire g30553;
  wire g30554;
  wire g30555;
  wire g30556;
  wire g30557;
  wire g30558;
  wire g30559;
  wire g3056;
  wire g30560;
  wire g30561;
  wire g30562;
  wire g30563;
  wire g30564;
  wire g30565;
  wire g30566;
  wire g30567;
  wire g30568;
  wire g30569;
  wire g3057;
  wire g30570;
  wire g30571;
  wire g30572;
  wire g30573;
  wire g30574;
  wire g30578;
  wire g30579;
  wire g3058;
  wire g30580;
  wire g30581;
  wire g30582;
  wire g30583;
  wire g30585;
  wire g30586;
  wire g30587;
  wire g3059;
  wire g30591;
  wire g30592;
  wire g3060;
  wire g30600;
  wire g3061;
  wire g3062;
  wire g3063;
  wire g30635;
  wire g30636;
  wire g30637;
  wire g30638;
  wire g30639;
  wire g3064;
  wire g30640;
  wire g30641;
  wire g30642;
  wire g30643;
  wire g30644;
  wire g30645;
  wire g30646;
  wire g30647;
  wire g30648;
  wire g30649;
  wire g3065;
  wire g30650;
  wire g30651;
  wire g30652;
  wire g30653;
  wire g30654;
  wire g30655;
  wire g30656;
  wire g30657;
  wire g30658;
  wire g30659;
  wire g3066;
  wire g30660;
  wire g30661;
  wire g30662;
  wire g30663;
  wire g30664;
  wire g30665;
  wire g30666;
  wire g30667;
  wire g30668;
  wire g30669;
  wire g3067;
  wire g30670;
  wire g30671;
  wire g30672;
  wire g30673;
  wire g30674;
  wire g30675;
  wire g30676;
  wire g30677;
  wire g30678;
  wire g30679;
  wire g3068;
  wire g30680;
  wire g30681;
  wire g30682;
  wire g30683;
  wire g30684;
  wire g30686;
  wire g30687;
  wire g30688;
  wire g30689;
  wire g3069;
  wire g30690;
  wire g30691;
  wire g30692;
  wire g30693;
  wire g30694;
  wire g30695;
  wire g30699;
  wire g3070;
  wire g30700;
  wire g30701;
  wire g30702;
  wire g30703;
  wire g30704;
  wire g30705;
  wire g30706;
  wire g30707;
  wire g30708;
  wire g30709;
  wire g3071;
  wire g30710;
  wire g30711;
  wire g30712;
  wire g30713;
  wire g30714;
  wire g30715;
  wire g30716;
  wire g30717;
  wire g30718;
  wire g30719;
  wire g3072;
  wire g30720;
  wire g30721;
  wire g30722;
  wire g30723;
  wire g30724;
  wire g30725;
  wire g30726;
  wire g30727;
  wire g30729;
  wire g3073;
  wire g30730;
  wire g30731;
  wire g30732;
  wire g30733;
  wire g30734;
  wire g30737;
  wire g30738;
  wire g30739;
  wire g3074;
  wire g30740;
  wire g30741;
  wire g30742;
  wire g30745;
  wire g30746;
  wire g30747;
  wire g30748;
  wire g30749;
  wire g3075;
  wire g30751;
  wire g30752;
  wire g30753;
  wire g30756;
  wire g3076;
  wire g30765;
  wire g30767;
  wire g30769;
  wire g3077;
  wire g30770;
  wire g30772;
  wire g30773;
  wire g30774;
  wire g30776;
  wire g30777;
  wire g30778;
  wire g3078;
  wire g30781;
  wire g30782;
  wire g30784;
  wire g3079;
  wire g30792;
  wire g30793;
  wire g30794;
  wire g30795;
  wire g30796;
  wire g30797;
  wire g30798;
  wire g30799;
  wire g3080;
  wire g30800;
  wire g30801;
  wire g30802;
  wire g30803;
  wire g30804;
  wire g30805;
  wire g30806;
  wire g30807;
  wire g30808;
  wire g30809;
  wire g30810;
  wire g30811;
  wire g30812;
  wire g30813;
  wire g30814;
  wire g30815;
  wire g30816;
  wire g30817;
  wire g30818;
  wire g30819;
  wire g30820;
  wire g30821;
  wire g30822;
  wire g30823;
  wire g30824;
  wire g30825;
  wire g30826;
  wire g30827;
  wire g30828;
  wire g30829;
  wire g3083;
  wire g30830;
  wire g30831;
  wire g30832;
  wire g30833;
  wire g30834;
  wire g30835;
  wire g30836;
  wire g30837;
  wire g30838;
  wire g30839;
  wire g3084;
  wire g30840;
  wire g30841;
  wire g30842;
  wire g30843;
  wire g30844;
  wire g30845;
  wire g30846;
  wire g30847;
  wire g30848;
  wire g30849;
  wire g3085;
  wire g30850;
  wire g30851;
  wire g30852;
  wire g30853;
  wire g30854;
  wire g30855;
  wire g30856;
  wire g30857;
  wire g30858;
  wire g30859;
  wire g3086;
  wire g30860;
  wire g30861;
  wire g30862;
  wire g30863;
  wire g30864;
  wire g30865;
  wire g30866;
  wire g30867;
  wire g30868;
  wire g30869;
  wire g3087;
  wire g30870;
  wire g30871;
  wire g30872;
  wire g30873;
  wire g30874;
  wire g30875;
  wire g30876;
  wire g30877;
  wire g30878;
  wire g30879;
  wire g3088;
  wire g30880;
  wire g30881;
  wire g30882;
  wire g30883;
  wire g30884;
  wire g30885;
  wire g30886;
  wire g30887;
  wire g30888;
  wire g30889;
  wire g30890;
  wire g30891;
  wire g30892;
  wire g30893;
  wire g30894;
  wire g30895;
  wire g30896;
  wire g30897;
  wire g30898;
  wire g30899;
  wire g309;
  wire g30900;
  wire g30901;
  wire g30902;
  wire g30903;
  wire g30904;
  wire g30905;
  wire g30906;
  wire g30907;
  wire g30908;
  wire g30909;
  wire g3091;
  wire g30910;
  wire g30911;
  wire g30912;
  wire g30913;
  wire g30914;
  wire g30915;
  wire g3092;
  wire g30928;
  wire g3093;
  wire g30937;
  wire g30938;
  wire g30939;
  wire g3094;
  wire g30940;
  wire g30941;
  wire g30942;
  wire g30943;
  wire g3095;
  wire g3096;
  wire g30962;
  wire g30963;
  wire g30964;
  wire g30965;
  wire g30966;
  wire g30967;
  wire g30968;
  wire g30969;
  wire g3097;
  wire g30971;
  wire g30972;
  wire g30973;
  wire g30974;
  wire g30975;
  wire g30976;
  wire g30977;
  wire g30978;
  wire g30979;
  wire g3098;
  wire g30980;
  wire g30981;
  wire g30982;
  wire g30983;
  wire g30984;
  wire g30985;
  wire g30986;
  wire g30987;
  wire g30988;
  wire g30989;
  wire g3099;
  wire g3100;
  wire g3101;
  wire g3102;
  wire g3103;
  wire g3104;
  wire g3105;
  wire g3106;
  wire g3107;
  wire g3108;
  wire g3109;
  wire g3110;
  wire g3111;
  wire g3112;
  wire g3113;
  wire g3114;
  wire g3117;
  wire g312;
  wire g3120;
  wire g3123;
  wire g3124;
  wire g3125;
  wire g3126;
  wire g3127;
  wire g3128;
  wire g3129;
  wire g313;
  wire g3132;
  wire g3133;
  wire g3134;
  wire g3135;
  wire g3136;
  wire g3139;
  wire g314;
  wire g3142;
  wire g3147;
  wire g315;
  wire g3151;
  wire g3155;
  wire g3158;
  wire g316;
  wire g3161;
  wire g3164;
  wire g3167;
  wire g317;
  wire g3170;
  wire g3173;
  wire g3176;
  wire g3179;
  wire g318;
  wire g3182;
  wire g3185;
  wire g3188;
  wire g319;
  wire g3191;
  wire g3194;
  wire g3197;
  wire g3198;
  wire g320;
  wire g3201;
  wire g3204;
  wire g3207;
  wire g321;
  wire g3210;
  wire g3211;
  input g3212;
  input g3213;
  input g3214;
  input g3215;
  input g3216;
  input g3217;
  input g3218;
  input g3219;
  wire g322;
  input g3220;
  input g3221;
  input g3222;
  input g3223;
  input g3224;
  input g3225;
  input g3226;
  input g3227;
  input g3228;
  input g3229;
  wire g323;
  input g3230;
  input g3231;
  input g3232;
  input g3233;
  input g3234;
  wire g3235;
  wire g3236;
  wire g3237;
  wire g3238;
  wire g3239;
  wire g324;
  wire g3240;
  wire g3241;
  wire g3242;
  wire g3243;
  wire g3244;
  wire g3245;
  wire g3246;
  wire g3247;
  wire g3248;
  wire g3249;
  wire g325;
  wire g3250;
  wire g3251;
  wire g3252;
  wire g3253;
  wire g3254;
  wire g33;
  wire g3306;
  wire g331;
  wire g3338;
  wire g3366;
  wire g337;
  wire g3398;
  wire g3410;
  wire g342;
  wire g343;
  wire g346;
  wire g3462;
  wire g349;
  wire g3494;
  wire g350;
  wire g351;
  wire g352;
  wire g3522;
  wire g353;
  wire g354;
  wire g3554;
  wire g3566;
  wire g357;
  wire g358;
  wire g36;
  wire g361;
  wire g3618;
  wire g364;
  wire g365;
  wire g3650;
  wire g366;
  wire g367;
  wire g3678;
  wire g368;
  wire g369;
  wire g3710;
  wire g372;
  wire g3722;
  wire g373;
  wire g376;
  wire g3774;
  wire g379;
  wire g380;
  wire g3806;
  wire g381;
  wire g382;
  wire g383;
  wire g3834;
  wire g384;
  wire g3866;
  wire g387;
  wire g3878;
  wire g388;
  wire g39;
  wire g3900;
  wire g391;
  wire g394;
  wire g395;
  wire g396;
  wire g397;
  wire g398;
  output g3993;
  wire g401;
  wire g402;
  wire g403;
  wire g404;
  wire g405;
  wire g408;
  output g4088;
  output g4090;
  wire g411;
  wire g414;
  wire g417;
  wire g42;
  wire g420;
  output g4200;
  wire g423;
  wire g426;
  wire g427;
  wire g428;
  wire g429;
  wire g432;
  output g4321;
  output g4323;
  wire g4338;
  wire g4339;
  wire g435;
  wire g438;
  wire g441;
  wire g444;
  output g4450;
  wire g447;
  wire g448;
  wire g449;
  wire g45;
  wire g450;
  wire g4507;
  wire g4508;
  wire g451;
  wire g452;
  wire g453;
  wire g454;
  wire g455;
  wire g458;
  output g4590;
  wire g461;
  wire g464;
  wire g465;
  wire g468;
  wire g4683;
  wire g4684;
  wire g471;
  wire g4735;
  wire g4736;
  wire g474;
  wire g477;
  wire g478;
  wire g479;
  wire g48;
  wire g480;
  wire g481;
  wire g484;
  wire g485;
  wire g486;
  wire g4860;
  wire g4861;
  wire g487;
  wire g488;
  wire g489;
  wire g490;
  wire g4911;
  wire g4912;
  wire g493;
  wire g496;
  wire g499;
  wire g5;
  wire g506;
  wire g507;
  wire g5070;
  wire g5071;
  input g51;
  wire g510;
  wire g513;
  wire g5141;
  wire g5199;
  wire g52;
  wire g520;
  wire g5200;
  wire g523;
  wire g5234;
  wire g524;
  wire g525;
  wire g528;
  wire g529;
  wire g5297;
  wire g530;
  wire g531;
  wire g532;
  wire g533;
  wire g5334;
  wire g534;
  wire g535;
  wire g536;
  wire g537;
  wire g538;
  output g5388;
  wire g5390;
  wire g5395;
  wire g5396;
  wire g5397;
  wire g5398;
  wire g5399;
  wire g5400;
  wire g5401;
  wire g5402;
  wire g5403;
  wire g5404;
  wire g5405;
  wire g5406;
  wire g5407;
  wire g5408;
  wire g5409;
  wire g541;
  wire g5411;
  wire g5412;
  wire g5413;
  wire g5414;
  wire g5415;
  wire g5416;
  wire g5417;
  wire g5418;
  wire g5419;
  wire g542;
  wire g5420;
  wire g5421;
  wire g5422;
  wire g5424;
  wire g5425;
  wire g5426;
  wire g5427;
  wire g543;
  output g5437;
  wire g5438;
  wire g544;
  wire g545;
  output g5472;
  wire g5473;
  wire g548;
  wire g549;
  wire g550;
  wire g5508;
  wire g551;
  output g5511;
  wire g5512;
  wire g554;
  wire g5547;
  wire g5548;
  output g5549;
  wire g5550;
  wire g5552;
  output g5555;
  wire g5556;
  wire g557;
  wire g558;
  wire g559;
  wire g5593;
  wire g5594;
  output g5595;
  wire g5596;
  wire g5598;
  wire g56;
  wire g5610;
  wire g5611;
  output g5612;
  wire g5613;
  wire g5615;
  wire g562;
  wire g5626;
  wire g5627;
  output g5629;
  input g563;
  wire g5635;
  wire g5636;
  output g5637;
  wire g5638;
  wire g564;
  wire g5645;
  output g5648;
  wire g565;
  wire g5654;
  wire g5655;
  output g5657;
  wire g566;
  wire g5665;
  wire g567;
  wire g568;
  wire g5683;
  output g5686;
  wire g569;
  wire g5692;
  wire g5693;
  output g5695;
  wire g570;
  wire g5701;
  wire g5703;
  wire g5707;
  wire g571;
  wire g5713;
  wire g5717;
  wire g572;
  wire g573;
  wire g5735;
  output g5738;
  wire g574;
  wire g5744;
  wire g5745;
  output g5747;
  wire g5749;
  wire g575;
  wire g5752;
  wire g576;
  wire g5761;
  wire g5765;
  wire g577;
  wire g5771;
  wire g5775;
  wire g578;
  wire g579;
  wire g5793;
  output g5796;
  wire g5799;
  wire g580;
  wire g5800;
  wire g5801;
  wire g5803;
  wire g581;
  wire g5811;
  wire g582;
  wire g5820;
  wire g5824;
  wire g583;
  wire g5830;
  wire g5834;
  wire g584;
  wire g5849;
  wire g585;
  wire g5850;
  wire g5852;
  wire g5856;
  wire g5859;
  wire g586;
  wire g5867;
  wire g587;
  wire g5876;
  wire g5880;
  wire g5886;
  wire g5889;
  wire g5893;
  wire g5899;
  wire g590;
  wire g5903;
  wire g5906;
  wire g5914;
  wire g5922;
  wire g5923;
  wire g5924;
  wire g593;
  wire g5932;
  wire g5938;
  wire g5942;
  wire g5945;
  wire g5951;
  wire g5952;
  wire g5953;
  wire g5958;
  wire g596;
  wire g5966;
  wire g5972;
  wire g5976;
  wire g5978;
  wire g5979;
  wire g5982;
  wire g5987;
  wire g599;
  wire g5995;
  wire g6000;
  wire g6014;
  wire g6015;
  wire g6019;
  wire g602;
  wire g6024;
  wire g6029;
  wire g6030;
  wire g6031;
  wire g6035;
  wire g6040;
  wire g6041;
  wire g6042;
  wire g6046;
  wire g6048;
  wire g605;
  wire g6051;
  wire g6052;
  wire g6053;
  wire g6054;
  wire g6055;
  wire g6056;
  wire g6057;
  wire g6058;
  wire g6059;
  wire g6060;
  wire g6061;
  wire g6062;
  wire g6063;
  wire g6064;
  wire g6065;
  wire g6066;
  wire g6067;
  wire g6079;
  wire g608;
  wire g6080;
  wire g6081;
  wire g6082;
  wire g6083;
  wire g6084;
  wire g6085;
  wire g6086;
  wire g6098;
  wire g6099;
  wire g61;
  wire g6100;
  wire g6101;
  wire g6102;
  wire g6103;
  wire g611;
  wire g6115;
  wire g6116;
  wire g6117;
  wire g6118;
  wire g6130;
  wire g6131;
  wire g6134;
  wire g6135;
  wire g6139;
  wire g614;
  wire g6145;
  wire g6153;
  wire g6156;
  wire g6166;
  wire g617;
  wire g6183;
  wire g6193;
  wire g620;
  wire g6204;
  wire g6215;
  output g6225;
  wire g623;
  wire g6230;
  output g6231;
  wire g6232;
  wire g626;
  wire g6288;
  wire g629;
  wire g6293;
  wire g630;
  wire g6304;
  output g6313;
  wire g6314;
  wire g633;
  wire g6367;
  output g6368;
  wire g6369;
  wire g640;
  wire g6425;
  wire g6430;
  wire g6441;
  output g6442;
  output g6447;
  wire g6448;
  wire g646;
  output g6485;
  wire g6486;
  wire g65;
  wire g6517;
  output g6518;
  wire g6519;
  wire g653;
  wire g6572;
  output g6573;
  wire g6574;
  wire g659;
  wire g660;
  wire g6630;
  wire g6635;
  wire g6636;
  wire g6641;
  output g6642;
  wire g6643;
  wire g666;
  output g6677;
  wire g6678;
  wire g6711;
  output g6712;
  wire g6713;
  wire g672;
  output g6750;
  wire g6751;
  wire g6781;
  output g6782;
  wire g6783;
  wire g679;
  wire g6836;
  output g6837;
  wire g6838;
  wire g686;
  wire g6894;
  output g6895;
  wire g6897;
  output g6911;
  wire g6912;
  wire g692;
  wire g6942;
  wire g6943;
  output g6944;
  wire g6945;
  output g6979;
  wire g698;
  wire g6980;
  wire g699;
  wire g70;
  wire g700;
  wire g701;
  wire g7013;
  output g7014;
  wire g7015;
  wire g702;
  wire g703;
  wire g704;
  wire g705;
  output g7052;
  wire g7053;
  wire g706;
  wire g707;
  wire g708;
  wire g7083;
  output g7084;
  wire g7085;
  wire g709;
  wire g710;
  wire g711;
  wire g712;
  wire g713;
  wire g7138;
  wire g7139;
  wire g714;
  wire g7140;
  wire g7141;
  wire g715;
  wire g7157;
  wire g716;
  output g7161;
  wire g7162;
  wire g717;
  wire g718;
  wire g719;
  wire g7192;
  wire g7193;
  output g7194;
  wire g7195;
  wire g720;
  wire g721;
  wire g722;
  output g7229;
  wire g723;
  wire g7230;
  wire g724;
  wire g725;
  wire g726;
  wire g7263;
  output g7264;
  wire g7265;
  wire g727;
  wire g728;
  wire g729;
  wire g730;
  output g7302;
  wire g7303;
  wire g731;
  wire g732;
  wire g733;
  wire g7333;
  output g7334;
  wire g7336;
  wire g7337;
  wire g734;
  wire g7346;
  wire g7348;
  wire g735;
  wire g7353;
  output g7357;
  wire g7358;
  wire g736;
  wire g737;
  wire g738;
  wire g7388;
  wire g7389;
  wire g739;
  output g7390;
  wire g7391;
  wire g74;
  wire g740;
  output g7425;
  wire g7426;
  wire g744;
  wire g7459;
  wire g7460;
  wire g7461;
  wire g7476;
  wire g7478;
  wire g7483;
  output g7487;
  wire g7488;
  wire g749;
  wire g7518;
  output g7519;
  wire g7521;
  wire g753;
  wire g7532;
  wire g7534;
  wire g7539;
  wire g7540;
  wire g7541;
  wire g7554;
  wire g7558;
  wire g7560;
  wire g7561;
  wire g7577;
  wire g758;
  wire g7581;
  wire g7582;
  wire g7591;
  wire g7594;
  wire g7606;
  wire g762;
  wire g767;
  wire g771;
  wire g776;
  wire g780;
  wire g785;
  wire g789;
  wire g79;
  wire g7901;
  output g7909;
  wire g7911;
  wire g793;
  wire g7936;
  output g7956;
  output g7961;
  wire g7963;
  wire g797;
  wire g7976;
  wire g8;
  output g8007;
  wire g801;
  output g8012;
  wire g8014;
  output g8021;
  output g8023;
  output g8030;
  wire g8031;
  wire g805;
  output g8082;
  output g8087;
  wire g8089;
  wire g809;
  output g8096;
  output g8106;
  wire g8107;
  wire g813;
  output g8167;
  wire g817;
  output g8175;
  wire g818;
  wire g819;
  wire g820;
  wire g821;
  wire g822;
  wire g823;
  output g8249;
  output g8251;
  output g8258;
  output g8259;
  wire g826;
  output g8260;
  output g8261;
  output g8262;
  output g8263;
  output g8264;
  output g8265;
  output g8266;
  output g8267;
  output g8268;
  output g8269;
  output g8270;
  output g8271;
  output g8272;
  output g8273;
  output g8274;
  output g8275;
  wire g8277;
  wire g8278;
  wire g8284;
  wire g8285;
  wire g8286;
  wire g8287;
  wire g829;
  wire g8293;
  wire g8294;
  wire g8295;
  wire g8296;
  wire g83;
  wire g830;
  wire g8302;
  wire g8303;
  wire g8304;
  wire g8305;
  wire g831;
  wire g8311;
  wire g8312;
  wire g8313;
  wire g8317;
  wire g832;
  wire g8321;
  wire g8324;
  wire g833;
  wire g8330;
  wire g8333;
  wire g8336;
  wire g834;
  wire g8341;
  wire g8344;
  wire g8347;
  wire g835;
  wire g8351;
  wire g8354;
  wire g8357;
  wire g836;
  wire g8363;
  wire g8366;
  wire g8369;
  wire g837;
  wire g8372;
  wire g8375;
  wire g838;
  wire g8382;
  wire g8388;
  wire g839;
  wire g8391;
  wire g8397;
  wire g840;
  wire g8400;
  wire g8403;
  wire g8408;
  wire g841;
  wire g8411;
  wire g8414;
  wire g8418;
  wire g842;
  wire g8421;
  wire g8424;
  wire g843;
  wire g8434;
  wire g844;
  wire g8440;
  wire g8443;
  wire g8449;
  wire g845;
  wire g8452;
  wire g8455;
  wire g846;
  wire g8460;
  wire g8469;
  wire g847;
  wire g8475;
  wire g8478;
  wire g848;
  wire g849;
  wire g8494;
  wire g850;
  wire g851;
  wire g852;
  wire g853;
  wire g856;
  wire g8569;
  wire g857;
  wire g8575;
  wire g8578;
  wire g8579;
  wire g858;
  wire g8580;
  wire g8587;
  wire g859;
  wire g8594;
  wire g860;
  wire g8602;
  wire g8605;
  wire g861;
  wire g8614;
  wire g8617;
  wire g862;
  wire g8620;
  wire g8622;
  wire g8627;
  wire g863;
  wire g8630;
  wire g8632;
  wire g8637;
  wire g864;
  wire g8640;
  wire g8643;
  wire g8646;
  wire g8649;
  wire g865;
  wire g8651;
  wire g8655;
  wire g8658;
  wire g8659;
  wire g866;
  wire g8662;
  wire g8665;
  wire g8667;
  wire g867;
  wire g8670;
  wire g8673;
  wire g8677;
  wire g8678;
  wire g868;
  wire g8681;
  wire g8684;
  wire g8689;
  wire g869;
  wire g8690;
  wire g8693;
  wire g8696;
  wire g8699;
  wire g870;
  wire g8700;
  wire g8707;
  wire g8708;
  wire g8711;
  wire g8714;
  wire g8718;
  wire g8719;
  wire g873;
  wire g8745;
  wire g8748;
  wire g8752;
  wire g8756;
  wire g8757;
  wire g876;
  wire g8763;
  wire g8766;
  wire g8769;
  wire g8770;
  wire g8771;
  wire g8775;
  wire g8779;
  wire g8780;
  wire g8785;
  wire g8788;
  wire g879;
  wire g8791;
  wire g8792;
  wire g8793;
  wire g8794;
  wire g8798;
  wire g88;
  wire g8802;
  wire g8805;
  wire g8808;
  wire g8809;
  wire g8810;
  wire g8811;
  wire g8812;
  wire g8813;
  wire g8817;
  wire g882;
  wire g8820;
  wire g8821;
  wire g8822;
  wire g8823;
  wire g8824;
  wire g8825;
  wire g8826;
  wire g8827;
  wire g8828;
  wire g8829;
  wire g8832;
  wire g8835;
  wire g8836;
  wire g8839;
  wire g8840;
  wire g8843;
  wire g8844;
  wire g8845;
  wire g8846;
  wire g8847;
  wire g885;
  wire g8850;
  wire g8851;
  wire g8852;
  wire g8853;
  wire g8856;
  wire g8859;
  wire g8860;
  wire g8862;
  wire g8863;
  wire g8866;
  wire g8867;
  wire g8870;
  wire g8871;
  wire g8872;
  wire g8873;
  wire g8874;
  wire g8877;
  wire g8878;
  wire g8879;
  wire g888;
  wire g8882;
  wire g8885;
  wire g8888;
  wire g8891;
  wire g8893;
  wire g8894;
  wire g8897;
  wire g8898;
  wire g8900;
  wire g8901;
  wire g8904;
  wire g8905;
  wire g8908;
  wire g8909;
  wire g891;
  wire g8910;
  wire g8911;
  wire g8912;
  wire g8915;
  wire g8918;
  wire g8921;
  wire g8924;
  wire g8925;
  wire g8928;
  wire g8931;
  wire g8933;
  wire g8934;
  wire g8937;
  wire g8938;
  wire g894;
  wire g8940;
  wire g8941;
  wire g8944;
  wire g8945;
  wire g8948;
  wire g8949;
  wire g8952;
  wire g8955;
  wire g8958;
  wire g8961;
  wire g8964;
  wire g8965;
  wire g8968;
  wire g897;
  wire g8971;
  wire g8973;
  wire g8974;
  wire g8977;
  wire g8978;
  wire g8980;
  wire g8984;
  wire g8987;
  wire g8990;
  wire g8993;
  wire g8996;
  wire g8997;
  wire g900;
  wire g9000;
  wire g9003;
  wire g9005;
  wire g9006;
  wire g9010;
  wire g9013;
  wire g9016;
  wire g9019;
  wire g9022;
  wire g9025;
  wire g9027;
  wire g903;
  wire g9035;
  wire g9038;
  wire g9041;
  wire g9044;
  wire g9050;
  wire g9058;
  wire g906;
  wire g9067;
  wire g9084;
  wire g909;
  wire g912;
  wire g9128;
  wire g9134;
  wire g9140;
  wire g9146;
  wire g9149;
  wire g915;
  wire g9150;
  wire g9159;
  wire g9160;
  wire g9161;
  wire g9170;
  wire g9173;
  wire g9174;
  wire g918;
  wire g9183;
  wire g9184;
  wire g9187;
  wire g9196;
  wire g9199;
  wire g92;
  wire g9202;
  wire g9203;
  wire g921;
  wire g9212;
  wire g9215;
  wire g9216;
  wire g9225;
  wire g9226;
  wire g9227;
  wire g9228;
  wire g9229;
  wire g9232;
  wire g924;
  wire g9242;
  wire g9245;
  wire g9248;
  wire g9257;
  wire g9260;
  wire g9263;
  wire g9264;
  wire g927;
  wire g9273;
  wire g9276;
  wire g9277;
  wire g9286;
  wire g9287;
  wire g9288;
  wire g9289;
  wire g9290;
  wire g9293;
  wire g930;
  wire g9303;
  wire g9306;
  wire g9309;
  wire g9310;
  wire g9320;
  wire g9323;
  wire g9326;
  wire g933;
  wire g9335;
  wire g9338;
  wire g9341;
  wire g9342;
  wire g9351;
  wire g9354;
  wire g9355;
  wire g9356;
  wire g936;
  wire g9368;
  wire g9371;
  wire g9374;
  wire g9384;
  wire g9387;
  wire g939;
  wire g9390;
  wire g9391;
  wire g9401;
  wire g9404;
  wire g9407;
  wire g9416;
  wire g9419;
  wire g942;
  wire g9422;
  wire g9423;
  wire g9424;
  wire g9425;
  wire g9426;
  wire g9427;
  wire g9443;
  wire g9446;
  wire g9449;
  wire g945;
  wire g9450;
  wire g9453;
  wire g9465;
  wire g9468;
  wire g9471;
  wire g948;
  wire g9481;
  wire g9484;
  wire g9487;
  wire g9488;
  wire g9498;
  wire g9501;
  wire g9504;
  wire g9505;
  wire g9506;
  wire g9507;
  wire g951;
  wire g9524;
  wire g9528;
  wire g9531;
  wire g954;
  wire g9569;
  wire g957;
  wire g9585;
  wire g9588;
  wire g9591;
  wire g9592;
  wire g9595;
  wire g960;
  wire g9607;
  wire g9610;
  wire g9613;
  wire g9623;
  wire g9626;
  wire g9629;
  wire g963;
  wire g9640;
  wire g9641;
  wire g9644;
  wire g9649;
  wire g966;
  wire g9666;
  wire g967;
  wire g9670;
  wire g9673;
  wire g968;
  wire g969;
  wire g97;
  wire g970;
  wire g971;
  wire g9711;
  wire g972;
  wire g9727;
  wire g973;
  wire g9730;
  wire g9733;
  wire g9734;
  wire g9737;
  wire g974;
  wire g9749;
  wire g975;
  wire g9752;
  wire g9755;
  wire g9756;
  wire g9757;
  wire g9758;
  wire g976;
  wire g9767;
  wire g977;
  wire g9770;
  wire g978;
  wire g9786;
  wire g9787;
  wire g9790;
  wire g9795;
  wire g9812;
  wire g9816;
  wire g9819;
  wire g985;
  wire g9857;
  wire g986;
  wire g9873;
  wire g9876;
  wire g9879;
  wire g9880;
  wire g9884;
  wire g9885;
  wire g9886;
  wire g9895;
  wire g9898;
  wire g9913;
  wire g9916;
  wire g992;
  wire g9932;
  wire g9933;
  wire g9936;
  wire g9941;
  wire g9958;
  wire g996;
  wire g9962;
  wire g9965;
  wire g999;
  al_inv _3592_ (
    .a(\DFF_72.Q ),
    .y(\DFF_304.D )
  );
  al_inv _3593_ (
    .a(\DFF_74.Q ),
    .y(\DFF_306.D )
  );
  al_inv _3594_ (
    .a(\DFF_76.Q ),
    .y(\DFF_308.D )
  );
  al_inv _3595_ (
    .a(\DFF_78.Q ),
    .y(\DFF_310.D )
  );
  al_inv _3596_ (
    .a(\DFF_80.Q ),
    .y(\DFF_312.D )
  );
  al_inv _3597_ (
    .a(\DFF_66.Q ),
    .y(\DFF_298.D )
  );
  al_inv _3598_ (
    .a(\DFF_68.Q ),
    .y(\DFF_300.D )
  );
  al_inv _3599_ (
    .a(\DFF_70.Q ),
    .y(\DFF_302.D )
  );
  al_inv _3600_ (
    .a(\DFF_54.Q ),
    .y(\DFF_654.D )
  );
  al_inv _3601_ (
    .a(\DFF_56.Q ),
    .y(\DFF_656.D )
  );
  al_inv _3602_ (
    .a(\DFF_58.Q ),
    .y(\DFF_658.D )
  );
  al_inv _3603_ (
    .a(\DFF_60.Q ),
    .y(\DFF_660.D )
  );
  al_inv _3604_ (
    .a(\DFF_62.Q ),
    .y(\DFF_662.D )
  );
  al_inv _3605_ (
    .a(\DFF_48.Q ),
    .y(\DFF_648.D )
  );
  al_inv _3606_ (
    .a(\DFF_50.Q ),
    .y(\DFF_650.D )
  );
  al_inv _3607_ (
    .a(\DFF_52.Q ),
    .y(\DFF_652.D )
  );
  al_inv _3608_ (
    .a(\DFF_41.Q ),
    .y(\DFF_1004.D )
  );
  al_inv _3609_ (
    .a(\DFF_42.Q ),
    .y(\DFF_1006.D )
  );
  al_inv _3610_ (
    .a(\DFF_43.Q ),
    .y(\DFF_1008.D )
  );
  al_inv _3611_ (
    .a(\DFF_44.Q ),
    .y(\DFF_1010.D )
  );
  al_inv _3612_ (
    .a(\DFF_45.Q ),
    .y(\DFF_1012.D )
  );
  al_inv _3613_ (
    .a(\DFF_38.Q ),
    .y(\DFF_998.D )
  );
  al_inv _3614_ (
    .a(\DFF_39.Q ),
    .y(\DFF_1000.D )
  );
  al_inv _3615_ (
    .a(\DFF_40.Q ),
    .y(\DFF_1002.D )
  );
  al_inv _3616_ (
    .a(\DFF_86.Q ),
    .y(\DFF_1354.D )
  );
  al_inv _3617_ (
    .a(\DFF_87.Q ),
    .y(\DFF_1356.D )
  );
  al_inv _3618_ (
    .a(\DFF_88.Q ),
    .y(\DFF_1358.D )
  );
  al_inv _3619_ (
    .a(\DFF_89.Q ),
    .y(\DFF_1360.D )
  );
  al_inv _3620_ (
    .a(\DFF_90.Q ),
    .y(\DFF_1362.D )
  );
  al_inv _3621_ (
    .a(\DFF_83.Q ),
    .y(\DFF_1348.D )
  );
  al_inv _3622_ (
    .a(\DFF_84.Q ),
    .y(\DFF_1350.D )
  );
  al_inv _3623_ (
    .a(\DFF_85.Q ),
    .y(\DFF_1352.D )
  );
  al_inv _3624_ (
    .a(\DFF_299.Q ),
    .y(\DFF_444.D )
  );
  al_inv _3625_ (
    .a(\DFF_301.Q ),
    .y(\DFF_445.D )
  );
  al_inv _3626_ (
    .a(\DFF_303.Q ),
    .y(\DFF_446.D )
  );
  al_inv _3627_ (
    .a(\DFF_305.Q ),
    .y(\DFF_447.D )
  );
  al_inv _3628_ (
    .a(\DFF_307.Q ),
    .y(\DFF_448.D )
  );
  al_inv _3629_ (
    .a(\DFF_309.Q ),
    .y(\DFF_449.D )
  );
  al_inv _3630_ (
    .a(\DFF_311.Q ),
    .y(\DFF_450.D )
  );
  al_inv _3631_ (
    .a(\DFF_313.Q ),
    .y(\DFF_451.D )
  );
  al_inv _3632_ (
    .a(\DFF_315.Q ),
    .y(\DFF_453.D )
  );
  al_inv _3633_ (
    .a(\DFF_649.Q ),
    .y(\DFF_794.D )
  );
  al_inv _3634_ (
    .a(\DFF_651.Q ),
    .y(\DFF_795.D )
  );
  al_inv _3635_ (
    .a(\DFF_653.Q ),
    .y(\DFF_796.D )
  );
  al_inv _3636_ (
    .a(\DFF_655.Q ),
    .y(\DFF_797.D )
  );
  al_inv _3637_ (
    .a(\DFF_657.Q ),
    .y(\DFF_798.D )
  );
  al_inv _3638_ (
    .a(\DFF_659.Q ),
    .y(\DFF_799.D )
  );
  al_inv _3639_ (
    .a(\DFF_661.Q ),
    .y(\DFF_800.D )
  );
  al_inv _3640_ (
    .a(\DFF_663.Q ),
    .y(\DFF_801.D )
  );
  al_inv _3641_ (
    .a(\DFF_665.Q ),
    .y(\DFF_803.D )
  );
  al_inv _3642_ (
    .a(\DFF_999.Q ),
    .y(\DFF_1144.D )
  );
  al_inv _3643_ (
    .a(\DFF_1001.Q ),
    .y(\DFF_1145.D )
  );
  al_inv _3644_ (
    .a(\DFF_1003.Q ),
    .y(\DFF_1146.D )
  );
  al_inv _3645_ (
    .a(\DFF_1005.Q ),
    .y(\DFF_1147.D )
  );
  al_inv _3646_ (
    .a(\DFF_1007.Q ),
    .y(\DFF_1148.D )
  );
  al_inv _3647_ (
    .a(\DFF_1009.Q ),
    .y(\DFF_1149.D )
  );
  al_inv _3648_ (
    .a(\DFF_1011.Q ),
    .y(\DFF_1150.D )
  );
  al_inv _3649_ (
    .a(\DFF_1013.Q ),
    .y(\DFF_1151.D )
  );
  al_inv _3650_ (
    .a(\DFF_1015.Q ),
    .y(\DFF_1153.D )
  );
  al_inv _3651_ (
    .a(\DFF_1349.Q ),
    .y(\DFF_1494.D )
  );
  al_inv _3652_ (
    .a(\DFF_1351.Q ),
    .y(\DFF_1495.D )
  );
  al_inv _3653_ (
    .a(\DFF_1353.Q ),
    .y(\DFF_1496.D )
  );
  al_inv _3654_ (
    .a(\DFF_1355.Q ),
    .y(\DFF_1497.D )
  );
  al_inv _3655_ (
    .a(\DFF_1357.Q ),
    .y(\DFF_1498.D )
  );
  al_inv _3656_ (
    .a(\DFF_1359.Q ),
    .y(\DFF_1499.D )
  );
  al_inv _3657_ (
    .a(\DFF_1361.Q ),
    .y(\DFF_1500.D )
  );
  al_inv _3658_ (
    .a(\DFF_1363.Q ),
    .y(\DFF_1501.D )
  );
  al_inv _3659_ (
    .a(\DFF_1365.Q ),
    .y(\DFF_1503.D )
  );
  al_nand3ftt _3660_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_317.Q ),
    .c(\DFF_316.Q ),
    .y(_0000_)
  );
  al_oai21 _3661_ (
    .a(\DFF_316.Q ),
    .b(\DFF_328.Q ),
    .c(_0000_),
    .y(\DFF_317.D )
  );
  al_or3 _3662_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_432.Q ),
    .c(\DFF_442.Q ),
    .y(_0001_)
  );
  al_aoi21ftf _3663_ (
    .a(\DFF_433.Q ),
    .b(\DFF_432.Q ),
    .c(_0001_),
    .y(\DFF_442.D )
  );
  al_oai21ftf _3664_ (
    .a(\DFF_400.Q ),
    .b(\DFF_1504.Q ),
    .c(\DFF_402.Q ),
    .y(_0002_)
  );
  al_aoi21ftf _3665_ (
    .a(\DFF_399.Q ),
    .b(\DFF_402.Q ),
    .c(_0002_),
    .y(\DFF_400.D )
  );
  al_and2ft _3666_ (
    .a(\DFF_1605.Q ),
    .b(\DFF_1603.Q ),
    .y(_0003_)
  );
  al_nand3fft _3667_ (
    .a(\DFF_1600.Q ),
    .b(\DFF_1602.Q ),
    .c(\DFF_1604.Q ),
    .y(_0004_)
  );
  al_and2 _3668_ (
    .a(\DFF_1601.Q ),
    .b(\DFF_1606.Q ),
    .y(_0005_)
  );
  al_and3ftt _3669_ (
    .a(_0004_),
    .b(_0003_),
    .c(_0005_),
    .y(_0006_)
  );
  al_and3fft _3670_ (
    .a(\DFF_1609.Q ),
    .b(\DFF_1610.Q ),
    .c(\DFF_1607.Q ),
    .y(_0007_)
  );
  al_and3 _3671_ (
    .a(\DFF_1608.Q ),
    .b(_0007_),
    .c(_0006_),
    .y(_0008_)
  );
  al_inv _3672_ (
    .a(_0008_),
    .y(_0009_)
  );
  al_mux2h _3673_ (
    .a(\DFF_359.Q ),
    .b(_0009_),
    .s(\DFF_1506.Q ),
    .y(\DFF_359.D )
  );
  al_inv _3674_ (
    .a(\DFF_459.Q ),
    .y(_0010_)
  );
  al_and3ftt _3675_ (
    .a(\DFF_458.Q ),
    .b(\DFF_452.Q ),
    .c(\DFF_443.Q ),
    .y(_0011_)
  );
  al_nand2 _3676_ (
    .a(\DFF_1505.Q ),
    .b(_0011_),
    .y(_0012_)
  );
  al_mux2l _3677_ (
    .a(\DFF_470.Q ),
    .b(_0010_),
    .s(_0012_),
    .y(\DFF_470.D )
  );
  al_nand2 _3678_ (
    .a(\DFF_1506.Q ),
    .b(_0011_),
    .y(_0013_)
  );
  al_mux2l _3679_ (
    .a(\DFF_471.Q ),
    .b(_0010_),
    .s(_0013_),
    .y(\DFF_471.D )
  );
  al_inv _3680_ (
    .a(\DFF_460.Q ),
    .y(_0014_)
  );
  al_nand2 _3681_ (
    .a(\DFF_1504.Q ),
    .b(_0011_),
    .y(_0015_)
  );
  al_mux2l _3682_ (
    .a(\DFF_472.Q ),
    .b(_0014_),
    .s(_0015_),
    .y(\DFF_472.D )
  );
  al_mux2l _3683_ (
    .a(\DFF_473.Q ),
    .b(_0014_),
    .s(_0012_),
    .y(\DFF_473.D )
  );
  al_mux2l _3684_ (
    .a(\DFF_474.Q ),
    .b(_0014_),
    .s(_0013_),
    .y(\DFF_474.D )
  );
  al_inv _3685_ (
    .a(\DFF_461.Q ),
    .y(_0016_)
  );
  al_mux2l _3686_ (
    .a(\DFF_475.Q ),
    .b(_0016_),
    .s(_0015_),
    .y(\DFF_475.D )
  );
  al_mux2l _3687_ (
    .a(\DFF_476.Q ),
    .b(_0016_),
    .s(_0012_),
    .y(\DFF_476.D )
  );
  al_mux2l _3688_ (
    .a(\DFF_477.Q ),
    .b(_0016_),
    .s(_0013_),
    .y(\DFF_477.D )
  );
  al_inv _3689_ (
    .a(\DFF_462.Q ),
    .y(_0017_)
  );
  al_mux2l _3690_ (
    .a(\DFF_478.Q ),
    .b(_0017_),
    .s(_0015_),
    .y(\DFF_478.D )
  );
  al_mux2l _3691_ (
    .a(\DFF_479.Q ),
    .b(_0017_),
    .s(_0012_),
    .y(\DFF_479.D )
  );
  al_mux2l _3692_ (
    .a(\DFF_480.Q ),
    .b(_0017_),
    .s(_0013_),
    .y(\DFF_480.D )
  );
  al_inv _3693_ (
    .a(\DFF_463.Q ),
    .y(_0018_)
  );
  al_mux2l _3694_ (
    .a(\DFF_481.Q ),
    .b(_0018_),
    .s(_0015_),
    .y(\DFF_481.D )
  );
  al_mux2l _3695_ (
    .a(\DFF_482.Q ),
    .b(_0018_),
    .s(_0012_),
    .y(\DFF_482.D )
  );
  al_mux2l _3696_ (
    .a(\DFF_483.Q ),
    .b(_0018_),
    .s(_0013_),
    .y(\DFF_483.D )
  );
  al_inv _3697_ (
    .a(\DFF_464.Q ),
    .y(_0019_)
  );
  al_mux2l _3698_ (
    .a(\DFF_484.Q ),
    .b(_0019_),
    .s(_0015_),
    .y(\DFF_484.D )
  );
  al_mux2l _3699_ (
    .a(\DFF_485.Q ),
    .b(_0019_),
    .s(_0012_),
    .y(\DFF_485.D )
  );
  al_mux2l _3700_ (
    .a(\DFF_486.Q ),
    .b(_0019_),
    .s(_0013_),
    .y(\DFF_486.D )
  );
  al_inv _3701_ (
    .a(\DFF_465.Q ),
    .y(_0020_)
  );
  al_mux2l _3702_ (
    .a(\DFF_487.Q ),
    .b(_0020_),
    .s(_0015_),
    .y(\DFF_487.D )
  );
  al_mux2l _3703_ (
    .a(\DFF_488.Q ),
    .b(_0020_),
    .s(_0012_),
    .y(\DFF_488.D )
  );
  al_mux2l _3704_ (
    .a(\DFF_489.Q ),
    .b(_0020_),
    .s(_0013_),
    .y(\DFF_489.D )
  );
  al_inv _3705_ (
    .a(\DFF_466.Q ),
    .y(_0021_)
  );
  al_mux2l _3706_ (
    .a(\DFF_490.Q ),
    .b(_0021_),
    .s(_0015_),
    .y(\DFF_490.D )
  );
  al_mux2l _3707_ (
    .a(\DFF_491.Q ),
    .b(_0021_),
    .s(_0012_),
    .y(\DFF_491.D )
  );
  al_mux2l _3708_ (
    .a(\DFF_492.Q ),
    .b(_0021_),
    .s(_0013_),
    .y(\DFF_492.D )
  );
  al_inv _3709_ (
    .a(\DFF_467.Q ),
    .y(_0022_)
  );
  al_mux2l _3710_ (
    .a(\DFF_493.Q ),
    .b(_0022_),
    .s(_0015_),
    .y(\DFF_493.D )
  );
  al_mux2l _3711_ (
    .a(\DFF_494.Q ),
    .b(_0022_),
    .s(_0012_),
    .y(\DFF_494.D )
  );
  al_mux2l _3712_ (
    .a(\DFF_495.Q ),
    .b(_0022_),
    .s(_0013_),
    .y(\DFF_495.D )
  );
  al_inv _3713_ (
    .a(\DFF_468.Q ),
    .y(_0023_)
  );
  al_mux2l _3714_ (
    .a(\DFF_496.Q ),
    .b(_0023_),
    .s(_0015_),
    .y(\DFF_496.D )
  );
  al_mux2l _3715_ (
    .a(\DFF_497.Q ),
    .b(_0023_),
    .s(_0012_),
    .y(\DFF_497.D )
  );
  al_mux2l _3716_ (
    .a(\DFF_498.Q ),
    .b(_0023_),
    .s(_0013_),
    .y(\DFF_498.D )
  );
  al_and2 _3717_ (
    .a(\DFF_457.Q ),
    .b(\DFF_1504.Q ),
    .y(_0024_)
  );
  al_inv _3718_ (
    .a(\DFF_1504.Q ),
    .y(_0025_)
  );
  al_nand2 _3719_ (
    .a(\DFF_424.Q ),
    .b(\DFF_1505.Q ),
    .y(_0026_)
  );
  al_ao21ttf _3720_ (
    .a(\DFF_425.Q ),
    .b(\DFF_1506.Q ),
    .c(_0026_),
    .y(_0027_)
  );
  al_aoi21ftt _3721_ (
    .a(_0025_),
    .b(\DFF_423.Q ),
    .c(_0027_),
    .y(_0028_)
  );
  al_mux2h _3722_ (
    .a(\DFF_499.Q ),
    .b(_0028_),
    .s(_0024_),
    .y(\DFF_499.D )
  );
  al_and2 _3723_ (
    .a(\DFF_457.Q ),
    .b(\DFF_1505.Q ),
    .y(_0029_)
  );
  al_mux2h _3724_ (
    .a(\DFF_500.Q ),
    .b(_0028_),
    .s(_0029_),
    .y(\DFF_500.D )
  );
  al_and2 _3725_ (
    .a(\DFF_457.Q ),
    .b(\DFF_1506.Q ),
    .y(_0030_)
  );
  al_mux2h _3726_ (
    .a(\DFF_501.Q ),
    .b(_0028_),
    .s(_0030_),
    .y(\DFF_501.D )
  );
  al_nand2 _3727_ (
    .a(\DFF_427.Q ),
    .b(\DFF_1505.Q ),
    .y(_0031_)
  );
  al_aoi21ttf _3728_ (
    .a(\DFF_428.Q ),
    .b(\DFF_1506.Q ),
    .c(_0031_),
    .y(_0032_)
  );
  al_aoi21ftf _3729_ (
    .a(_0025_),
    .b(\DFF_426.Q ),
    .c(_0032_),
    .y(_0033_)
  );
  al_mux2h _3730_ (
    .a(\DFF_502.Q ),
    .b(_0033_),
    .s(_0024_),
    .y(\DFF_502.D )
  );
  al_mux2h _3731_ (
    .a(\DFF_503.Q ),
    .b(_0033_),
    .s(_0029_),
    .y(\DFF_503.D )
  );
  al_mux2h _3732_ (
    .a(\DFF_504.Q ),
    .b(_0033_),
    .s(_0030_),
    .y(\DFF_504.D )
  );
  al_mux2h _3733_ (
    .a(\DFF_709.Q ),
    .b(_0009_),
    .s(\DFF_1506.Q ),
    .y(\DFF_709.D )
  );
  al_and3ftt _3734_ (
    .a(\DFF_808.Q ),
    .b(\DFF_809.Q ),
    .c(\DFF_1506.Q ),
    .y(_0034_)
  );
  al_and2 _3735_ (
    .a(\DFF_807.Q ),
    .b(\DFF_1505.Q ),
    .y(_0035_)
  );
  al_oai21ftf _3736_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_808.Q ),
    .c(\DFF_809.Q ),
    .y(_0036_)
  );
  al_and3fft _3737_ (
    .a(_0034_),
    .b(_0035_),
    .c(_0036_),
    .y(\DFF_809.D )
  );
  al_inv _3738_ (
    .a(\DFF_809.Q ),
    .y(_0037_)
  );
  al_and3ftt _3739_ (
    .a(\DFF_808.Q ),
    .b(\DFF_802.Q ),
    .c(\DFF_793.Q ),
    .y(_0038_)
  );
  al_nand2 _3740_ (
    .a(\DFF_1504.Q ),
    .b(_0038_),
    .y(_0039_)
  );
  al_mux2l _3741_ (
    .a(\DFF_819.Q ),
    .b(_0037_),
    .s(_0039_),
    .y(\DFF_819.D )
  );
  al_nand2 _3742_ (
    .a(\DFF_1505.Q ),
    .b(_0038_),
    .y(_0040_)
  );
  al_mux2l _3743_ (
    .a(\DFF_820.Q ),
    .b(_0037_),
    .s(_0040_),
    .y(\DFF_820.D )
  );
  al_nand2 _3744_ (
    .a(\DFF_1506.Q ),
    .b(_0038_),
    .y(_0041_)
  );
  al_mux2l _3745_ (
    .a(\DFF_821.Q ),
    .b(_0037_),
    .s(_0041_),
    .y(\DFF_821.D )
  );
  al_inv _3746_ (
    .a(\DFF_810.Q ),
    .y(_0042_)
  );
  al_mux2l _3747_ (
    .a(\DFF_822.Q ),
    .b(_0042_),
    .s(_0039_),
    .y(\DFF_822.D )
  );
  al_mux2l _3748_ (
    .a(\DFF_823.Q ),
    .b(_0042_),
    .s(_0040_),
    .y(\DFF_823.D )
  );
  al_mux2l _3749_ (
    .a(\DFF_824.Q ),
    .b(_0042_),
    .s(_0041_),
    .y(\DFF_824.D )
  );
  al_inv _3750_ (
    .a(\DFF_811.Q ),
    .y(_0043_)
  );
  al_mux2l _3751_ (
    .a(\DFF_825.Q ),
    .b(_0043_),
    .s(_0039_),
    .y(\DFF_825.D )
  );
  al_mux2l _3752_ (
    .a(\DFF_826.Q ),
    .b(_0043_),
    .s(_0040_),
    .y(\DFF_826.D )
  );
  al_mux2l _3753_ (
    .a(\DFF_827.Q ),
    .b(_0043_),
    .s(_0041_),
    .y(\DFF_827.D )
  );
  al_inv _3754_ (
    .a(\DFF_812.Q ),
    .y(_0044_)
  );
  al_mux2l _3755_ (
    .a(\DFF_828.Q ),
    .b(_0044_),
    .s(_0039_),
    .y(\DFF_828.D )
  );
  al_mux2l _3756_ (
    .a(\DFF_829.Q ),
    .b(_0044_),
    .s(_0040_),
    .y(\DFF_829.D )
  );
  al_mux2l _3757_ (
    .a(\DFF_830.Q ),
    .b(_0044_),
    .s(_0041_),
    .y(\DFF_830.D )
  );
  al_inv _3758_ (
    .a(\DFF_813.Q ),
    .y(_0045_)
  );
  al_mux2l _3759_ (
    .a(\DFF_831.Q ),
    .b(_0045_),
    .s(_0039_),
    .y(\DFF_831.D )
  );
  al_mux2l _3760_ (
    .a(\DFF_832.Q ),
    .b(_0045_),
    .s(_0040_),
    .y(\DFF_832.D )
  );
  al_mux2l _3761_ (
    .a(\DFF_833.Q ),
    .b(_0045_),
    .s(_0041_),
    .y(\DFF_833.D )
  );
  al_inv _3762_ (
    .a(\DFF_814.Q ),
    .y(_0046_)
  );
  al_mux2l _3763_ (
    .a(\DFF_834.Q ),
    .b(_0046_),
    .s(_0039_),
    .y(\DFF_834.D )
  );
  al_mux2l _3764_ (
    .a(\DFF_835.Q ),
    .b(_0046_),
    .s(_0040_),
    .y(\DFF_835.D )
  );
  al_mux2l _3765_ (
    .a(\DFF_836.Q ),
    .b(_0046_),
    .s(_0041_),
    .y(\DFF_836.D )
  );
  al_inv _3766_ (
    .a(\DFF_815.Q ),
    .y(_0047_)
  );
  al_mux2l _3767_ (
    .a(\DFF_837.Q ),
    .b(_0047_),
    .s(_0039_),
    .y(\DFF_837.D )
  );
  al_mux2l _3768_ (
    .a(\DFF_838.Q ),
    .b(_0047_),
    .s(_0040_),
    .y(\DFF_838.D )
  );
  al_mux2l _3769_ (
    .a(\DFF_839.Q ),
    .b(_0047_),
    .s(_0041_),
    .y(\DFF_839.D )
  );
  al_inv _3770_ (
    .a(\DFF_816.Q ),
    .y(_0048_)
  );
  al_mux2l _3771_ (
    .a(\DFF_840.Q ),
    .b(_0048_),
    .s(_0039_),
    .y(\DFF_840.D )
  );
  al_mux2l _3772_ (
    .a(\DFF_841.Q ),
    .b(_0048_),
    .s(_0040_),
    .y(\DFF_841.D )
  );
  al_mux2l _3773_ (
    .a(\DFF_842.Q ),
    .b(_0048_),
    .s(_0041_),
    .y(\DFF_842.D )
  );
  al_inv _3774_ (
    .a(\DFF_817.Q ),
    .y(_0049_)
  );
  al_mux2l _3775_ (
    .a(\DFF_843.Q ),
    .b(_0049_),
    .s(_0039_),
    .y(\DFF_843.D )
  );
  al_mux2l _3776_ (
    .a(\DFF_844.Q ),
    .b(_0049_),
    .s(_0040_),
    .y(\DFF_844.D )
  );
  al_mux2l _3777_ (
    .a(\DFF_845.Q ),
    .b(_0049_),
    .s(_0041_),
    .y(\DFF_845.D )
  );
  al_inv _3778_ (
    .a(\DFF_818.Q ),
    .y(_0050_)
  );
  al_mux2l _3779_ (
    .a(\DFF_846.Q ),
    .b(_0050_),
    .s(_0039_),
    .y(\DFF_846.D )
  );
  al_mux2l _3780_ (
    .a(\DFF_847.Q ),
    .b(_0050_),
    .s(_0040_),
    .y(\DFF_847.D )
  );
  al_mux2l _3781_ (
    .a(\DFF_848.Q ),
    .b(_0050_),
    .s(_0041_),
    .y(\DFF_848.D )
  );
  al_and2 _3782_ (
    .a(\DFF_807.Q ),
    .b(\DFF_1504.Q ),
    .y(_0051_)
  );
  al_nand2 _3783_ (
    .a(\DFF_774.Q ),
    .b(\DFF_1505.Q ),
    .y(_0052_)
  );
  al_aoi21ttf _3784_ (
    .a(\DFF_775.Q ),
    .b(\DFF_1506.Q ),
    .c(_0052_),
    .y(_0053_)
  );
  al_ao21ftf _3785_ (
    .a(_0025_),
    .b(\DFF_773.Q ),
    .c(_0053_),
    .y(_0054_)
  );
  al_inv _3786_ (
    .a(_0054_),
    .y(_0055_)
  );
  al_mux2h _3787_ (
    .a(\DFF_849.Q ),
    .b(_0055_),
    .s(_0051_),
    .y(\DFF_849.D )
  );
  al_mux2h _3788_ (
    .a(\DFF_850.Q ),
    .b(_0055_),
    .s(_0035_),
    .y(\DFF_850.D )
  );
  al_and2 _3789_ (
    .a(\DFF_807.Q ),
    .b(\DFF_1506.Q ),
    .y(_0056_)
  );
  al_mux2h _3790_ (
    .a(\DFF_851.Q ),
    .b(_0055_),
    .s(_0056_),
    .y(\DFF_851.D )
  );
  al_nand2 _3791_ (
    .a(\DFF_777.Q ),
    .b(\DFF_1505.Q ),
    .y(_0057_)
  );
  al_aoi21ttf _3792_ (
    .a(\DFF_778.Q ),
    .b(\DFF_1506.Q ),
    .c(_0057_),
    .y(_0058_)
  );
  al_ao21ftf _3793_ (
    .a(_0025_),
    .b(\DFF_776.Q ),
    .c(_0058_),
    .y(_0059_)
  );
  al_inv _3794_ (
    .a(_0059_),
    .y(_0060_)
  );
  al_mux2h _3795_ (
    .a(\DFF_852.Q ),
    .b(_0060_),
    .s(_0051_),
    .y(\DFF_852.D )
  );
  al_mux2h _3796_ (
    .a(\DFF_853.Q ),
    .b(_0060_),
    .s(_0035_),
    .y(\DFF_853.D )
  );
  al_mux2h _3797_ (
    .a(\DFF_854.Q ),
    .b(_0060_),
    .s(_0056_),
    .y(\DFF_854.D )
  );
  al_mux2h _3798_ (
    .a(\DFF_1059.Q ),
    .b(_0009_),
    .s(\DFF_1506.Q ),
    .y(\DFF_1059.D )
  );
  al_and3ftt _3799_ (
    .a(\DFF_1158.Q ),
    .b(\DFF_1159.Q ),
    .c(\DFF_1506.Q ),
    .y(_0061_)
  );
  al_and2 _3800_ (
    .a(\DFF_1157.Q ),
    .b(\DFF_1505.Q ),
    .y(_0062_)
  );
  al_oai21ftf _3801_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_1158.Q ),
    .c(\DFF_1159.Q ),
    .y(_0063_)
  );
  al_and3fft _3802_ (
    .a(_0061_),
    .b(_0062_),
    .c(_0063_),
    .y(\DFF_1159.D )
  );
  al_inv _3803_ (
    .a(\DFF_1159.Q ),
    .y(_0064_)
  );
  al_and3ftt _3804_ (
    .a(\DFF_1158.Q ),
    .b(\DFF_1152.Q ),
    .c(\DFF_1143.Q ),
    .y(_0065_)
  );
  al_nand2 _3805_ (
    .a(\DFF_1504.Q ),
    .b(_0065_),
    .y(_0066_)
  );
  al_mux2l _3806_ (
    .a(\DFF_1169.Q ),
    .b(_0064_),
    .s(_0066_),
    .y(\DFF_1169.D )
  );
  al_nand2 _3807_ (
    .a(\DFF_1505.Q ),
    .b(_0065_),
    .y(_0067_)
  );
  al_mux2l _3808_ (
    .a(\DFF_1170.Q ),
    .b(_0064_),
    .s(_0067_),
    .y(\DFF_1170.D )
  );
  al_nand2 _3809_ (
    .a(\DFF_1506.Q ),
    .b(_0065_),
    .y(_0068_)
  );
  al_mux2l _3810_ (
    .a(\DFF_1171.Q ),
    .b(_0064_),
    .s(_0068_),
    .y(\DFF_1171.D )
  );
  al_inv _3811_ (
    .a(\DFF_1160.Q ),
    .y(_0069_)
  );
  al_mux2l _3812_ (
    .a(\DFF_1172.Q ),
    .b(_0069_),
    .s(_0066_),
    .y(\DFF_1172.D )
  );
  al_mux2l _3813_ (
    .a(\DFF_1173.Q ),
    .b(_0069_),
    .s(_0067_),
    .y(\DFF_1173.D )
  );
  al_mux2l _3814_ (
    .a(\DFF_1174.Q ),
    .b(_0069_),
    .s(_0068_),
    .y(\DFF_1174.D )
  );
  al_inv _3815_ (
    .a(\DFF_1161.Q ),
    .y(_0070_)
  );
  al_mux2l _3816_ (
    .a(\DFF_1175.Q ),
    .b(_0070_),
    .s(_0066_),
    .y(\DFF_1175.D )
  );
  al_mux2l _3817_ (
    .a(\DFF_1176.Q ),
    .b(_0070_),
    .s(_0067_),
    .y(\DFF_1176.D )
  );
  al_mux2l _3818_ (
    .a(\DFF_1177.Q ),
    .b(_0070_),
    .s(_0068_),
    .y(\DFF_1177.D )
  );
  al_inv _3819_ (
    .a(\DFF_1162.Q ),
    .y(_0071_)
  );
  al_mux2l _3820_ (
    .a(\DFF_1178.Q ),
    .b(_0071_),
    .s(_0066_),
    .y(\DFF_1178.D )
  );
  al_mux2l _3821_ (
    .a(\DFF_1179.Q ),
    .b(_0071_),
    .s(_0067_),
    .y(\DFF_1179.D )
  );
  al_mux2l _3822_ (
    .a(\DFF_1180.Q ),
    .b(_0071_),
    .s(_0068_),
    .y(\DFF_1180.D )
  );
  al_inv _3823_ (
    .a(\DFF_1163.Q ),
    .y(_0072_)
  );
  al_mux2l _3824_ (
    .a(\DFF_1181.Q ),
    .b(_0072_),
    .s(_0066_),
    .y(\DFF_1181.D )
  );
  al_mux2l _3825_ (
    .a(\DFF_1182.Q ),
    .b(_0072_),
    .s(_0067_),
    .y(\DFF_1182.D )
  );
  al_mux2l _3826_ (
    .a(\DFF_1183.Q ),
    .b(_0072_),
    .s(_0068_),
    .y(\DFF_1183.D )
  );
  al_inv _3827_ (
    .a(\DFF_1164.Q ),
    .y(_0073_)
  );
  al_mux2l _3828_ (
    .a(\DFF_1184.Q ),
    .b(_0073_),
    .s(_0066_),
    .y(\DFF_1184.D )
  );
  al_mux2l _3829_ (
    .a(\DFF_1185.Q ),
    .b(_0073_),
    .s(_0067_),
    .y(\DFF_1185.D )
  );
  al_mux2l _3830_ (
    .a(\DFF_1186.Q ),
    .b(_0073_),
    .s(_0068_),
    .y(\DFF_1186.D )
  );
  al_inv _3831_ (
    .a(\DFF_1165.Q ),
    .y(_0074_)
  );
  al_mux2l _3832_ (
    .a(\DFF_1187.Q ),
    .b(_0074_),
    .s(_0066_),
    .y(\DFF_1187.D )
  );
  al_mux2l _3833_ (
    .a(\DFF_1188.Q ),
    .b(_0074_),
    .s(_0067_),
    .y(\DFF_1188.D )
  );
  al_mux2l _3834_ (
    .a(\DFF_1189.Q ),
    .b(_0074_),
    .s(_0068_),
    .y(\DFF_1189.D )
  );
  al_inv _3835_ (
    .a(\DFF_1166.Q ),
    .y(_0075_)
  );
  al_mux2l _3836_ (
    .a(\DFF_1190.Q ),
    .b(_0075_),
    .s(_0066_),
    .y(\DFF_1190.D )
  );
  al_mux2l _3837_ (
    .a(\DFF_1191.Q ),
    .b(_0075_),
    .s(_0067_),
    .y(\DFF_1191.D )
  );
  al_mux2l _3838_ (
    .a(\DFF_1192.Q ),
    .b(_0075_),
    .s(_0068_),
    .y(\DFF_1192.D )
  );
  al_inv _3839_ (
    .a(\DFF_1167.Q ),
    .y(_0076_)
  );
  al_mux2l _3840_ (
    .a(\DFF_1193.Q ),
    .b(_0076_),
    .s(_0066_),
    .y(\DFF_1193.D )
  );
  al_mux2l _3841_ (
    .a(\DFF_1194.Q ),
    .b(_0076_),
    .s(_0067_),
    .y(\DFF_1194.D )
  );
  al_mux2l _3842_ (
    .a(\DFF_1195.Q ),
    .b(_0076_),
    .s(_0068_),
    .y(\DFF_1195.D )
  );
  al_inv _3843_ (
    .a(\DFF_1168.Q ),
    .y(_0077_)
  );
  al_mux2l _3844_ (
    .a(\DFF_1196.Q ),
    .b(_0077_),
    .s(_0066_),
    .y(\DFF_1196.D )
  );
  al_mux2l _3845_ (
    .a(\DFF_1197.Q ),
    .b(_0077_),
    .s(_0067_),
    .y(\DFF_1197.D )
  );
  al_mux2l _3846_ (
    .a(\DFF_1198.Q ),
    .b(_0077_),
    .s(_0068_),
    .y(\DFF_1198.D )
  );
  al_and2 _3847_ (
    .a(\DFF_1157.Q ),
    .b(\DFF_1504.Q ),
    .y(_0078_)
  );
  al_nand2 _3848_ (
    .a(\DFF_1124.Q ),
    .b(\DFF_1505.Q ),
    .y(_0079_)
  );
  al_aoi21ttf _3849_ (
    .a(\DFF_1125.Q ),
    .b(\DFF_1506.Q ),
    .c(_0079_),
    .y(_0080_)
  );
  al_ao21ftf _3850_ (
    .a(_0025_),
    .b(\DFF_1123.Q ),
    .c(_0080_),
    .y(_0081_)
  );
  al_inv _3851_ (
    .a(_0081_),
    .y(_0082_)
  );
  al_mux2h _3852_ (
    .a(\DFF_1199.Q ),
    .b(_0082_),
    .s(_0078_),
    .y(\DFF_1199.D )
  );
  al_mux2h _3853_ (
    .a(\DFF_1200.Q ),
    .b(_0082_),
    .s(_0062_),
    .y(\DFF_1200.D )
  );
  al_and2 _3854_ (
    .a(\DFF_1157.Q ),
    .b(\DFF_1506.Q ),
    .y(_0083_)
  );
  al_mux2h _3855_ (
    .a(\DFF_1201.Q ),
    .b(_0082_),
    .s(_0083_),
    .y(\DFF_1201.D )
  );
  al_nand2 _3856_ (
    .a(\DFF_1127.Q ),
    .b(\DFF_1505.Q ),
    .y(_0084_)
  );
  al_aoi21ttf _3857_ (
    .a(\DFF_1128.Q ),
    .b(\DFF_1506.Q ),
    .c(_0084_),
    .y(_0085_)
  );
  al_aoi21ftf _3858_ (
    .a(_0025_),
    .b(\DFF_1126.Q ),
    .c(_0085_),
    .y(_0086_)
  );
  al_mux2h _3859_ (
    .a(\DFF_1202.Q ),
    .b(_0086_),
    .s(_0078_),
    .y(\DFF_1202.D )
  );
  al_mux2h _3860_ (
    .a(\DFF_1203.Q ),
    .b(_0086_),
    .s(_0062_),
    .y(\DFF_1203.D )
  );
  al_mux2h _3861_ (
    .a(\DFF_1204.Q ),
    .b(_0086_),
    .s(_0083_),
    .y(\DFF_1204.D )
  );
  al_mux2h _3862_ (
    .a(\DFF_1409.Q ),
    .b(_0009_),
    .s(\DFF_1506.Q ),
    .y(\DFF_1409.D )
  );
  al_and3ftt _3863_ (
    .a(\DFF_1508.Q ),
    .b(\DFF_1509.Q ),
    .c(\DFF_1506.Q ),
    .y(_0087_)
  );
  al_and2 _3864_ (
    .a(\DFF_1507.Q ),
    .b(\DFF_1505.Q ),
    .y(_0088_)
  );
  al_oai21ftf _3865_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_1508.Q ),
    .c(\DFF_1509.Q ),
    .y(_0089_)
  );
  al_and3fft _3866_ (
    .a(_0087_),
    .b(_0088_),
    .c(_0089_),
    .y(\DFF_1509.D )
  );
  al_inv _3867_ (
    .a(\DFF_1509.Q ),
    .y(_0090_)
  );
  al_and3ftt _3868_ (
    .a(\DFF_1508.Q ),
    .b(\DFF_1502.Q ),
    .c(\DFF_1493.Q ),
    .y(_0091_)
  );
  al_nand2 _3869_ (
    .a(\DFF_1504.Q ),
    .b(_0091_),
    .y(_0092_)
  );
  al_mux2l _3870_ (
    .a(\DFF_1519.Q ),
    .b(_0090_),
    .s(_0092_),
    .y(\DFF_1519.D )
  );
  al_nand2 _3871_ (
    .a(\DFF_1505.Q ),
    .b(_0091_),
    .y(_0093_)
  );
  al_mux2l _3872_ (
    .a(\DFF_1520.Q ),
    .b(_0090_),
    .s(_0093_),
    .y(\DFF_1520.D )
  );
  al_nand2 _3873_ (
    .a(\DFF_1506.Q ),
    .b(_0091_),
    .y(_0094_)
  );
  al_mux2l _3874_ (
    .a(\DFF_1521.Q ),
    .b(_0090_),
    .s(_0094_),
    .y(\DFF_1521.D )
  );
  al_inv _3875_ (
    .a(\DFF_1510.Q ),
    .y(_0095_)
  );
  al_mux2l _3876_ (
    .a(\DFF_1522.Q ),
    .b(_0095_),
    .s(_0092_),
    .y(\DFF_1522.D )
  );
  al_mux2l _3877_ (
    .a(\DFF_1523.Q ),
    .b(_0095_),
    .s(_0093_),
    .y(\DFF_1523.D )
  );
  al_mux2l _3878_ (
    .a(\DFF_1524.Q ),
    .b(_0095_),
    .s(_0094_),
    .y(\DFF_1524.D )
  );
  al_inv _3879_ (
    .a(\DFF_1511.Q ),
    .y(_0096_)
  );
  al_mux2l _3880_ (
    .a(\DFF_1525.Q ),
    .b(_0096_),
    .s(_0092_),
    .y(\DFF_1525.D )
  );
  al_mux2l _3881_ (
    .a(\DFF_1526.Q ),
    .b(_0096_),
    .s(_0093_),
    .y(\DFF_1526.D )
  );
  al_mux2l _3882_ (
    .a(\DFF_1527.Q ),
    .b(_0096_),
    .s(_0094_),
    .y(\DFF_1527.D )
  );
  al_inv _3883_ (
    .a(\DFF_1512.Q ),
    .y(_0097_)
  );
  al_mux2l _3884_ (
    .a(\DFF_1528.Q ),
    .b(_0097_),
    .s(_0092_),
    .y(\DFF_1528.D )
  );
  al_mux2l _3885_ (
    .a(\DFF_1529.Q ),
    .b(_0097_),
    .s(_0093_),
    .y(\DFF_1529.D )
  );
  al_mux2l _3886_ (
    .a(\DFF_1530.Q ),
    .b(_0097_),
    .s(_0094_),
    .y(\DFF_1530.D )
  );
  al_inv _3887_ (
    .a(\DFF_1513.Q ),
    .y(_0098_)
  );
  al_mux2l _3888_ (
    .a(\DFF_1531.Q ),
    .b(_0098_),
    .s(_0092_),
    .y(\DFF_1531.D )
  );
  al_mux2l _3889_ (
    .a(\DFF_1532.Q ),
    .b(_0098_),
    .s(_0093_),
    .y(\DFF_1532.D )
  );
  al_mux2l _3890_ (
    .a(\DFF_1533.Q ),
    .b(_0098_),
    .s(_0094_),
    .y(\DFF_1533.D )
  );
  al_inv _3891_ (
    .a(\DFF_1514.Q ),
    .y(_0099_)
  );
  al_mux2l _3892_ (
    .a(\DFF_1534.Q ),
    .b(_0099_),
    .s(_0092_),
    .y(\DFF_1534.D )
  );
  al_mux2l _3893_ (
    .a(\DFF_1535.Q ),
    .b(_0099_),
    .s(_0093_),
    .y(\DFF_1535.D )
  );
  al_mux2l _3894_ (
    .a(\DFF_1536.Q ),
    .b(_0099_),
    .s(_0094_),
    .y(\DFF_1536.D )
  );
  al_inv _3895_ (
    .a(\DFF_1515.Q ),
    .y(_0100_)
  );
  al_mux2l _3896_ (
    .a(\DFF_1537.Q ),
    .b(_0100_),
    .s(_0092_),
    .y(\DFF_1537.D )
  );
  al_mux2l _3897_ (
    .a(\DFF_1538.Q ),
    .b(_0100_),
    .s(_0093_),
    .y(\DFF_1538.D )
  );
  al_mux2l _3898_ (
    .a(\DFF_1539.Q ),
    .b(_0100_),
    .s(_0094_),
    .y(\DFF_1539.D )
  );
  al_inv _3899_ (
    .a(\DFF_1516.Q ),
    .y(_0101_)
  );
  al_mux2l _3900_ (
    .a(\DFF_1540.Q ),
    .b(_0101_),
    .s(_0092_),
    .y(\DFF_1540.D )
  );
  al_mux2l _3901_ (
    .a(\DFF_1541.Q ),
    .b(_0101_),
    .s(_0093_),
    .y(\DFF_1541.D )
  );
  al_mux2l _3902_ (
    .a(\DFF_1542.Q ),
    .b(_0101_),
    .s(_0094_),
    .y(\DFF_1542.D )
  );
  al_inv _3903_ (
    .a(\DFF_1517.Q ),
    .y(_0102_)
  );
  al_mux2l _3904_ (
    .a(\DFF_1543.Q ),
    .b(_0102_),
    .s(_0092_),
    .y(\DFF_1543.D )
  );
  al_mux2l _3905_ (
    .a(\DFF_1544.Q ),
    .b(_0102_),
    .s(_0093_),
    .y(\DFF_1544.D )
  );
  al_mux2l _3906_ (
    .a(\DFF_1545.Q ),
    .b(_0102_),
    .s(_0094_),
    .y(\DFF_1545.D )
  );
  al_inv _3907_ (
    .a(\DFF_1518.Q ),
    .y(_0103_)
  );
  al_mux2l _3908_ (
    .a(\DFF_1546.Q ),
    .b(_0103_),
    .s(_0092_),
    .y(\DFF_1546.D )
  );
  al_mux2l _3909_ (
    .a(\DFF_1547.Q ),
    .b(_0103_),
    .s(_0093_),
    .y(\DFF_1547.D )
  );
  al_mux2l _3910_ (
    .a(\DFF_1548.Q ),
    .b(_0103_),
    .s(_0094_),
    .y(\DFF_1548.D )
  );
  al_and2 _3911_ (
    .a(\DFF_1507.Q ),
    .b(\DFF_1504.Q ),
    .y(_0104_)
  );
  al_nand2 _3912_ (
    .a(\DFF_1474.Q ),
    .b(\DFF_1505.Q ),
    .y(_0105_)
  );
  al_aoi21ttf _3913_ (
    .a(\DFF_1475.Q ),
    .b(\DFF_1506.Q ),
    .c(_0105_),
    .y(_0106_)
  );
  al_aoi21ftf _3914_ (
    .a(_0025_),
    .b(\DFF_1473.Q ),
    .c(_0106_),
    .y(_0107_)
  );
  al_mux2h _3915_ (
    .a(\DFF_1549.Q ),
    .b(_0107_),
    .s(_0104_),
    .y(\DFF_1549.D )
  );
  al_mux2h _3916_ (
    .a(\DFF_1550.Q ),
    .b(_0107_),
    .s(_0088_),
    .y(\DFF_1550.D )
  );
  al_and2 _3917_ (
    .a(\DFF_1507.Q ),
    .b(\DFF_1506.Q ),
    .y(_0108_)
  );
  al_mux2h _3918_ (
    .a(\DFF_1551.Q ),
    .b(_0107_),
    .s(_0108_),
    .y(\DFF_1551.D )
  );
  al_nand2 _3919_ (
    .a(\DFF_1477.Q ),
    .b(\DFF_1505.Q ),
    .y(_0109_)
  );
  al_aoi21ttf _3920_ (
    .a(\DFF_1478.Q ),
    .b(\DFF_1506.Q ),
    .c(_0109_),
    .y(_0110_)
  );
  al_aoi21ftf _3921_ (
    .a(_0025_),
    .b(\DFF_1476.Q ),
    .c(_0110_),
    .y(_0111_)
  );
  al_mux2h _3922_ (
    .a(\DFF_1552.Q ),
    .b(_0111_),
    .s(_0104_),
    .y(\DFF_1552.D )
  );
  al_mux2h _3923_ (
    .a(\DFF_1553.Q ),
    .b(_0111_),
    .s(_0088_),
    .y(\DFF_1553.D )
  );
  al_mux2h _3924_ (
    .a(\DFF_1554.Q ),
    .b(_0111_),
    .s(_0108_),
    .y(\DFF_1554.D )
  );
  al_inv _3925_ (
    .a(\DFF_19.Q ),
    .y(_0112_)
  );
  al_inv _3926_ (
    .a(g3231),
    .y(_0113_)
  );
  al_and2ft _3927_ (
    .a(\DFF_32.Q ),
    .b(\DFF_33.Q ),
    .y(_0114_)
  );
  al_nand2ft _3928_ (
    .a(\DFF_33.Q ),
    .b(\DFF_32.Q ),
    .y(_0115_)
  );
  al_and2ft _3929_ (
    .a(\DFF_31.Q ),
    .b(\DFF_30.Q ),
    .y(_0116_)
  );
  al_nand2ft _3930_ (
    .a(\DFF_30.Q ),
    .b(\DFF_31.Q ),
    .y(_0117_)
  );
  al_nand2ft _3931_ (
    .a(_0116_),
    .b(_0117_),
    .y(_0118_)
  );
  al_aoi21ftf _3932_ (
    .a(_0114_),
    .b(_0115_),
    .c(_0118_),
    .y(_0119_)
  );
  al_and3fft _3933_ (
    .a(_0114_),
    .b(_0118_),
    .c(_0115_),
    .y(_0120_)
  );
  al_and2ft _3934_ (
    .a(\DFF_34.Q ),
    .b(\DFF_35.Q ),
    .y(_0121_)
  );
  al_nand2ft _3935_ (
    .a(\DFF_35.Q ),
    .b(\DFF_34.Q ),
    .y(_0122_)
  );
  al_nand2 _3936_ (
    .a(\DFF_36.Q ),
    .b(\DFF_37.Q ),
    .y(_0123_)
  );
  al_nor2 _3937_ (
    .a(\DFF_36.Q ),
    .b(\DFF_37.Q ),
    .y(_0124_)
  );
  al_nand2ft _3938_ (
    .a(_0124_),
    .b(_0123_),
    .y(_0125_)
  );
  al_or3ftt _3939_ (
    .a(_0122_),
    .b(_0121_),
    .c(_0125_),
    .y(_0126_)
  );
  al_aoi21ftf _3940_ (
    .a(_0121_),
    .b(_0122_),
    .c(_0125_),
    .y(_0127_)
  );
  al_nand2ft _3941_ (
    .a(_0127_),
    .b(_0126_),
    .y(_0128_)
  );
  al_nand3fft _3942_ (
    .a(_0119_),
    .b(_0120_),
    .c(_0128_),
    .y(_0129_)
  );
  al_oai21ttf _3943_ (
    .a(_0119_),
    .b(_0120_),
    .c(_0128_),
    .y(_0130_)
  );
  al_and2 _3944_ (
    .a(_0129_),
    .b(_0130_),
    .y(_0131_)
  );
  al_and3 _3945_ (
    .a(\DFF_157.Q ),
    .b(_0113_),
    .c(_0131_),
    .y(_0132_)
  );
  al_ao21ftt _3946_ (
    .a(g3231),
    .b(\DFF_157.Q ),
    .c(_0131_),
    .y(_0133_)
  );
  al_nand2ft _3947_ (
    .a(_0132_),
    .b(_0133_),
    .y(_0134_)
  );
  al_mux2h _3948_ (
    .a(\DFF_63.Q ),
    .b(_0134_),
    .s(_0112_),
    .y(\DFF_63.D )
  );
  al_and2ft _3949_ (
    .a(\DFF_23.Q ),
    .b(\DFF_24.Q ),
    .y(_0135_)
  );
  al_nand2ft _3950_ (
    .a(\DFF_24.Q ),
    .b(\DFF_23.Q ),
    .y(_0136_)
  );
  al_and2ft _3951_ (
    .a(\DFF_22.Q ),
    .b(\DFF_21.Q ),
    .y(_0137_)
  );
  al_nand2ft _3952_ (
    .a(\DFF_21.Q ),
    .b(\DFF_22.Q ),
    .y(_0138_)
  );
  al_nand2ft _3953_ (
    .a(_0137_),
    .b(_0138_),
    .y(_0139_)
  );
  al_aoi21ftf _3954_ (
    .a(_0135_),
    .b(_0136_),
    .c(_0139_),
    .y(_0140_)
  );
  al_and3fft _3955_ (
    .a(_0135_),
    .b(_0139_),
    .c(_0136_),
    .y(_0141_)
  );
  al_and2ft _3956_ (
    .a(\DFF_28.Q ),
    .b(\DFF_25.Q ),
    .y(_0142_)
  );
  al_nand2ft _3957_ (
    .a(\DFF_25.Q ),
    .b(\DFF_28.Q ),
    .y(_0143_)
  );
  al_nand2 _3958_ (
    .a(\DFF_26.Q ),
    .b(\DFF_27.Q ),
    .y(_0144_)
  );
  al_nor2 _3959_ (
    .a(\DFF_26.Q ),
    .b(\DFF_27.Q ),
    .y(_0145_)
  );
  al_nand2ft _3960_ (
    .a(_0145_),
    .b(_0144_),
    .y(_0146_)
  );
  al_or3ftt _3961_ (
    .a(_0143_),
    .b(_0142_),
    .c(_0146_),
    .y(_0147_)
  );
  al_aoi21ftf _3962_ (
    .a(_0142_),
    .b(_0143_),
    .c(_0146_),
    .y(_0148_)
  );
  al_nand2ft _3963_ (
    .a(_0148_),
    .b(_0147_),
    .y(_0149_)
  );
  al_nand3fft _3964_ (
    .a(_0140_),
    .b(_0141_),
    .c(_0149_),
    .y(_0150_)
  );
  al_oai21ttf _3965_ (
    .a(_0140_),
    .b(_0141_),
    .c(_0149_),
    .y(_0151_)
  );
  al_and2 _3966_ (
    .a(_0150_),
    .b(_0151_),
    .y(_0152_)
  );
  al_and3 _3967_ (
    .a(\DFF_157.Q ),
    .b(_0113_),
    .c(_0152_),
    .y(_0153_)
  );
  al_ao21ftt _3968_ (
    .a(g3231),
    .b(\DFF_157.Q ),
    .c(_0152_),
    .y(_0154_)
  );
  al_nand2ft _3969_ (
    .a(_0153_),
    .b(_0154_),
    .y(_0155_)
  );
  al_mux2h _3970_ (
    .a(\DFF_46.Q ),
    .b(_0155_),
    .s(\DFF_19.Q ),
    .y(\DFF_46.D )
  );
  al_mux2h _3971_ (
    .a(\DFF_91.Q ),
    .b(_0134_),
    .s(\DFF_19.Q ),
    .y(\DFF_91.D )
  );
  al_mux2h _3972_ (
    .a(\DFF_81.Q ),
    .b(_0155_),
    .s(_0112_),
    .y(\DFF_81.D )
  );
  al_and2ft _3973_ (
    .a(g3234),
    .b(\DFF_1563.Q ),
    .y(\DFF_1561.D )
  );
  al_and2ft _3974_ (
    .a(g3234),
    .b(\DFF_1561.Q ),
    .y(\DFF_1562.D )
  );
  al_and2 _3975_ (
    .a(\DFF_1302.Q ),
    .b(\DFF_1427.Q ),
    .y(_0156_)
  );
  al_mux2l _3976_ (
    .a(\DFF_312.D ),
    .b(\DFF_164.Q ),
    .s(_0156_),
    .y(\DFF_164.D )
  );
  al_and2 _3977_ (
    .a(\DFF_1302.Q ),
    .b(\DFF_1428.Q ),
    .y(_0157_)
  );
  al_mux2l _3978_ (
    .a(\DFF_312.D ),
    .b(\DFF_165.Q ),
    .s(_0157_),
    .y(\DFF_165.D )
  );
  al_and2 _3979_ (
    .a(\DFF_1302.Q ),
    .b(\DFF_1429.Q ),
    .y(_0158_)
  );
  al_mux2l _3980_ (
    .a(\DFF_312.D ),
    .b(\DFF_166.Q ),
    .s(_0158_),
    .y(\DFF_166.D )
  );
  al_mux2l _3981_ (
    .a(\DFF_310.D ),
    .b(\DFF_167.Q ),
    .s(_0156_),
    .y(\DFF_167.D )
  );
  al_mux2l _3982_ (
    .a(\DFF_310.D ),
    .b(\DFF_168.Q ),
    .s(_0157_),
    .y(\DFF_168.D )
  );
  al_mux2l _3983_ (
    .a(\DFF_310.D ),
    .b(\DFF_169.Q ),
    .s(_0158_),
    .y(\DFF_169.D )
  );
  al_mux2l _3984_ (
    .a(\DFF_308.D ),
    .b(\DFF_170.Q ),
    .s(_0156_),
    .y(\DFF_170.D )
  );
  al_mux2l _3985_ (
    .a(\DFF_308.D ),
    .b(\DFF_171.Q ),
    .s(_0157_),
    .y(\DFF_171.D )
  );
  al_mux2l _3986_ (
    .a(\DFF_308.D ),
    .b(\DFF_172.Q ),
    .s(_0158_),
    .y(\DFF_172.D )
  );
  al_mux2l _3987_ (
    .a(\DFF_306.D ),
    .b(\DFF_173.Q ),
    .s(_0156_),
    .y(\DFF_173.D )
  );
  al_mux2l _3988_ (
    .a(\DFF_306.D ),
    .b(\DFF_174.Q ),
    .s(_0157_),
    .y(\DFF_174.D )
  );
  al_mux2l _3989_ (
    .a(\DFF_306.D ),
    .b(\DFF_175.Q ),
    .s(_0158_),
    .y(\DFF_175.D )
  );
  al_mux2l _3990_ (
    .a(\DFF_304.D ),
    .b(\DFF_176.Q ),
    .s(_0156_),
    .y(\DFF_176.D )
  );
  al_mux2l _3991_ (
    .a(\DFF_304.D ),
    .b(\DFF_177.Q ),
    .s(_0157_),
    .y(\DFF_177.D )
  );
  al_mux2l _3992_ (
    .a(\DFF_304.D ),
    .b(\DFF_178.Q ),
    .s(_0158_),
    .y(\DFF_178.D )
  );
  al_mux2l _3993_ (
    .a(\DFF_302.D ),
    .b(\DFF_179.Q ),
    .s(_0156_),
    .y(\DFF_179.D )
  );
  al_mux2l _3994_ (
    .a(\DFF_302.D ),
    .b(\DFF_180.Q ),
    .s(_0157_),
    .y(\DFF_180.D )
  );
  al_mux2l _3995_ (
    .a(\DFF_302.D ),
    .b(\DFF_181.Q ),
    .s(_0158_),
    .y(\DFF_181.D )
  );
  al_mux2l _3996_ (
    .a(\DFF_300.D ),
    .b(\DFF_182.Q ),
    .s(_0156_),
    .y(\DFF_182.D )
  );
  al_mux2l _3997_ (
    .a(\DFF_300.D ),
    .b(\DFF_183.Q ),
    .s(_0157_),
    .y(\DFF_183.D )
  );
  al_mux2l _3998_ (
    .a(\DFF_300.D ),
    .b(\DFF_184.Q ),
    .s(_0158_),
    .y(\DFF_184.D )
  );
  al_mux2l _3999_ (
    .a(\DFF_298.D ),
    .b(\DFF_185.Q ),
    .s(_0156_),
    .y(\DFF_185.D )
  );
  al_mux2l _4000_ (
    .a(\DFF_298.D ),
    .b(\DFF_186.Q ),
    .s(_0157_),
    .y(\DFF_186.D )
  );
  al_mux2l _4001_ (
    .a(\DFF_298.D ),
    .b(\DFF_187.Q ),
    .s(_0158_),
    .y(\DFF_187.D )
  );
  al_nand2ft _4002_ (
    .a(\DFF_201.Q ),
    .b(\DFF_1428.Q ),
    .y(_0159_)
  );
  al_ao21ftf _4003_ (
    .a(\DFF_202.Q ),
    .b(\DFF_1429.Q ),
    .c(_0159_),
    .y(_0160_)
  );
  al_ao21ftt _4004_ (
    .a(\DFF_200.Q ),
    .b(\DFF_1427.Q ),
    .c(_0160_),
    .y(_0161_)
  );
  al_inv _4005_ (
    .a(_0161_),
    .y(_0162_)
  );
  al_mux2h _4006_ (
    .a(\DFF_188.Q ),
    .b(_0162_),
    .s(_0156_),
    .y(\DFF_188.D )
  );
  al_mux2h _4007_ (
    .a(\DFF_189.Q ),
    .b(_0162_),
    .s(_0157_),
    .y(\DFF_189.D )
  );
  al_mux2h _4008_ (
    .a(\DFF_190.Q ),
    .b(_0162_),
    .s(_0158_),
    .y(\DFF_190.D )
  );
  al_nand2ft _4009_ (
    .a(\DFF_198.Q ),
    .b(\DFF_1428.Q ),
    .y(_0163_)
  );
  al_ao21ftf _4010_ (
    .a(\DFF_199.Q ),
    .b(\DFF_1429.Q ),
    .c(_0163_),
    .y(_0164_)
  );
  al_ao21ftt _4011_ (
    .a(\DFF_197.Q ),
    .b(\DFF_1427.Q ),
    .c(_0164_),
    .y(_0165_)
  );
  al_inv _4012_ (
    .a(_0165_),
    .y(_0166_)
  );
  al_mux2h _4013_ (
    .a(\DFF_191.Q ),
    .b(_0166_),
    .s(_0156_),
    .y(\DFF_191.D )
  );
  al_mux2h _4014_ (
    .a(\DFF_192.Q ),
    .b(_0166_),
    .s(_0157_),
    .y(\DFF_192.D )
  );
  al_mux2h _4015_ (
    .a(\DFF_193.Q ),
    .b(_0166_),
    .s(_0158_),
    .y(\DFF_193.D )
  );
  al_nand2 _4016_ (
    .a(\DFF_269.Q ),
    .b(\DFF_1428.Q ),
    .y(_0167_)
  );
  al_nand2 _4017_ (
    .a(\DFF_268.Q ),
    .b(\DFF_1427.Q ),
    .y(_0168_)
  );
  al_and2 _4018_ (
    .a(\DFF_270.Q ),
    .b(\DFF_1429.Q ),
    .y(_0169_)
  );
  al_and3ftt _4019_ (
    .a(_0169_),
    .b(_0167_),
    .c(_0168_),
    .y(_0170_)
  );
  al_mux2h _4020_ (
    .a(\DFF_389.Q ),
    .b(_0170_),
    .s(\DFF_1427.Q ),
    .y(\DFF_389.D )
  );
  al_mux2h _4021_ (
    .a(\DFF_390.Q ),
    .b(_0170_),
    .s(\DFF_1428.Q ),
    .y(\DFF_390.D )
  );
  al_mux2h _4022_ (
    .a(\DFF_391.Q ),
    .b(_0170_),
    .s(\DFF_1429.Q ),
    .y(\DFF_391.D )
  );
  al_nand2 _4023_ (
    .a(\DFF_278.Q ),
    .b(\DFF_1428.Q ),
    .y(_0171_)
  );
  al_and2 _4024_ (
    .a(\DFF_277.Q ),
    .b(\DFF_1427.Q ),
    .y(_0172_)
  );
  al_and2 _4025_ (
    .a(\DFF_279.Q ),
    .b(\DFF_1429.Q ),
    .y(_0173_)
  );
  al_and3fft _4026_ (
    .a(_0172_),
    .b(_0173_),
    .c(_0171_),
    .y(_0174_)
  );
  al_inv _4027_ (
    .a(_0174_),
    .y(_0175_)
  );
  al_mux2h _4028_ (
    .a(\DFF_380.Q ),
    .b(_0175_),
    .s(\DFF_1427.Q ),
    .y(\DFF_380.D )
  );
  al_mux2h _4029_ (
    .a(\DFF_381.Q ),
    .b(_0175_),
    .s(\DFF_1428.Q ),
    .y(\DFF_381.D )
  );
  al_mux2h _4030_ (
    .a(\DFF_382.Q ),
    .b(_0175_),
    .s(\DFF_1429.Q ),
    .y(\DFF_382.D )
  );
  al_inv _4031_ (
    .a(\DFF_1604.Q ),
    .y(_0176_)
  );
  al_or3 _4032_ (
    .a(\DFF_1603.Q ),
    .b(\DFF_1606.Q ),
    .c(\DFF_1605.Q ),
    .y(_0177_)
  );
  al_and3fft _4033_ (
    .a(\DFF_1602.Q ),
    .b(_0177_),
    .c(_0176_),
    .y(_0178_)
  );
  al_inv _4034_ (
    .a(_0178_),
    .y(_0179_)
  );
  al_ao21ftt _4035_ (
    .a(_0025_),
    .b(\DFF_423.Q ),
    .c(_0027_),
    .y(_0180_)
  );
  al_nand2 _4036_ (
    .a(\DFF_430.Q ),
    .b(\DFF_1505.Q ),
    .y(_0181_)
  );
  al_aoi21ttf _4037_ (
    .a(\DFF_431.Q ),
    .b(\DFF_1506.Q ),
    .c(_0181_),
    .y(_0182_)
  );
  al_aoi21ftf _4038_ (
    .a(_0025_),
    .b(\DFF_429.Q ),
    .c(_0182_),
    .y(_0183_)
  );
  al_nand3 _4039_ (
    .a(\DFF_361.Q ),
    .b(_0180_),
    .c(_0183_),
    .y(_0184_)
  );
  al_or2 _4040_ (
    .a(_0033_),
    .b(_0183_),
    .y(_0185_)
  );
  al_aoi21ftf _4041_ (
    .a(_0179_),
    .b(_0184_),
    .c(_0185_),
    .y(\DFF_433.D )
  );
  al_and3ftt _4042_ (
    .a(\DFF_458.Q ),
    .b(\DFF_459.Q ),
    .c(\DFF_1506.Q ),
    .y(_0186_)
  );
  al_oa21ttf _4043_ (
    .a(\DFF_460.Q ),
    .b(_0186_),
    .c(_0029_),
    .y(_0187_)
  );
  al_aoi21ftf _4044_ (
    .a(_0014_),
    .b(_0186_),
    .c(_0187_),
    .y(\DFF_460.D )
  );
  al_aoi21ftt _4045_ (
    .a(\DFF_508.Q ),
    .b(_0015_),
    .c(_0024_),
    .y(\DFF_508.D )
  );
  al_aoi21ftt _4046_ (
    .a(\DFF_509.Q ),
    .b(_0012_),
    .c(_0029_),
    .y(\DFF_509.D )
  );
  al_aoi21ftt _4047_ (
    .a(\DFF_510.Q ),
    .b(_0013_),
    .c(_0030_),
    .y(\DFF_510.D )
  );
  al_mux2l _4048_ (
    .a(\DFF_662.D ),
    .b(\DFF_514.Q ),
    .s(_0156_),
    .y(\DFF_514.D )
  );
  al_mux2l _4049_ (
    .a(\DFF_662.D ),
    .b(\DFF_515.Q ),
    .s(_0157_),
    .y(\DFF_515.D )
  );
  al_mux2l _4050_ (
    .a(\DFF_662.D ),
    .b(\DFF_516.Q ),
    .s(_0158_),
    .y(\DFF_516.D )
  );
  al_mux2l _4051_ (
    .a(\DFF_660.D ),
    .b(\DFF_517.Q ),
    .s(_0156_),
    .y(\DFF_517.D )
  );
  al_mux2l _4052_ (
    .a(\DFF_660.D ),
    .b(\DFF_518.Q ),
    .s(_0157_),
    .y(\DFF_518.D )
  );
  al_mux2l _4053_ (
    .a(\DFF_660.D ),
    .b(\DFF_519.Q ),
    .s(_0158_),
    .y(\DFF_519.D )
  );
  al_mux2l _4054_ (
    .a(\DFF_658.D ),
    .b(\DFF_520.Q ),
    .s(_0156_),
    .y(\DFF_520.D )
  );
  al_mux2l _4055_ (
    .a(\DFF_658.D ),
    .b(\DFF_521.Q ),
    .s(_0157_),
    .y(\DFF_521.D )
  );
  al_mux2l _4056_ (
    .a(\DFF_658.D ),
    .b(\DFF_522.Q ),
    .s(_0158_),
    .y(\DFF_522.D )
  );
  al_mux2l _4057_ (
    .a(\DFF_656.D ),
    .b(\DFF_523.Q ),
    .s(_0156_),
    .y(\DFF_523.D )
  );
  al_mux2l _4058_ (
    .a(\DFF_656.D ),
    .b(\DFF_524.Q ),
    .s(_0157_),
    .y(\DFF_524.D )
  );
  al_mux2l _4059_ (
    .a(\DFF_656.D ),
    .b(\DFF_525.Q ),
    .s(_0158_),
    .y(\DFF_525.D )
  );
  al_mux2l _4060_ (
    .a(\DFF_654.D ),
    .b(\DFF_526.Q ),
    .s(_0156_),
    .y(\DFF_526.D )
  );
  al_mux2l _4061_ (
    .a(\DFF_654.D ),
    .b(\DFF_527.Q ),
    .s(_0157_),
    .y(\DFF_527.D )
  );
  al_mux2l _4062_ (
    .a(\DFF_654.D ),
    .b(\DFF_528.Q ),
    .s(_0158_),
    .y(\DFF_528.D )
  );
  al_mux2l _4063_ (
    .a(\DFF_652.D ),
    .b(\DFF_529.Q ),
    .s(_0156_),
    .y(\DFF_529.D )
  );
  al_mux2l _4064_ (
    .a(\DFF_652.D ),
    .b(\DFF_530.Q ),
    .s(_0157_),
    .y(\DFF_530.D )
  );
  al_mux2l _4065_ (
    .a(\DFF_652.D ),
    .b(\DFF_531.Q ),
    .s(_0158_),
    .y(\DFF_531.D )
  );
  al_mux2l _4066_ (
    .a(\DFF_650.D ),
    .b(\DFF_532.Q ),
    .s(_0156_),
    .y(\DFF_532.D )
  );
  al_mux2l _4067_ (
    .a(\DFF_650.D ),
    .b(\DFF_533.Q ),
    .s(_0157_),
    .y(\DFF_533.D )
  );
  al_mux2l _4068_ (
    .a(\DFF_650.D ),
    .b(\DFF_534.Q ),
    .s(_0158_),
    .y(\DFF_534.D )
  );
  al_mux2l _4069_ (
    .a(\DFF_648.D ),
    .b(\DFF_535.Q ),
    .s(_0156_),
    .y(\DFF_535.D )
  );
  al_mux2l _4070_ (
    .a(\DFF_648.D ),
    .b(\DFF_536.Q ),
    .s(_0157_),
    .y(\DFF_536.D )
  );
  al_mux2l _4071_ (
    .a(\DFF_648.D ),
    .b(\DFF_537.Q ),
    .s(_0158_),
    .y(\DFF_537.D )
  );
  al_nand2ft _4072_ (
    .a(\DFF_551.Q ),
    .b(\DFF_1428.Q ),
    .y(_0188_)
  );
  al_and2ft _4073_ (
    .a(\DFF_550.Q ),
    .b(\DFF_1427.Q ),
    .y(_0189_)
  );
  al_nand2ft _4074_ (
    .a(\DFF_552.Q ),
    .b(\DFF_1429.Q ),
    .y(_0190_)
  );
  al_and3ftt _4075_ (
    .a(_0189_),
    .b(_0188_),
    .c(_0190_),
    .y(_0191_)
  );
  al_mux2h _4076_ (
    .a(\DFF_538.Q ),
    .b(_0191_),
    .s(_0156_),
    .y(\DFF_538.D )
  );
  al_mux2h _4077_ (
    .a(\DFF_539.Q ),
    .b(_0191_),
    .s(_0157_),
    .y(\DFF_539.D )
  );
  al_mux2h _4078_ (
    .a(\DFF_540.Q ),
    .b(_0191_),
    .s(_0158_),
    .y(\DFF_540.D )
  );
  al_nand2ft _4079_ (
    .a(\DFF_548.Q ),
    .b(\DFF_1428.Q ),
    .y(_0192_)
  );
  al_and2ft _4080_ (
    .a(\DFF_547.Q ),
    .b(\DFF_1427.Q ),
    .y(_0193_)
  );
  al_nand2ft _4081_ (
    .a(\DFF_549.Q ),
    .b(\DFF_1429.Q ),
    .y(_0194_)
  );
  al_and3ftt _4082_ (
    .a(_0193_),
    .b(_0192_),
    .c(_0194_),
    .y(_0195_)
  );
  al_mux2h _4083_ (
    .a(\DFF_541.Q ),
    .b(_0195_),
    .s(_0156_),
    .y(\DFF_541.D )
  );
  al_mux2h _4084_ (
    .a(\DFF_542.Q ),
    .b(_0195_),
    .s(_0157_),
    .y(\DFF_542.D )
  );
  al_mux2h _4085_ (
    .a(\DFF_543.Q ),
    .b(_0195_),
    .s(_0158_),
    .y(\DFF_543.D )
  );
  al_and2 _4086_ (
    .a(\DFF_619.Q ),
    .b(\DFF_1428.Q ),
    .y(_0196_)
  );
  al_and2 _4087_ (
    .a(\DFF_618.Q ),
    .b(\DFF_1427.Q ),
    .y(_0197_)
  );
  al_and2 _4088_ (
    .a(\DFF_620.Q ),
    .b(\DFF_1429.Q ),
    .y(_0198_)
  );
  al_or3 _4089_ (
    .a(_0196_),
    .b(_0197_),
    .c(_0198_),
    .y(\DFF_666.D )
  );
  al_inv _4090_ (
    .a(\DFF_666.D ),
    .y(_0199_)
  );
  al_mux2h _4091_ (
    .a(\DFF_739.Q ),
    .b(_0199_),
    .s(\DFF_1427.Q ),
    .y(\DFF_739.D )
  );
  al_mux2h _4092_ (
    .a(\DFF_740.Q ),
    .b(_0199_),
    .s(\DFF_1428.Q ),
    .y(\DFF_740.D )
  );
  al_mux2h _4093_ (
    .a(\DFF_741.Q ),
    .b(_0199_),
    .s(\DFF_1429.Q ),
    .y(\DFF_741.D )
  );
  al_nand2 _4094_ (
    .a(\DFF_628.Q ),
    .b(\DFF_1428.Q ),
    .y(_0200_)
  );
  al_and2 _4095_ (
    .a(\DFF_627.Q ),
    .b(\DFF_1427.Q ),
    .y(_0201_)
  );
  al_and2 _4096_ (
    .a(\DFF_629.Q ),
    .b(\DFF_1429.Q ),
    .y(_0202_)
  );
  al_and3fft _4097_ (
    .a(_0201_),
    .b(_0202_),
    .c(_0200_),
    .y(_0203_)
  );
  al_inv _4098_ (
    .a(_0203_),
    .y(_0204_)
  );
  al_mux2h _4099_ (
    .a(\DFF_730.Q ),
    .b(_0204_),
    .s(\DFF_1427.Q ),
    .y(\DFF_730.D )
  );
  al_mux2h _4100_ (
    .a(\DFF_731.Q ),
    .b(_0204_),
    .s(\DFF_1428.Q ),
    .y(\DFF_731.D )
  );
  al_mux2h _4101_ (
    .a(\DFF_732.Q ),
    .b(_0204_),
    .s(\DFF_1429.Q ),
    .y(\DFF_732.D )
  );
  al_nand2 _4102_ (
    .a(\DFF_780.Q ),
    .b(\DFF_1505.Q ),
    .y(_0205_)
  );
  al_aoi21ttf _4103_ (
    .a(\DFF_781.Q ),
    .b(\DFF_1506.Q ),
    .c(_0205_),
    .y(_0206_)
  );
  al_aoi21ftf _4104_ (
    .a(_0025_),
    .b(\DFF_779.Q ),
    .c(_0206_),
    .y(_0207_)
  );
  al_nand3 _4105_ (
    .a(\DFF_711.Q ),
    .b(_0054_),
    .c(_0207_),
    .y(_0208_)
  );
  al_nand2ft _4106_ (
    .a(_0207_),
    .b(_0059_),
    .y(_0209_)
  );
  al_aoi21ftf _4107_ (
    .a(_0179_),
    .b(_0208_),
    .c(_0209_),
    .y(\DFF_783.D )
  );
  al_oa21ttf _4108_ (
    .a(\DFF_810.Q ),
    .b(_0034_),
    .c(_0035_),
    .y(_0210_)
  );
  al_aoi21ftf _4109_ (
    .a(_0042_),
    .b(_0034_),
    .c(_0210_),
    .y(\DFF_810.D )
  );
  al_aoi21ftt _4110_ (
    .a(\DFF_858.Q ),
    .b(_0039_),
    .c(_0051_),
    .y(\DFF_858.D )
  );
  al_aoi21ftt _4111_ (
    .a(\DFF_859.Q ),
    .b(_0040_),
    .c(_0035_),
    .y(\DFF_859.D )
  );
  al_aoi21ftt _4112_ (
    .a(\DFF_860.Q ),
    .b(_0041_),
    .c(_0056_),
    .y(\DFF_860.D )
  );
  al_mux2l _4113_ (
    .a(\DFF_1012.D ),
    .b(\DFF_864.Q ),
    .s(_0156_),
    .y(\DFF_864.D )
  );
  al_mux2l _4114_ (
    .a(\DFF_1012.D ),
    .b(\DFF_865.Q ),
    .s(_0157_),
    .y(\DFF_865.D )
  );
  al_mux2l _4115_ (
    .a(\DFF_1012.D ),
    .b(\DFF_866.Q ),
    .s(_0158_),
    .y(\DFF_866.D )
  );
  al_mux2l _4116_ (
    .a(\DFF_1010.D ),
    .b(\DFF_867.Q ),
    .s(_0156_),
    .y(\DFF_867.D )
  );
  al_mux2l _4117_ (
    .a(\DFF_1010.D ),
    .b(\DFF_868.Q ),
    .s(_0157_),
    .y(\DFF_868.D )
  );
  al_mux2l _4118_ (
    .a(\DFF_1010.D ),
    .b(\DFF_869.Q ),
    .s(_0158_),
    .y(\DFF_869.D )
  );
  al_mux2l _4119_ (
    .a(\DFF_1008.D ),
    .b(\DFF_870.Q ),
    .s(_0156_),
    .y(\DFF_870.D )
  );
  al_mux2l _4120_ (
    .a(\DFF_1008.D ),
    .b(\DFF_871.Q ),
    .s(_0157_),
    .y(\DFF_871.D )
  );
  al_mux2l _4121_ (
    .a(\DFF_1008.D ),
    .b(\DFF_872.Q ),
    .s(_0158_),
    .y(\DFF_872.D )
  );
  al_mux2l _4122_ (
    .a(\DFF_1006.D ),
    .b(\DFF_873.Q ),
    .s(_0156_),
    .y(\DFF_873.D )
  );
  al_mux2l _4123_ (
    .a(\DFF_1006.D ),
    .b(\DFF_874.Q ),
    .s(_0157_),
    .y(\DFF_874.D )
  );
  al_mux2l _4124_ (
    .a(\DFF_1006.D ),
    .b(\DFF_875.Q ),
    .s(_0158_),
    .y(\DFF_875.D )
  );
  al_mux2l _4125_ (
    .a(\DFF_1004.D ),
    .b(\DFF_876.Q ),
    .s(_0156_),
    .y(\DFF_876.D )
  );
  al_mux2l _4126_ (
    .a(\DFF_1004.D ),
    .b(\DFF_877.Q ),
    .s(_0157_),
    .y(\DFF_877.D )
  );
  al_mux2l _4127_ (
    .a(\DFF_1004.D ),
    .b(\DFF_878.Q ),
    .s(_0158_),
    .y(\DFF_878.D )
  );
  al_mux2l _4128_ (
    .a(\DFF_1002.D ),
    .b(\DFF_879.Q ),
    .s(_0156_),
    .y(\DFF_879.D )
  );
  al_mux2l _4129_ (
    .a(\DFF_1002.D ),
    .b(\DFF_880.Q ),
    .s(_0157_),
    .y(\DFF_880.D )
  );
  al_mux2l _4130_ (
    .a(\DFF_1002.D ),
    .b(\DFF_881.Q ),
    .s(_0158_),
    .y(\DFF_881.D )
  );
  al_mux2l _4131_ (
    .a(\DFF_1000.D ),
    .b(\DFF_882.Q ),
    .s(_0156_),
    .y(\DFF_882.D )
  );
  al_mux2l _4132_ (
    .a(\DFF_1000.D ),
    .b(\DFF_883.Q ),
    .s(_0157_),
    .y(\DFF_883.D )
  );
  al_mux2l _4133_ (
    .a(\DFF_1000.D ),
    .b(\DFF_884.Q ),
    .s(_0158_),
    .y(\DFF_884.D )
  );
  al_mux2l _4134_ (
    .a(\DFF_998.D ),
    .b(\DFF_885.Q ),
    .s(_0156_),
    .y(\DFF_885.D )
  );
  al_mux2l _4135_ (
    .a(\DFF_998.D ),
    .b(\DFF_886.Q ),
    .s(_0157_),
    .y(\DFF_886.D )
  );
  al_mux2l _4136_ (
    .a(\DFF_998.D ),
    .b(\DFF_887.Q ),
    .s(_0158_),
    .y(\DFF_887.D )
  );
  al_nand2ft _4137_ (
    .a(\DFF_901.Q ),
    .b(\DFF_1428.Q ),
    .y(_0211_)
  );
  al_and2ft _4138_ (
    .a(\DFF_900.Q ),
    .b(\DFF_1427.Q ),
    .y(_0212_)
  );
  al_nand2ft _4139_ (
    .a(\DFF_902.Q ),
    .b(\DFF_1429.Q ),
    .y(_0213_)
  );
  al_and3ftt _4140_ (
    .a(_0212_),
    .b(_0211_),
    .c(_0213_),
    .y(_0214_)
  );
  al_mux2h _4141_ (
    .a(\DFF_888.Q ),
    .b(_0214_),
    .s(_0156_),
    .y(\DFF_888.D )
  );
  al_mux2h _4142_ (
    .a(\DFF_889.Q ),
    .b(_0214_),
    .s(_0157_),
    .y(\DFF_889.D )
  );
  al_mux2h _4143_ (
    .a(\DFF_890.Q ),
    .b(_0214_),
    .s(_0158_),
    .y(\DFF_890.D )
  );
  al_and2ft _4144_ (
    .a(\DFF_897.Q ),
    .b(\DFF_1427.Q ),
    .y(_0215_)
  );
  al_nand2ft _4145_ (
    .a(\DFF_898.Q ),
    .b(\DFF_1428.Q ),
    .y(_0216_)
  );
  al_ao21ftf _4146_ (
    .a(\DFF_899.Q ),
    .b(\DFF_1429.Q ),
    .c(_0216_),
    .y(_0217_)
  );
  al_nor2 _4147_ (
    .a(_0215_),
    .b(_0217_),
    .y(_0218_)
  );
  al_mux2h _4148_ (
    .a(\DFF_891.Q ),
    .b(_0218_),
    .s(_0156_),
    .y(\DFF_891.D )
  );
  al_mux2h _4149_ (
    .a(\DFF_892.Q ),
    .b(_0218_),
    .s(_0157_),
    .y(\DFF_892.D )
  );
  al_mux2h _4150_ (
    .a(\DFF_893.Q ),
    .b(_0218_),
    .s(_0158_),
    .y(\DFF_893.D )
  );
  al_nand2 _4151_ (
    .a(\DFF_969.Q ),
    .b(\DFF_1428.Q ),
    .y(_0219_)
  );
  al_nand2 _4152_ (
    .a(\DFF_968.Q ),
    .b(\DFF_1427.Q ),
    .y(_0220_)
  );
  al_and2 _4153_ (
    .a(\DFF_970.Q ),
    .b(\DFF_1429.Q ),
    .y(_0221_)
  );
  al_and3ftt _4154_ (
    .a(_0221_),
    .b(_0219_),
    .c(_0220_),
    .y(_0222_)
  );
  al_mux2h _4155_ (
    .a(\DFF_1089.Q ),
    .b(_0222_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1089.D )
  );
  al_mux2h _4156_ (
    .a(\DFF_1090.Q ),
    .b(_0222_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1090.D )
  );
  al_mux2h _4157_ (
    .a(\DFF_1091.Q ),
    .b(_0222_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1091.D )
  );
  al_nand2 _4158_ (
    .a(\DFF_978.Q ),
    .b(\DFF_1428.Q ),
    .y(_0223_)
  );
  al_and2 _4159_ (
    .a(\DFF_977.Q ),
    .b(\DFF_1427.Q ),
    .y(_0224_)
  );
  al_and2 _4160_ (
    .a(\DFF_979.Q ),
    .b(\DFF_1429.Q ),
    .y(_0225_)
  );
  al_and3fft _4161_ (
    .a(_0224_),
    .b(_0225_),
    .c(_0223_),
    .y(_0226_)
  );
  al_inv _4162_ (
    .a(_0226_),
    .y(_0227_)
  );
  al_mux2h _4163_ (
    .a(\DFF_1080.Q ),
    .b(_0227_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1080.D )
  );
  al_mux2h _4164_ (
    .a(\DFF_1081.Q ),
    .b(_0227_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1081.D )
  );
  al_mux2h _4165_ (
    .a(\DFF_1082.Q ),
    .b(_0227_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1082.D )
  );
  al_nand2 _4166_ (
    .a(\DFF_1130.Q ),
    .b(\DFF_1505.Q ),
    .y(_0228_)
  );
  al_aoi21ttf _4167_ (
    .a(\DFF_1131.Q ),
    .b(\DFF_1506.Q ),
    .c(_0228_),
    .y(_0229_)
  );
  al_aoi21ftf _4168_ (
    .a(_0025_),
    .b(\DFF_1129.Q ),
    .c(_0229_),
    .y(_0230_)
  );
  al_nand3 _4169_ (
    .a(\DFF_1061.Q ),
    .b(_0081_),
    .c(_0230_),
    .y(_0231_)
  );
  al_or2 _4170_ (
    .a(_0086_),
    .b(_0230_),
    .y(_0232_)
  );
  al_aoi21ftf _4171_ (
    .a(_0179_),
    .b(_0231_),
    .c(_0232_),
    .y(\DFF_1133.D )
  );
  al_oa21ttf _4172_ (
    .a(\DFF_1160.Q ),
    .b(_0061_),
    .c(_0062_),
    .y(_0233_)
  );
  al_aoi21ftf _4173_ (
    .a(_0069_),
    .b(_0061_),
    .c(_0233_),
    .y(\DFF_1160.D )
  );
  al_aoi21ftt _4174_ (
    .a(\DFF_1208.Q ),
    .b(_0066_),
    .c(_0078_),
    .y(\DFF_1208.D )
  );
  al_aoi21ftt _4175_ (
    .a(\DFF_1209.Q ),
    .b(_0067_),
    .c(_0062_),
    .y(\DFF_1209.D )
  );
  al_aoi21ftt _4176_ (
    .a(\DFF_1210.Q ),
    .b(_0068_),
    .c(_0083_),
    .y(\DFF_1210.D )
  );
  al_mux2l _4177_ (
    .a(\DFF_1362.D ),
    .b(\DFF_1214.Q ),
    .s(_0156_),
    .y(\DFF_1214.D )
  );
  al_mux2l _4178_ (
    .a(\DFF_1362.D ),
    .b(\DFF_1215.Q ),
    .s(_0157_),
    .y(\DFF_1215.D )
  );
  al_mux2l _4179_ (
    .a(\DFF_1362.D ),
    .b(\DFF_1216.Q ),
    .s(_0158_),
    .y(\DFF_1216.D )
  );
  al_mux2l _4180_ (
    .a(\DFF_1360.D ),
    .b(\DFF_1217.Q ),
    .s(_0156_),
    .y(\DFF_1217.D )
  );
  al_mux2l _4181_ (
    .a(\DFF_1360.D ),
    .b(\DFF_1218.Q ),
    .s(_0157_),
    .y(\DFF_1218.D )
  );
  al_mux2l _4182_ (
    .a(\DFF_1360.D ),
    .b(\DFF_1219.Q ),
    .s(_0158_),
    .y(\DFF_1219.D )
  );
  al_mux2l _4183_ (
    .a(\DFF_1358.D ),
    .b(\DFF_1220.Q ),
    .s(_0156_),
    .y(\DFF_1220.D )
  );
  al_mux2l _4184_ (
    .a(\DFF_1358.D ),
    .b(\DFF_1221.Q ),
    .s(_0157_),
    .y(\DFF_1221.D )
  );
  al_mux2l _4185_ (
    .a(\DFF_1358.D ),
    .b(\DFF_1222.Q ),
    .s(_0158_),
    .y(\DFF_1222.D )
  );
  al_mux2l _4186_ (
    .a(\DFF_1356.D ),
    .b(\DFF_1223.Q ),
    .s(_0156_),
    .y(\DFF_1223.D )
  );
  al_mux2l _4187_ (
    .a(\DFF_1356.D ),
    .b(\DFF_1224.Q ),
    .s(_0157_),
    .y(\DFF_1224.D )
  );
  al_mux2l _4188_ (
    .a(\DFF_1356.D ),
    .b(\DFF_1225.Q ),
    .s(_0158_),
    .y(\DFF_1225.D )
  );
  al_mux2l _4189_ (
    .a(\DFF_1354.D ),
    .b(\DFF_1226.Q ),
    .s(_0156_),
    .y(\DFF_1226.D )
  );
  al_mux2l _4190_ (
    .a(\DFF_1354.D ),
    .b(\DFF_1227.Q ),
    .s(_0157_),
    .y(\DFF_1227.D )
  );
  al_mux2l _4191_ (
    .a(\DFF_1354.D ),
    .b(\DFF_1228.Q ),
    .s(_0158_),
    .y(\DFF_1228.D )
  );
  al_mux2l _4192_ (
    .a(\DFF_1352.D ),
    .b(\DFF_1229.Q ),
    .s(_0156_),
    .y(\DFF_1229.D )
  );
  al_mux2l _4193_ (
    .a(\DFF_1352.D ),
    .b(\DFF_1230.Q ),
    .s(_0157_),
    .y(\DFF_1230.D )
  );
  al_mux2l _4194_ (
    .a(\DFF_1352.D ),
    .b(\DFF_1231.Q ),
    .s(_0158_),
    .y(\DFF_1231.D )
  );
  al_mux2l _4195_ (
    .a(\DFF_1350.D ),
    .b(\DFF_1232.Q ),
    .s(_0156_),
    .y(\DFF_1232.D )
  );
  al_mux2l _4196_ (
    .a(\DFF_1350.D ),
    .b(\DFF_1233.Q ),
    .s(_0157_),
    .y(\DFF_1233.D )
  );
  al_mux2l _4197_ (
    .a(\DFF_1350.D ),
    .b(\DFF_1234.Q ),
    .s(_0158_),
    .y(\DFF_1234.D )
  );
  al_mux2l _4198_ (
    .a(\DFF_1348.D ),
    .b(\DFF_1235.Q ),
    .s(_0156_),
    .y(\DFF_1235.D )
  );
  al_mux2l _4199_ (
    .a(\DFF_1348.D ),
    .b(\DFF_1236.Q ),
    .s(_0157_),
    .y(\DFF_1236.D )
  );
  al_mux2l _4200_ (
    .a(\DFF_1348.D ),
    .b(\DFF_1237.Q ),
    .s(_0158_),
    .y(\DFF_1237.D )
  );
  al_nand2ft _4201_ (
    .a(\DFF_1251.Q ),
    .b(\DFF_1428.Q ),
    .y(_0234_)
  );
  al_aoi21ftf _4202_ (
    .a(\DFF_1252.Q ),
    .b(\DFF_1429.Q ),
    .c(_0234_),
    .y(_0235_)
  );
  al_ao21ftf _4203_ (
    .a(\DFF_1250.Q ),
    .b(\DFF_1427.Q ),
    .c(_0235_),
    .y(_0236_)
  );
  al_inv _4204_ (
    .a(_0236_),
    .y(_0237_)
  );
  al_mux2h _4205_ (
    .a(\DFF_1238.Q ),
    .b(_0237_),
    .s(_0156_),
    .y(\DFF_1238.D )
  );
  al_mux2h _4206_ (
    .a(\DFF_1239.Q ),
    .b(_0237_),
    .s(_0157_),
    .y(\DFF_1239.D )
  );
  al_mux2h _4207_ (
    .a(\DFF_1240.Q ),
    .b(_0237_),
    .s(_0158_),
    .y(\DFF_1240.D )
  );
  al_nand2ft _4208_ (
    .a(\DFF_1248.Q ),
    .b(\DFF_1428.Q ),
    .y(_0238_)
  );
  al_ao21ftf _4209_ (
    .a(\DFF_1249.Q ),
    .b(\DFF_1429.Q ),
    .c(_0238_),
    .y(_0239_)
  );
  al_ao21ftt _4210_ (
    .a(\DFF_1247.Q ),
    .b(\DFF_1427.Q ),
    .c(_0239_),
    .y(_0240_)
  );
  al_inv _4211_ (
    .a(_0240_),
    .y(_0241_)
  );
  al_mux2h _4212_ (
    .a(\DFF_1241.Q ),
    .b(_0241_),
    .s(_0156_),
    .y(\DFF_1241.D )
  );
  al_mux2h _4213_ (
    .a(\DFF_1242.Q ),
    .b(_0241_),
    .s(_0157_),
    .y(\DFF_1242.D )
  );
  al_mux2h _4214_ (
    .a(\DFF_1243.Q ),
    .b(_0241_),
    .s(_0158_),
    .y(\DFF_1243.D )
  );
  al_nand2 _4215_ (
    .a(\DFF_1319.Q ),
    .b(\DFF_1428.Q ),
    .y(_0242_)
  );
  al_nand2 _4216_ (
    .a(\DFF_1318.Q ),
    .b(\DFF_1427.Q ),
    .y(_0243_)
  );
  al_and2 _4217_ (
    .a(\DFF_1320.Q ),
    .b(\DFF_1429.Q ),
    .y(_0244_)
  );
  al_and3ftt _4218_ (
    .a(_0244_),
    .b(_0242_),
    .c(_0243_),
    .y(_0245_)
  );
  al_mux2h _4219_ (
    .a(\DFF_1439.Q ),
    .b(_0245_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1439.D )
  );
  al_mux2h _4220_ (
    .a(\DFF_1440.Q ),
    .b(_0245_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1440.D )
  );
  al_mux2h _4221_ (
    .a(\DFF_1441.Q ),
    .b(_0245_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1441.D )
  );
  al_inv _4222_ (
    .a(\DFF_1428.Q ),
    .y(_0246_)
  );
  al_nand2 _4223_ (
    .a(\DFF_1329.Q ),
    .b(\DFF_1429.Q ),
    .y(_0247_)
  );
  al_aoi21ttf _4224_ (
    .a(\DFF_1327.Q ),
    .b(\DFF_1427.Q ),
    .c(_0247_),
    .y(_0248_)
  );
  al_ao21ftf _4225_ (
    .a(_0246_),
    .b(\DFF_1328.Q ),
    .c(_0248_),
    .y(_0249_)
  );
  al_mux2h _4226_ (
    .a(\DFF_1430.Q ),
    .b(_0249_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1430.D )
  );
  al_mux2h _4227_ (
    .a(\DFF_1431.Q ),
    .b(_0249_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1431.D )
  );
  al_mux2h _4228_ (
    .a(\DFF_1432.Q ),
    .b(_0249_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1432.D )
  );
  al_nand2 _4229_ (
    .a(\DFF_1480.Q ),
    .b(\DFF_1505.Q ),
    .y(_0250_)
  );
  al_aoi21ttf _4230_ (
    .a(\DFF_1481.Q ),
    .b(\DFF_1506.Q ),
    .c(_0250_),
    .y(_0251_)
  );
  al_aoi21ftf _4231_ (
    .a(_0025_),
    .b(\DFF_1479.Q ),
    .c(_0251_),
    .y(_0252_)
  );
  al_or3fft _4232_ (
    .a(\DFF_1411.Q ),
    .b(_0252_),
    .c(_0107_),
    .y(_0253_)
  );
  al_or2 _4233_ (
    .a(_0111_),
    .b(_0252_),
    .y(_0254_)
  );
  al_aoi21ftf _4234_ (
    .a(_0179_),
    .b(_0253_),
    .c(_0254_),
    .y(\DFF_1483.D )
  );
  al_oa21ttf _4235_ (
    .a(\DFF_1510.Q ),
    .b(_0087_),
    .c(_0088_),
    .y(_0255_)
  );
  al_aoi21ftf _4236_ (
    .a(_0095_),
    .b(_0087_),
    .c(_0255_),
    .y(\DFF_1510.D )
  );
  al_aoi21ftt _4237_ (
    .a(\DFF_1558.Q ),
    .b(_0092_),
    .c(_0104_),
    .y(\DFF_1558.D )
  );
  al_aoi21ftt _4238_ (
    .a(\DFF_1559.Q ),
    .b(_0093_),
    .c(_0088_),
    .y(\DFF_1559.D )
  );
  al_aoi21ftt _4239_ (
    .a(\DFF_1560.Q ),
    .b(_0094_),
    .c(_0108_),
    .y(\DFF_1560.D )
  );
  al_nor2 _4240_ (
    .a(\DFF_6.Q ),
    .b(\DFF_9.Q ),
    .y(_0256_)
  );
  al_and2ft _4241_ (
    .a(\DFF_4.Q ),
    .b(\DFF_10.Q ),
    .y(_0257_)
  );
  al_and3 _4242_ (
    .a(\DFF_7.Q ),
    .b(\DFF_8.Q ),
    .c(_0257_),
    .y(_0258_)
  );
  al_and2 _4243_ (
    .a(\DFF_5.Q ),
    .b(\DFF_3.Q ),
    .y(_0259_)
  );
  al_nand3 _4244_ (
    .a(_0256_),
    .b(_0259_),
    .c(_0258_),
    .y(_0260_)
  );
  al_and2ft _4245_ (
    .a(\DFF_17.Q ),
    .b(_0260_),
    .y(_0261_)
  );
  al_ao21 _4246_ (
    .a(\DFF_4.Q ),
    .b(\DFF_3.Q ),
    .c(\DFF_5.Q ),
    .y(_0262_)
  );
  al_and3 _4247_ (
    .a(\DFF_4.Q ),
    .b(\DFF_5.Q ),
    .c(\DFF_3.Q ),
    .y(_0263_)
  );
  al_and3ftt _4248_ (
    .a(_0263_),
    .b(_0262_),
    .c(_0261_),
    .y(\DFF_5.D )
  );
  al_and2ft _4249_ (
    .a(\DFF_284.Q ),
    .b(\DFF_1428.Q ),
    .y(_0264_)
  );
  al_and2ft _4250_ (
    .a(\DFF_283.Q ),
    .b(\DFF_1427.Q ),
    .y(_0265_)
  );
  al_nand2ft _4251_ (
    .a(\DFF_285.Q ),
    .b(\DFF_1429.Q ),
    .y(_0266_)
  );
  al_nand3fft _4252_ (
    .a(_0264_),
    .b(_0265_),
    .c(_0266_),
    .y(_0267_)
  );
  al_nand2ft _4253_ (
    .a(\DFF_290.Q ),
    .b(\DFF_1428.Q ),
    .y(_0268_)
  );
  al_aoi21ftf _4254_ (
    .a(\DFF_291.Q ),
    .b(\DFF_1429.Q ),
    .c(_0268_),
    .y(_0269_)
  );
  al_aoi21ftf _4255_ (
    .a(\DFF_289.Q ),
    .b(\DFF_1427.Q ),
    .c(_0269_),
    .y(_0270_)
  );
  al_nand2ft _4256_ (
    .a(\DFF_287.Q ),
    .b(\DFF_1428.Q ),
    .y(_0271_)
  );
  al_aoi21ftf _4257_ (
    .a(\DFF_288.Q ),
    .b(\DFF_1429.Q ),
    .c(_0271_),
    .y(_0272_)
  );
  al_ao21ftf _4258_ (
    .a(\DFF_286.Q ),
    .b(\DFF_1427.Q ),
    .c(_0272_),
    .y(_0273_)
  );
  al_and3fft _4259_ (
    .a(_0267_),
    .b(_0270_),
    .c(_0273_),
    .y(_0274_)
  );
  al_mux2h _4260_ (
    .a(\DFF_384.Q ),
    .b(_0274_),
    .s(\DFF_1428.Q ),
    .y(\DFF_384.D )
  );
  al_mux2h _4261_ (
    .a(\DFF_385.Q ),
    .b(_0274_),
    .s(\DFF_1429.Q ),
    .y(\DFF_385.D )
  );
  al_and3fft _4262_ (
    .a(_0267_),
    .b(_0273_),
    .c(_0270_),
    .y(_0275_)
  );
  al_mux2h _4263_ (
    .a(\DFF_392.Q ),
    .b(_0275_),
    .s(\DFF_1427.Q ),
    .y(\DFF_392.D )
  );
  al_mux2h _4264_ (
    .a(\DFF_393.Q ),
    .b(_0275_),
    .s(\DFF_1428.Q ),
    .y(\DFF_393.D )
  );
  al_mux2h _4265_ (
    .a(\DFF_394.Q ),
    .b(_0275_),
    .s(\DFF_1429.Q ),
    .y(\DFF_394.D )
  );
  al_nor3ftt _4266_ (
    .a(_0267_),
    .b(_0273_),
    .c(_0270_),
    .y(_0276_)
  );
  al_mux2h _4267_ (
    .a(\DFF_386.Q ),
    .b(_0276_),
    .s(\DFF_1427.Q ),
    .y(\DFF_386.D )
  );
  al_mux2h _4268_ (
    .a(\DFF_387.Q ),
    .b(_0276_),
    .s(\DFF_1428.Q ),
    .y(\DFF_387.D )
  );
  al_mux2h _4269_ (
    .a(\DFF_388.Q ),
    .b(_0276_),
    .s(\DFF_1429.Q ),
    .y(\DFF_388.D )
  );
  al_mux2h _4270_ (
    .a(\DFF_383.Q ),
    .b(_0274_),
    .s(\DFF_1427.Q ),
    .y(\DFF_383.D )
  );
  al_and3 _4271_ (
    .a(\DFF_460.Q ),
    .b(\DFF_461.Q ),
    .c(_0186_),
    .y(_0277_)
  );
  al_ao21 _4272_ (
    .a(\DFF_460.Q ),
    .b(_0186_),
    .c(\DFF_461.Q ),
    .y(_0278_)
  );
  al_and3fft _4273_ (
    .a(_0029_),
    .b(_0277_),
    .c(_0278_),
    .y(\DFF_461.D )
  );
  al_nand2ft _4274_ (
    .a(\DFF_633.Q ),
    .b(\DFF_1427.Q ),
    .y(_0279_)
  );
  al_aoi21ftf _4275_ (
    .a(\DFF_635.Q ),
    .b(\DFF_1429.Q ),
    .c(_0279_),
    .y(_0280_)
  );
  al_aoi21ftf _4276_ (
    .a(\DFF_634.Q ),
    .b(\DFF_1428.Q ),
    .c(_0280_),
    .y(_0281_)
  );
  al_nand2ft _4277_ (
    .a(\DFF_640.Q ),
    .b(\DFF_1428.Q ),
    .y(_0282_)
  );
  al_aoi21ftf _4278_ (
    .a(\DFF_641.Q ),
    .b(\DFF_1429.Q ),
    .c(_0282_),
    .y(_0283_)
  );
  al_aoi21ftf _4279_ (
    .a(\DFF_639.Q ),
    .b(\DFF_1427.Q ),
    .c(_0283_),
    .y(_0284_)
  );
  al_nand2ft _4280_ (
    .a(\DFF_637.Q ),
    .b(\DFF_1428.Q ),
    .y(_0285_)
  );
  al_aoi21ftf _4281_ (
    .a(\DFF_638.Q ),
    .b(\DFF_1429.Q ),
    .c(_0285_),
    .y(_0286_)
  );
  al_ao21ftf _4282_ (
    .a(\DFF_636.Q ),
    .b(\DFF_1427.Q ),
    .c(_0286_),
    .y(_0287_)
  );
  al_and3ftt _4283_ (
    .a(_0284_),
    .b(_0281_),
    .c(_0287_),
    .y(_0288_)
  );
  al_mux2h _4284_ (
    .a(\DFF_734.Q ),
    .b(_0288_),
    .s(\DFF_1428.Q ),
    .y(\DFF_734.D )
  );
  al_mux2h _4285_ (
    .a(\DFF_735.Q ),
    .b(_0288_),
    .s(\DFF_1429.Q ),
    .y(\DFF_735.D )
  );
  al_nand3ftt _4286_ (
    .a(_0287_),
    .b(_0281_),
    .c(_0284_),
    .y(_0289_)
  );
  al_inv _4287_ (
    .a(_0289_),
    .y(_0290_)
  );
  al_mux2h _4288_ (
    .a(\DFF_742.Q ),
    .b(_0290_),
    .s(\DFF_1427.Q ),
    .y(\DFF_742.D )
  );
  al_mux2h _4289_ (
    .a(\DFF_743.Q ),
    .b(_0290_),
    .s(\DFF_1428.Q ),
    .y(\DFF_743.D )
  );
  al_mux2h _4290_ (
    .a(\DFF_744.Q ),
    .b(_0290_),
    .s(\DFF_1429.Q ),
    .y(\DFF_744.D )
  );
  al_or2 _4291_ (
    .a(_0287_),
    .b(_0284_),
    .y(_0291_)
  );
  al_nor2 _4292_ (
    .a(_0281_),
    .b(_0291_),
    .y(_0292_)
  );
  al_mux2h _4293_ (
    .a(\DFF_736.Q ),
    .b(_0292_),
    .s(\DFF_1427.Q ),
    .y(\DFF_736.D )
  );
  al_mux2h _4294_ (
    .a(\DFF_737.Q ),
    .b(_0292_),
    .s(\DFF_1428.Q ),
    .y(\DFF_737.D )
  );
  al_mux2h _4295_ (
    .a(\DFF_738.Q ),
    .b(_0292_),
    .s(\DFF_1429.Q ),
    .y(\DFF_738.D )
  );
  al_mux2h _4296_ (
    .a(\DFF_733.Q ),
    .b(_0288_),
    .s(\DFF_1427.Q ),
    .y(\DFF_733.D )
  );
  al_and3 _4297_ (
    .a(\DFF_810.Q ),
    .b(\DFF_811.Q ),
    .c(_0034_),
    .y(_0293_)
  );
  al_ao21 _4298_ (
    .a(\DFF_810.Q ),
    .b(_0034_),
    .c(\DFF_811.Q ),
    .y(_0294_)
  );
  al_and3fft _4299_ (
    .a(_0035_),
    .b(_0293_),
    .c(_0294_),
    .y(\DFF_811.D )
  );
  al_nand2ft _4300_ (
    .a(\DFF_984.Q ),
    .b(\DFF_1428.Q ),
    .y(_0295_)
  );
  al_nand2ft _4301_ (
    .a(\DFF_983.Q ),
    .b(\DFF_1427.Q ),
    .y(_0296_)
  );
  al_and2ft _4302_ (
    .a(\DFF_985.Q ),
    .b(\DFF_1429.Q ),
    .y(_0297_)
  );
  al_and3ftt _4303_ (
    .a(_0297_),
    .b(_0295_),
    .c(_0296_),
    .y(_0298_)
  );
  al_nand2ft _4304_ (
    .a(\DFF_990.Q ),
    .b(\DFF_1428.Q ),
    .y(_0299_)
  );
  al_aoi21ftf _4305_ (
    .a(\DFF_991.Q ),
    .b(\DFF_1429.Q ),
    .c(_0299_),
    .y(_0300_)
  );
  al_aoi21ftf _4306_ (
    .a(\DFF_989.Q ),
    .b(\DFF_1427.Q ),
    .c(_0300_),
    .y(_0301_)
  );
  al_nand2ft _4307_ (
    .a(\DFF_988.Q ),
    .b(\DFF_1429.Q ),
    .y(_0302_)
  );
  al_aoi21ftf _4308_ (
    .a(\DFF_986.Q ),
    .b(\DFF_1427.Q ),
    .c(_0302_),
    .y(_0303_)
  );
  al_ao21ftf _4309_ (
    .a(\DFF_987.Q ),
    .b(\DFF_1428.Q ),
    .c(_0303_),
    .y(_0304_)
  );
  al_nor3fft _4310_ (
    .a(_0298_),
    .b(_0304_),
    .c(_0301_),
    .y(_0305_)
  );
  al_mux2h _4311_ (
    .a(\DFF_1084.Q ),
    .b(_0305_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1084.D )
  );
  al_mux2h _4312_ (
    .a(\DFF_1085.Q ),
    .b(_0305_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1085.D )
  );
  al_ao21ftf _4313_ (
    .a(\DFF_989.Q ),
    .b(\DFF_1427.Q ),
    .c(_0300_),
    .y(_0306_)
  );
  al_nor3ftt _4314_ (
    .a(_0298_),
    .b(_0306_),
    .c(_0304_),
    .y(_0307_)
  );
  al_mux2h _4315_ (
    .a(\DFF_1092.Q ),
    .b(_0307_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1092.D )
  );
  al_mux2h _4316_ (
    .a(\DFF_1093.Q ),
    .b(_0307_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1093.D )
  );
  al_mux2h _4317_ (
    .a(\DFF_1094.Q ),
    .b(_0307_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1094.D )
  );
  al_and3fft _4318_ (
    .a(_0298_),
    .b(_0304_),
    .c(_0306_),
    .y(_0308_)
  );
  al_mux2h _4319_ (
    .a(\DFF_1086.Q ),
    .b(_0308_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1086.D )
  );
  al_mux2h _4320_ (
    .a(\DFF_1087.Q ),
    .b(_0308_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1087.D )
  );
  al_mux2h _4321_ (
    .a(\DFF_1088.Q ),
    .b(_0308_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1088.D )
  );
  al_mux2h _4322_ (
    .a(\DFF_1083.Q ),
    .b(_0305_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1083.D )
  );
  al_and3 _4323_ (
    .a(\DFF_1160.Q ),
    .b(\DFF_1161.Q ),
    .c(_0061_),
    .y(_0309_)
  );
  al_ao21 _4324_ (
    .a(\DFF_1160.Q ),
    .b(_0061_),
    .c(\DFF_1161.Q ),
    .y(_0310_)
  );
  al_and3fft _4325_ (
    .a(_0062_),
    .b(_0309_),
    .c(_0310_),
    .y(\DFF_1161.D )
  );
  al_and2ft _4326_ (
    .a(\DFF_1334.Q ),
    .b(\DFF_1428.Q ),
    .y(_0311_)
  );
  al_and2ft _4327_ (
    .a(\DFF_1333.Q ),
    .b(\DFF_1427.Q ),
    .y(_0312_)
  );
  al_nand2ft _4328_ (
    .a(\DFF_1335.Q ),
    .b(\DFF_1429.Q ),
    .y(_0313_)
  );
  al_nand3fft _4329_ (
    .a(_0311_),
    .b(_0312_),
    .c(_0313_),
    .y(_0314_)
  );
  al_nand2ft _4330_ (
    .a(\DFF_1340.Q ),
    .b(\DFF_1428.Q ),
    .y(_0315_)
  );
  al_aoi21ftf _4331_ (
    .a(\DFF_1341.Q ),
    .b(\DFF_1429.Q ),
    .c(_0315_),
    .y(_0316_)
  );
  al_aoi21ftf _4332_ (
    .a(\DFF_1339.Q ),
    .b(\DFF_1427.Q ),
    .c(_0316_),
    .y(_0317_)
  );
  al_nand2ft _4333_ (
    .a(\DFF_1337.Q ),
    .b(\DFF_1428.Q ),
    .y(_0318_)
  );
  al_aoi21ftf _4334_ (
    .a(\DFF_1338.Q ),
    .b(\DFF_1429.Q ),
    .c(_0318_),
    .y(_0319_)
  );
  al_ao21ftf _4335_ (
    .a(\DFF_1336.Q ),
    .b(\DFF_1427.Q ),
    .c(_0319_),
    .y(_0320_)
  );
  al_and3fft _4336_ (
    .a(_0314_),
    .b(_0317_),
    .c(_0320_),
    .y(_0321_)
  );
  al_mux2h _4337_ (
    .a(\DFF_1434.Q ),
    .b(_0321_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1434.D )
  );
  al_mux2h _4338_ (
    .a(\DFF_1435.Q ),
    .b(_0321_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1435.D )
  );
  al_and3fft _4339_ (
    .a(_0314_),
    .b(_0320_),
    .c(_0317_),
    .y(_0322_)
  );
  al_mux2h _4340_ (
    .a(\DFF_1442.Q ),
    .b(_0322_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1442.D )
  );
  al_mux2h _4341_ (
    .a(\DFF_1443.Q ),
    .b(_0322_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1443.D )
  );
  al_mux2h _4342_ (
    .a(\DFF_1444.Q ),
    .b(_0322_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1444.D )
  );
  al_nor3ftt _4343_ (
    .a(_0314_),
    .b(_0320_),
    .c(_0317_),
    .y(_0323_)
  );
  al_mux2h _4344_ (
    .a(\DFF_1436.Q ),
    .b(_0323_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1436.D )
  );
  al_mux2h _4345_ (
    .a(\DFF_1437.Q ),
    .b(_0323_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1437.D )
  );
  al_mux2h _4346_ (
    .a(\DFF_1438.Q ),
    .b(_0323_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1438.D )
  );
  al_mux2h _4347_ (
    .a(\DFF_1433.Q ),
    .b(_0321_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1433.D )
  );
  al_and3 _4348_ (
    .a(\DFF_1510.Q ),
    .b(\DFF_1511.Q ),
    .c(_0087_),
    .y(_0324_)
  );
  al_ao21 _4349_ (
    .a(\DFF_1510.Q ),
    .b(_0087_),
    .c(\DFF_1511.Q ),
    .y(_0325_)
  );
  al_and3fft _4350_ (
    .a(_0088_),
    .b(_0324_),
    .c(_0325_),
    .y(\DFF_1511.D )
  );
  al_inv _4351_ (
    .a(\DFF_11.Q ),
    .y(_0326_)
  );
  al_nor2 _4352_ (
    .a(_0326_),
    .b(_0260_),
    .y(_0327_)
  );
  al_and3fft _4353_ (
    .a(\DFF_12.Q ),
    .b(\DFF_13.Q ),
    .c(\DFF_14.Q ),
    .y(_0328_)
  );
  al_aoi21 _4354_ (
    .a(_0328_),
    .b(_0327_),
    .c(\DFF_17.Q ),
    .y(_0329_)
  );
  al_and3fft _4355_ (
    .a(_0326_),
    .b(_0260_),
    .c(\DFF_12.Q ),
    .y(_0330_)
  );
  al_oai21ftf _4356_ (
    .a(\DFF_11.Q ),
    .b(_0260_),
    .c(\DFF_12.Q ),
    .y(_0331_)
  );
  al_and3ftt _4357_ (
    .a(_0330_),
    .b(_0331_),
    .c(_0329_),
    .y(\DFF_12.D )
  );
  al_or2 _4358_ (
    .a(\DFF_6.Q ),
    .b(_0263_),
    .y(_0332_)
  );
  al_and2 _4359_ (
    .a(\DFF_6.Q ),
    .b(_0263_),
    .y(_0333_)
  );
  al_and3ftt _4360_ (
    .a(_0333_),
    .b(_0332_),
    .c(_0261_),
    .y(\DFF_6.D )
  );
  al_and3 _4361_ (
    .a(\DFF_1607.Q ),
    .b(\DFF_1563.Q ),
    .c(_0006_),
    .y(_0334_)
  );
  al_and3fft _4362_ (
    .a(\DFF_1609.Q ),
    .b(\DFF_1608.Q ),
    .c(\DFF_1610.Q ),
    .y(_0335_)
  );
  al_aoi21 _4363_ (
    .a(_0335_),
    .b(_0334_),
    .c(g3234),
    .y(_0336_)
  );
  al_and2 _4364_ (
    .a(\DFF_1608.Q ),
    .b(_0334_),
    .y(_0337_)
  );
  al_or2 _4365_ (
    .a(\DFF_1608.Q ),
    .b(_0334_),
    .y(_0338_)
  );
  al_and3ftt _4366_ (
    .a(_0337_),
    .b(_0338_),
    .c(_0336_),
    .y(\DFF_1608.D )
  );
  al_aoi21 _4367_ (
    .a(\DFF_1563.Q ),
    .b(_0006_),
    .c(g3234),
    .y(_0339_)
  );
  al_and3 _4368_ (
    .a(\DFF_1600.Q ),
    .b(\DFF_1601.Q ),
    .c(\DFF_1563.Q ),
    .y(_0340_)
  );
  al_nand2 _4369_ (
    .a(\DFF_1602.Q ),
    .b(_0340_),
    .y(_0341_)
  );
  al_or2 _4370_ (
    .a(\DFF_1602.Q ),
    .b(_0340_),
    .y(_0342_)
  );
  al_and3 _4371_ (
    .a(_0341_),
    .b(_0342_),
    .c(_0339_),
    .y(\DFF_1602.D )
  );
  al_inv _4372_ (
    .a(\DFF_236.Q ),
    .y(_0343_)
  );
  al_inv _4373_ (
    .a(\DFF_1429.Q ),
    .y(_0344_)
  );
  al_or3 _4374_ (
    .a(\DFF_7.Q ),
    .b(\DFF_8.Q ),
    .c(\DFF_10.Q ),
    .y(_0345_)
  );
  al_aoi21ftt _4375_ (
    .a(_0345_),
    .b(_0256_),
    .c(_0344_),
    .y(_0346_)
  );
  al_aoi21ttf _4376_ (
    .a(\DFF_1302.Q ),
    .b(\DFF_1429.Q ),
    .c(\DFF_236.Q ),
    .y(_0347_)
  );
  al_mux2l _4377_ (
    .a(_0343_),
    .b(_0347_),
    .s(_0346_),
    .y(\DFF_236.D )
  );
  al_mux2h _4378_ (
    .a(\DFF_317.Q ),
    .b(\DFF_453.D ),
    .s(g3229),
    .y(\DFF_452.D )
  );
  al_and2 _4379_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_368.Q ),
    .y(_0348_)
  );
  al_and2 _4380_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_366.Q ),
    .y(_0349_)
  );
  al_and2 _4381_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_370.Q ),
    .y(_0350_)
  );
  al_or3 _4382_ (
    .a(_0348_),
    .b(_0349_),
    .c(_0350_),
    .y(_0351_)
  );
  al_nand2 _4383_ (
    .a(\DFF_364.Q ),
    .b(\DFF_160.Q ),
    .y(_0352_)
  );
  al_inv _4384_ (
    .a(\DFF_1505.Q ),
    .y(_0353_)
  );
  al_nand2 _4385_ (
    .a(\DFF_417.Q ),
    .b(\DFF_1504.Q ),
    .y(_0354_)
  );
  al_aoi21ttf _4386_ (
    .a(\DFF_419.Q ),
    .b(\DFF_1506.Q ),
    .c(_0354_),
    .y(_0355_)
  );
  al_aoi21ftf _4387_ (
    .a(_0353_),
    .b(\DFF_418.Q ),
    .c(_0355_),
    .y(_0356_)
  );
  al_ao21ftf _4388_ (
    .a(_0352_),
    .b(_0351_),
    .c(_0356_),
    .y(_0357_)
  );
  al_and2ft _4389_ (
    .a(_0008_),
    .b(_0357_),
    .y(_0358_)
  );
  al_mux2h _4390_ (
    .a(\DFF_417.Q ),
    .b(_0358_),
    .s(\DFF_1504.Q ),
    .y(\DFF_417.D )
  );
  al_mux2h _4391_ (
    .a(\DFF_418.Q ),
    .b(_0358_),
    .s(\DFF_1505.Q ),
    .y(\DFF_418.D )
  );
  al_mux2h _4392_ (
    .a(\DFF_419.Q ),
    .b(_0358_),
    .s(\DFF_1506.Q ),
    .y(\DFF_419.D )
  );
  al_and2 _4393_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_374.Q ),
    .y(_0359_)
  );
  al_and2 _4394_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_372.Q ),
    .y(_0360_)
  );
  al_and2 _4395_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_376.Q ),
    .y(_0361_)
  );
  al_or3 _4396_ (
    .a(_0359_),
    .b(_0360_),
    .c(_0361_),
    .y(_0362_)
  );
  al_nand2 _4397_ (
    .a(\DFF_397.Q ),
    .b(\DFF_160.Q ),
    .y(_0363_)
  );
  al_nand2 _4398_ (
    .a(\DFF_420.Q ),
    .b(\DFF_1504.Q ),
    .y(_0364_)
  );
  al_aoi21ttf _4399_ (
    .a(\DFF_422.Q ),
    .b(\DFF_1506.Q ),
    .c(_0364_),
    .y(_0365_)
  );
  al_aoi21ftf _4400_ (
    .a(_0353_),
    .b(\DFF_421.Q ),
    .c(_0365_),
    .y(_0366_)
  );
  al_ao21ftf _4401_ (
    .a(_0363_),
    .b(_0362_),
    .c(_0366_),
    .y(_0367_)
  );
  al_and2ft _4402_ (
    .a(_0008_),
    .b(_0367_),
    .y(_0368_)
  );
  al_mux2h _4403_ (
    .a(\DFF_420.Q ),
    .b(_0368_),
    .s(\DFF_1504.Q ),
    .y(\DFF_420.D )
  );
  al_mux2h _4404_ (
    .a(\DFF_421.Q ),
    .b(_0368_),
    .s(\DFF_1505.Q ),
    .y(\DFF_421.D )
  );
  al_mux2h _4405_ (
    .a(\DFF_422.Q ),
    .b(_0368_),
    .s(\DFF_1506.Q ),
    .y(\DFF_422.D )
  );
  al_oa21ftf _4406_ (
    .a(_0017_),
    .b(_0277_),
    .c(_0029_),
    .y(_0369_)
  );
  al_aoi21ftf _4407_ (
    .a(_0017_),
    .b(_0277_),
    .c(_0369_),
    .y(\DFF_462.D )
  );
  al_inv _4408_ (
    .a(\DFF_586.Q ),
    .y(_0370_)
  );
  al_aoi21ttf _4409_ (
    .a(\DFF_1302.Q ),
    .b(\DFF_1429.Q ),
    .c(\DFF_586.Q ),
    .y(_0371_)
  );
  al_mux2l _4410_ (
    .a(_0370_),
    .b(_0371_),
    .s(_0346_),
    .y(\DFF_586.D )
  );
  al_mux2h _4411_ (
    .a(\DFF_667.Q ),
    .b(\DFF_803.D ),
    .s(g3229),
    .y(\DFF_802.D )
  );
  al_and2 _4412_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_718.Q ),
    .y(_0372_)
  );
  al_and2 _4413_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_716.Q ),
    .y(_0373_)
  );
  al_and2 _4414_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_720.Q ),
    .y(_0374_)
  );
  al_or3 _4415_ (
    .a(_0372_),
    .b(_0373_),
    .c(_0374_),
    .y(_0375_)
  );
  al_nand2 _4416_ (
    .a(\DFF_714.Q ),
    .b(\DFF_160.Q ),
    .y(_0376_)
  );
  al_nand2 _4417_ (
    .a(\DFF_767.Q ),
    .b(\DFF_1504.Q ),
    .y(_0377_)
  );
  al_aoi21ttf _4418_ (
    .a(\DFF_769.Q ),
    .b(\DFF_1506.Q ),
    .c(_0377_),
    .y(_0378_)
  );
  al_aoi21ftf _4419_ (
    .a(_0353_),
    .b(\DFF_768.Q ),
    .c(_0378_),
    .y(_0379_)
  );
  al_ao21ftf _4420_ (
    .a(_0376_),
    .b(_0375_),
    .c(_0379_),
    .y(_0380_)
  );
  al_and2ft _4421_ (
    .a(_0008_),
    .b(_0380_),
    .y(_0381_)
  );
  al_mux2h _4422_ (
    .a(\DFF_767.Q ),
    .b(_0381_),
    .s(\DFF_1504.Q ),
    .y(\DFF_767.D )
  );
  al_mux2h _4423_ (
    .a(\DFF_768.Q ),
    .b(_0381_),
    .s(\DFF_1505.Q ),
    .y(\DFF_768.D )
  );
  al_mux2h _4424_ (
    .a(\DFF_769.Q ),
    .b(_0381_),
    .s(\DFF_1506.Q ),
    .y(\DFF_769.D )
  );
  al_and2 _4425_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_724.Q ),
    .y(_0382_)
  );
  al_and2 _4426_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_722.Q ),
    .y(_0383_)
  );
  al_and2 _4427_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_726.Q ),
    .y(_0384_)
  );
  al_or3 _4428_ (
    .a(_0382_),
    .b(_0383_),
    .c(_0384_),
    .y(_0385_)
  );
  al_nand2 _4429_ (
    .a(\DFF_747.Q ),
    .b(\DFF_160.Q ),
    .y(_0386_)
  );
  al_nand2 _4430_ (
    .a(\DFF_770.Q ),
    .b(\DFF_1504.Q ),
    .y(_0387_)
  );
  al_aoi21ttf _4431_ (
    .a(\DFF_772.Q ),
    .b(\DFF_1506.Q ),
    .c(_0387_),
    .y(_0388_)
  );
  al_aoi21ftf _4432_ (
    .a(_0353_),
    .b(\DFF_771.Q ),
    .c(_0388_),
    .y(_0389_)
  );
  al_ao21ftf _4433_ (
    .a(_0386_),
    .b(_0385_),
    .c(_0389_),
    .y(_0390_)
  );
  al_and2ft _4434_ (
    .a(_0008_),
    .b(_0390_),
    .y(_0391_)
  );
  al_mux2h _4435_ (
    .a(\DFF_770.Q ),
    .b(_0391_),
    .s(\DFF_1504.Q ),
    .y(\DFF_770.D )
  );
  al_mux2h _4436_ (
    .a(\DFF_771.Q ),
    .b(_0391_),
    .s(\DFF_1505.Q ),
    .y(\DFF_771.D )
  );
  al_mux2h _4437_ (
    .a(\DFF_772.Q ),
    .b(_0391_),
    .s(\DFF_1506.Q ),
    .y(\DFF_772.D )
  );
  al_oa21ftf _4438_ (
    .a(_0044_),
    .b(_0293_),
    .c(_0035_),
    .y(_0392_)
  );
  al_aoi21ftf _4439_ (
    .a(_0044_),
    .b(_0293_),
    .c(_0392_),
    .y(\DFF_812.D )
  );
  al_or3 _4440_ (
    .a(\DFF_6.Q ),
    .b(\DFF_9.Q ),
    .c(_0345_),
    .y(_0393_)
  );
  al_and3 _4441_ (
    .a(\DFF_936.Q ),
    .b(\DFF_1429.Q ),
    .c(_0393_),
    .y(_0394_)
  );
  al_ao21ttf _4442_ (
    .a(\DFF_1302.Q ),
    .b(\DFF_1429.Q ),
    .c(\DFF_936.Q ),
    .y(_0395_)
  );
  al_aoi21ftt _4443_ (
    .a(_0346_),
    .b(_0395_),
    .c(_0394_),
    .y(\DFF_936.D )
  );
  al_mux2h _4444_ (
    .a(\DFF_1017.Q ),
    .b(\DFF_1153.D ),
    .s(g3229),
    .y(\DFF_1152.D )
  );
  al_and2 _4445_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_1068.Q ),
    .y(_0396_)
  );
  al_and2 _4446_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_1066.Q ),
    .y(_0397_)
  );
  al_and2 _4447_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_1070.Q ),
    .y(_0398_)
  );
  al_or3 _4448_ (
    .a(_0396_),
    .b(_0397_),
    .c(_0398_),
    .y(_0399_)
  );
  al_nand2 _4449_ (
    .a(\DFF_1064.Q ),
    .b(\DFF_160.Q ),
    .y(_0400_)
  );
  al_nand2 _4450_ (
    .a(\DFF_1117.Q ),
    .b(\DFF_1504.Q ),
    .y(_0401_)
  );
  al_aoi21ttf _4451_ (
    .a(\DFF_1119.Q ),
    .b(\DFF_1506.Q ),
    .c(_0401_),
    .y(_0402_)
  );
  al_aoi21ftf _4452_ (
    .a(_0353_),
    .b(\DFF_1118.Q ),
    .c(_0402_),
    .y(_0403_)
  );
  al_ao21ftf _4453_ (
    .a(_0400_),
    .b(_0399_),
    .c(_0403_),
    .y(_0404_)
  );
  al_and2ft _4454_ (
    .a(_0008_),
    .b(_0404_),
    .y(_0405_)
  );
  al_mux2h _4455_ (
    .a(\DFF_1117.Q ),
    .b(_0405_),
    .s(\DFF_1504.Q ),
    .y(\DFF_1117.D )
  );
  al_mux2h _4456_ (
    .a(\DFF_1118.Q ),
    .b(_0405_),
    .s(\DFF_1505.Q ),
    .y(\DFF_1118.D )
  );
  al_mux2h _4457_ (
    .a(\DFF_1119.Q ),
    .b(_0405_),
    .s(\DFF_1506.Q ),
    .y(\DFF_1119.D )
  );
  al_and2 _4458_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_1074.Q ),
    .y(_0406_)
  );
  al_and2 _4459_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_1072.Q ),
    .y(_0407_)
  );
  al_and2 _4460_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_1076.Q ),
    .y(_0408_)
  );
  al_or3 _4461_ (
    .a(_0406_),
    .b(_0407_),
    .c(_0408_),
    .y(_0409_)
  );
  al_nand2 _4462_ (
    .a(\DFF_1097.Q ),
    .b(\DFF_160.Q ),
    .y(_0410_)
  );
  al_nand2 _4463_ (
    .a(\DFF_1120.Q ),
    .b(\DFF_1504.Q ),
    .y(_0411_)
  );
  al_aoi21ttf _4464_ (
    .a(\DFF_1122.Q ),
    .b(\DFF_1506.Q ),
    .c(_0411_),
    .y(_0412_)
  );
  al_aoi21ftf _4465_ (
    .a(_0353_),
    .b(\DFF_1121.Q ),
    .c(_0412_),
    .y(_0413_)
  );
  al_ao21ftf _4466_ (
    .a(_0410_),
    .b(_0409_),
    .c(_0413_),
    .y(_0414_)
  );
  al_and2ft _4467_ (
    .a(_0008_),
    .b(_0414_),
    .y(_0415_)
  );
  al_mux2h _4468_ (
    .a(\DFF_1120.Q ),
    .b(_0415_),
    .s(\DFF_1504.Q ),
    .y(\DFF_1120.D )
  );
  al_mux2h _4469_ (
    .a(\DFF_1121.Q ),
    .b(_0415_),
    .s(\DFF_1505.Q ),
    .y(\DFF_1121.D )
  );
  al_mux2h _4470_ (
    .a(\DFF_1122.Q ),
    .b(_0415_),
    .s(\DFF_1506.Q ),
    .y(\DFF_1122.D )
  );
  al_oa21ftf _4471_ (
    .a(_0071_),
    .b(_0309_),
    .c(_0062_),
    .y(_0416_)
  );
  al_aoi21ftf _4472_ (
    .a(_0071_),
    .b(_0309_),
    .c(_0416_),
    .y(\DFF_1162.D )
  );
  al_and3 _4473_ (
    .a(\DFF_1286.Q ),
    .b(\DFF_1429.Q ),
    .c(_0393_),
    .y(_0417_)
  );
  al_ao21ttf _4474_ (
    .a(\DFF_1302.Q ),
    .b(\DFF_1429.Q ),
    .c(\DFF_1286.Q ),
    .y(_0418_)
  );
  al_aoi21ftt _4475_ (
    .a(_0346_),
    .b(_0418_),
    .c(_0417_),
    .y(\DFF_1286.D )
  );
  al_mux2h _4476_ (
    .a(\DFF_1367.Q ),
    .b(\DFF_1503.D ),
    .s(g3229),
    .y(\DFF_1502.D )
  );
  al_and2 _4477_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_1418.Q ),
    .y(_0419_)
  );
  al_and2 _4478_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_1416.Q ),
    .y(_0420_)
  );
  al_and2 _4479_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_1420.Q ),
    .y(_0421_)
  );
  al_or3 _4480_ (
    .a(_0419_),
    .b(_0420_),
    .c(_0421_),
    .y(_0422_)
  );
  al_nand2 _4481_ (
    .a(\DFF_1414.Q ),
    .b(\DFF_160.Q ),
    .y(_0423_)
  );
  al_nand2 _4482_ (
    .a(\DFF_1467.Q ),
    .b(\DFF_1504.Q ),
    .y(_0424_)
  );
  al_aoi21ttf _4483_ (
    .a(\DFF_1469.Q ),
    .b(\DFF_1506.Q ),
    .c(_0424_),
    .y(_0425_)
  );
  al_aoi21ftf _4484_ (
    .a(_0353_),
    .b(\DFF_1468.Q ),
    .c(_0425_),
    .y(_0426_)
  );
  al_ao21ftf _4485_ (
    .a(_0423_),
    .b(_0422_),
    .c(_0426_),
    .y(_0427_)
  );
  al_and2ft _4486_ (
    .a(_0008_),
    .b(_0427_),
    .y(_0428_)
  );
  al_mux2h _4487_ (
    .a(\DFF_1467.Q ),
    .b(_0428_),
    .s(\DFF_1504.Q ),
    .y(\DFF_1467.D )
  );
  al_mux2h _4488_ (
    .a(\DFF_1468.Q ),
    .b(_0428_),
    .s(\DFF_1505.Q ),
    .y(\DFF_1468.D )
  );
  al_mux2h _4489_ (
    .a(\DFF_1469.Q ),
    .b(_0428_),
    .s(\DFF_1506.Q ),
    .y(\DFF_1469.D )
  );
  al_and2 _4490_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_1424.Q ),
    .y(_0429_)
  );
  al_and2 _4491_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_1422.Q ),
    .y(_0430_)
  );
  al_and2 _4492_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_1426.Q ),
    .y(_0431_)
  );
  al_or3 _4493_ (
    .a(_0429_),
    .b(_0430_),
    .c(_0431_),
    .y(_0432_)
  );
  al_nand2 _4494_ (
    .a(\DFF_1447.Q ),
    .b(\DFF_160.Q ),
    .y(_0433_)
  );
  al_nand2 _4495_ (
    .a(\DFF_1470.Q ),
    .b(\DFF_1504.Q ),
    .y(_0434_)
  );
  al_aoi21ttf _4496_ (
    .a(\DFF_1472.Q ),
    .b(\DFF_1506.Q ),
    .c(_0434_),
    .y(_0435_)
  );
  al_aoi21ftf _4497_ (
    .a(_0353_),
    .b(\DFF_1471.Q ),
    .c(_0435_),
    .y(_0436_)
  );
  al_ao21ftf _4498_ (
    .a(_0433_),
    .b(_0432_),
    .c(_0436_),
    .y(_0437_)
  );
  al_and2ft _4499_ (
    .a(_0008_),
    .b(_0437_),
    .y(_0438_)
  );
  al_mux2h _4500_ (
    .a(\DFF_1470.Q ),
    .b(_0438_),
    .s(\DFF_1504.Q ),
    .y(\DFF_1470.D )
  );
  al_mux2h _4501_ (
    .a(\DFF_1471.Q ),
    .b(_0438_),
    .s(\DFF_1505.Q ),
    .y(\DFF_1471.D )
  );
  al_mux2h _4502_ (
    .a(\DFF_1472.Q ),
    .b(_0438_),
    .s(\DFF_1506.Q ),
    .y(\DFF_1472.D )
  );
  al_oa21ftf _4503_ (
    .a(_0097_),
    .b(_0324_),
    .c(_0088_),
    .y(_0439_)
  );
  al_aoi21ftf _4504_ (
    .a(_0097_),
    .b(_0324_),
    .c(_0439_),
    .y(\DFF_1512.D )
  );
  al_nand3 _4505_ (
    .a(\DFF_6.Q ),
    .b(\DFF_7.Q ),
    .c(_0263_),
    .y(_0440_)
  );
  al_ao21 _4506_ (
    .a(\DFF_6.Q ),
    .b(_0263_),
    .c(\DFF_7.Q ),
    .y(_0441_)
  );
  al_and3 _4507_ (
    .a(_0440_),
    .b(_0441_),
    .c(_0261_),
    .y(\DFF_7.D )
  );
  al_or2 _4508_ (
    .a(\DFF_13.Q ),
    .b(_0330_),
    .y(_0442_)
  );
  al_and2 _4509_ (
    .a(\DFF_13.Q ),
    .b(_0330_),
    .y(_0443_)
  );
  al_and3ftt _4510_ (
    .a(_0443_),
    .b(_0442_),
    .c(_0329_),
    .y(\DFF_13.D )
  );
  al_and3 _4511_ (
    .a(\DFF_1602.Q ),
    .b(\DFF_1603.Q ),
    .c(_0340_),
    .y(_0444_)
  );
  al_ao21 _4512_ (
    .a(\DFF_1602.Q ),
    .b(_0340_),
    .c(\DFF_1603.Q ),
    .y(_0445_)
  );
  al_and3ftt _4513_ (
    .a(_0444_),
    .b(_0445_),
    .c(_0339_),
    .y(\DFF_1603.D )
  );
  al_ao21 _4514_ (
    .a(\DFF_1608.Q ),
    .b(_0334_),
    .c(\DFF_1609.Q ),
    .y(_0446_)
  );
  al_and3 _4515_ (
    .a(\DFF_1609.Q ),
    .b(\DFF_1608.Q ),
    .c(_0334_),
    .y(_0447_)
  );
  al_and3ftt _4516_ (
    .a(_0447_),
    .b(_0446_),
    .c(_0336_),
    .y(\DFF_1609.D )
  );
  al_and3 _4517_ (
    .a(\DFF_236.Q ),
    .b(\DFF_237.Q ),
    .c(_0346_),
    .y(_0448_)
  );
  al_and3ftt _4518_ (
    .a(_0345_),
    .b(_0158_),
    .c(_0256_),
    .y(_0449_)
  );
  al_ao21 _4519_ (
    .a(\DFF_236.Q ),
    .b(_0346_),
    .c(\DFF_237.Q ),
    .y(_0450_)
  );
  al_and3fft _4520_ (
    .a(_0449_),
    .b(_0448_),
    .c(_0450_),
    .y(\DFF_237.D )
  );
  al_nor2 _4521_ (
    .a(\DFF_11.Q ),
    .b(\DFF_12.Q ),
    .y(_0451_)
  );
  al_and2ft _4522_ (
    .a(\DFF_14.Q ),
    .b(\DFF_4.Q ),
    .y(_0452_)
  );
  al_nand3ftt _4523_ (
    .a(\DFF_5.Q ),
    .b(\DFF_13.Q ),
    .c(_0452_),
    .y(_0453_)
  );
  al_nor3ftt _4524_ (
    .a(_0451_),
    .b(_0453_),
    .c(_0393_),
    .y(\DFF_1296.D )
  );
  al_nand2 _4525_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_1296.D ),
    .y(_0454_)
  );
  al_and2 _4526_ (
    .a(\DFF_72.Q ),
    .b(\DFF_66.Q ),
    .y(_0455_)
  );
  al_and3ftt _4527_ (
    .a(\DFF_70.Q ),
    .b(\DFF_300.D ),
    .c(_0455_),
    .y(_0456_)
  );
  al_mux2l _4528_ (
    .a(\DFF_194.Q ),
    .b(_0456_),
    .s(_0454_),
    .y(\DFF_194.D )
  );
  al_nand2 _4529_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_1296.D ),
    .y(_0457_)
  );
  al_mux2l _4530_ (
    .a(\DFF_195.Q ),
    .b(_0456_),
    .s(_0457_),
    .y(\DFF_195.D )
  );
  al_nand2 _4531_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_1296.D ),
    .y(_0458_)
  );
  al_mux2l _4532_ (
    .a(\DFF_196.Q ),
    .b(_0456_),
    .s(_0458_),
    .y(\DFF_196.D )
  );
  al_mux2l _4533_ (
    .a(\DFF_197.Q ),
    .b(\DFF_310.D ),
    .s(_0454_),
    .y(\DFF_197.D )
  );
  al_mux2l _4534_ (
    .a(\DFF_198.Q ),
    .b(\DFF_310.D ),
    .s(_0457_),
    .y(\DFF_198.D )
  );
  al_mux2l _4535_ (
    .a(\DFF_199.Q ),
    .b(\DFF_310.D ),
    .s(_0458_),
    .y(\DFF_199.D )
  );
  al_mux2l _4536_ (
    .a(\DFF_200.Q ),
    .b(\DFF_312.D ),
    .s(_0454_),
    .y(\DFF_200.D )
  );
  al_mux2l _4537_ (
    .a(\DFF_201.Q ),
    .b(\DFF_312.D ),
    .s(_0457_),
    .y(\DFF_201.D )
  );
  al_mux2l _4538_ (
    .a(\DFF_202.Q ),
    .b(\DFF_312.D ),
    .s(_0458_),
    .y(\DFF_202.D )
  );
  al_nand2 _4539_ (
    .a(\DFF_80.Q ),
    .b(\DFF_68.Q ),
    .y(_0459_)
  );
  al_nand2 _4540_ (
    .a(\DFF_78.Q ),
    .b(\DFF_70.Q ),
    .y(_0460_)
  );
  al_and3 _4541_ (
    .a(\DFF_74.Q ),
    .b(\DFF_76.Q ),
    .c(_0455_),
    .y(_0461_)
  );
  al_nand3fft _4542_ (
    .a(_0459_),
    .b(_0460_),
    .c(_0461_),
    .y(_0462_)
  );
  al_mux2l _4543_ (
    .a(\DFF_203.Q ),
    .b(_0462_),
    .s(_0454_),
    .y(\DFF_203.D )
  );
  al_mux2l _4544_ (
    .a(\DFF_204.Q ),
    .b(_0462_),
    .s(_0457_),
    .y(\DFF_204.D )
  );
  al_mux2l _4545_ (
    .a(\DFF_205.Q ),
    .b(_0462_),
    .s(_0458_),
    .y(\DFF_205.D )
  );
  al_inv _4546_ (
    .a(_0029_),
    .y(_0463_)
  );
  al_and3 _4547_ (
    .a(\DFF_462.Q ),
    .b(\DFF_463.Q ),
    .c(_0277_),
    .y(_0464_)
  );
  al_aoi21 _4548_ (
    .a(\DFF_462.Q ),
    .b(_0277_),
    .c(\DFF_463.Q ),
    .y(_0465_)
  );
  al_nor3ftt _4549_ (
    .a(_0463_),
    .b(_0464_),
    .c(_0465_),
    .y(\DFF_463.D )
  );
  al_nand2ft _4550_ (
    .a(\DFF_491.Q ),
    .b(\DFF_1505.Q ),
    .y(_0466_)
  );
  al_aoi21ftf _4551_ (
    .a(\DFF_492.Q ),
    .b(\DFF_1506.Q ),
    .c(_0466_),
    .y(_0467_)
  );
  al_aoi21ftf _4552_ (
    .a(\DFF_490.Q ),
    .b(\DFF_1504.Q ),
    .c(_0467_),
    .y(_0468_)
  );
  al_and2 _4553_ (
    .a(_0021_),
    .b(_0468_),
    .y(_0469_)
  );
  al_or2 _4554_ (
    .a(_0021_),
    .b(_0468_),
    .y(_0470_)
  );
  al_nand2ft _4555_ (
    .a(_0469_),
    .b(_0470_),
    .y(_0471_)
  );
  al_nand2ft _4556_ (
    .a(\DFF_485.Q ),
    .b(\DFF_1505.Q ),
    .y(_0472_)
  );
  al_aoi21ftf _4557_ (
    .a(\DFF_486.Q ),
    .b(\DFF_1506.Q ),
    .c(_0472_),
    .y(_0473_)
  );
  al_ao21ftf _4558_ (
    .a(\DFF_484.Q ),
    .b(\DFF_1504.Q ),
    .c(_0473_),
    .y(_0474_)
  );
  al_nand2 _4559_ (
    .a(_0019_),
    .b(_0474_),
    .y(_0475_)
  );
  al_or2 _4560_ (
    .a(_0019_),
    .b(_0474_),
    .y(_0476_)
  );
  al_and3 _4561_ (
    .a(_0475_),
    .b(_0476_),
    .c(_0471_),
    .y(_0477_)
  );
  al_nand2ft _4562_ (
    .a(\DFF_477.Q ),
    .b(\DFF_1506.Q ),
    .y(_0478_)
  );
  al_aoi21ftf _4563_ (
    .a(\DFF_475.Q ),
    .b(\DFF_1504.Q ),
    .c(_0478_),
    .y(_0479_)
  );
  al_ao21ftf _4564_ (
    .a(\DFF_476.Q ),
    .b(\DFF_1505.Q ),
    .c(_0479_),
    .y(_0480_)
  );
  al_nand2 _4565_ (
    .a(_0016_),
    .b(_0480_),
    .y(_0481_)
  );
  al_nand2ft _4566_ (
    .a(\DFF_470.Q ),
    .b(\DFF_1505.Q ),
    .y(_0482_)
  );
  al_aoi21ftf _4567_ (
    .a(\DFF_471.Q ),
    .b(\DFF_1506.Q ),
    .c(_0482_),
    .y(_0483_)
  );
  al_ao21ftf _4568_ (
    .a(\DFF_469.Q ),
    .b(\DFF_1504.Q ),
    .c(_0483_),
    .y(_0484_)
  );
  al_aoi21ftf _4569_ (
    .a(_0484_),
    .b(\DFF_459.Q ),
    .c(_0481_),
    .y(_0485_)
  );
  al_nand2 _4570_ (
    .a(_0010_),
    .b(_0484_),
    .y(_0486_)
  );
  al_nand2ft _4571_ (
    .a(\DFF_494.Q ),
    .b(\DFF_1505.Q ),
    .y(_0487_)
  );
  al_aoi21ftf _4572_ (
    .a(\DFF_495.Q ),
    .b(\DFF_1506.Q ),
    .c(_0487_),
    .y(_0488_)
  );
  al_ao21ftf _4573_ (
    .a(\DFF_493.Q ),
    .b(\DFF_1504.Q ),
    .c(_0488_),
    .y(_0489_)
  );
  al_aoi21ftf _4574_ (
    .a(\DFF_467.Q ),
    .b(_0489_),
    .c(_0486_),
    .y(_0490_)
  );
  al_and3 _4575_ (
    .a(_0485_),
    .b(_0490_),
    .c(_0477_),
    .y(_0491_)
  );
  al_nand2ft _4576_ (
    .a(\DFF_479.Q ),
    .b(\DFF_1505.Q ),
    .y(_0492_)
  );
  al_aoi21ftf _4577_ (
    .a(\DFF_480.Q ),
    .b(\DFF_1506.Q ),
    .c(_0492_),
    .y(_0493_)
  );
  al_ao21ftf _4578_ (
    .a(\DFF_478.Q ),
    .b(\DFF_1504.Q ),
    .c(_0493_),
    .y(_0494_)
  );
  al_or2 _4579_ (
    .a(\DFF_462.Q ),
    .b(_0494_),
    .y(_0495_)
  );
  al_and2 _4580_ (
    .a(\DFF_462.Q ),
    .b(_0494_),
    .y(_0496_)
  );
  al_nand2ft _4581_ (
    .a(_0496_),
    .b(_0495_),
    .y(_0497_)
  );
  al_nand2ft _4582_ (
    .a(\DFF_473.Q ),
    .b(\DFF_1505.Q ),
    .y(_0498_)
  );
  al_aoi21ftf _4583_ (
    .a(\DFF_474.Q ),
    .b(\DFF_1506.Q ),
    .c(_0498_),
    .y(_0499_)
  );
  al_ao21ftf _4584_ (
    .a(\DFF_472.Q ),
    .b(\DFF_1504.Q ),
    .c(_0499_),
    .y(_0500_)
  );
  al_nand2 _4585_ (
    .a(_0014_),
    .b(_0500_),
    .y(_0501_)
  );
  al_or2 _4586_ (
    .a(_0014_),
    .b(_0500_),
    .y(_0502_)
  );
  al_and3 _4587_ (
    .a(_0501_),
    .b(_0502_),
    .c(_0497_),
    .y(_0503_)
  );
  al_nand2ft _4588_ (
    .a(\DFF_497.Q ),
    .b(\DFF_1505.Q ),
    .y(_0504_)
  );
  al_aoi21ftf _4589_ (
    .a(\DFF_498.Q ),
    .b(\DFF_1506.Q ),
    .c(_0504_),
    .y(_0505_)
  );
  al_ao21ftf _4590_ (
    .a(\DFF_496.Q ),
    .b(\DFF_1504.Q ),
    .c(_0505_),
    .y(_0506_)
  );
  al_nand2 _4591_ (
    .a(_0023_),
    .b(_0506_),
    .y(_0507_)
  );
  al_or2 _4592_ (
    .a(_0023_),
    .b(_0506_),
    .y(_0508_)
  );
  al_nand2ft _4593_ (
    .a(\DFF_482.Q ),
    .b(\DFF_1505.Q ),
    .y(_0509_)
  );
  al_aoi21ftf _4594_ (
    .a(\DFF_483.Q ),
    .b(\DFF_1506.Q ),
    .c(_0509_),
    .y(_0510_)
  );
  al_aoi21ftf _4595_ (
    .a(\DFF_481.Q ),
    .b(\DFF_1504.Q ),
    .c(_0510_),
    .y(_0511_)
  );
  al_nand2 _4596_ (
    .a(\DFF_463.Q ),
    .b(_0511_),
    .y(_0512_)
  );
  al_aoi21ftf _4597_ (
    .a(_0480_),
    .b(\DFF_461.Q ),
    .c(_0512_),
    .y(_0513_)
  );
  al_and3 _4598_ (
    .a(_0507_),
    .b(_0508_),
    .c(_0513_),
    .y(_0514_)
  );
  al_nand2ft _4599_ (
    .a(\DFF_488.Q ),
    .b(\DFF_1505.Q ),
    .y(_0515_)
  );
  al_aoi21ftf _4600_ (
    .a(\DFF_489.Q ),
    .b(\DFF_1506.Q ),
    .c(_0515_),
    .y(_0516_)
  );
  al_ao21ftf _4601_ (
    .a(\DFF_487.Q ),
    .b(\DFF_1504.Q ),
    .c(_0516_),
    .y(_0517_)
  );
  al_and2 _4602_ (
    .a(_0020_),
    .b(_0517_),
    .y(_0518_)
  );
  al_nor2 _4603_ (
    .a(_0020_),
    .b(_0517_),
    .y(_0519_)
  );
  al_ao21ftf _4604_ (
    .a(\DFF_481.Q ),
    .b(\DFF_1504.Q ),
    .c(_0510_),
    .y(_0520_)
  );
  al_nand2 _4605_ (
    .a(_0018_),
    .b(_0520_),
    .y(_0521_)
  );
  al_aoi21ftf _4606_ (
    .a(_0489_),
    .b(\DFF_467.Q ),
    .c(_0521_),
    .y(_0522_)
  );
  al_nand3fft _4607_ (
    .a(_0518_),
    .b(_0519_),
    .c(_0522_),
    .y(_0523_)
  );
  al_and3ftt _4608_ (
    .a(_0523_),
    .b(_0514_),
    .c(_0503_),
    .y(_0524_)
  );
  al_nand2ft _4609_ (
    .a(\DFF_502.Q ),
    .b(\DFF_1504.Q ),
    .y(_0525_)
  );
  al_aoi21ftf _4610_ (
    .a(\DFF_504.Q ),
    .b(\DFF_1506.Q ),
    .c(_0525_),
    .y(_0526_)
  );
  al_aoi21ftf _4611_ (
    .a(\DFF_503.Q ),
    .b(\DFF_1505.Q ),
    .c(_0526_),
    .y(_0527_)
  );
  al_nand2ft _4612_ (
    .a(\DFF_500.Q ),
    .b(\DFF_1505.Q ),
    .y(_0528_)
  );
  al_nand2ft _4613_ (
    .a(\DFF_499.Q ),
    .b(\DFF_1504.Q ),
    .y(_0529_)
  );
  al_aoi21ftf _4614_ (
    .a(\DFF_501.Q ),
    .b(\DFF_1506.Q ),
    .c(_0529_),
    .y(_0530_)
  );
  al_nand3 _4615_ (
    .a(_0528_),
    .b(_0530_),
    .c(_0527_),
    .y(_0531_)
  );
  al_aoi21 _4616_ (
    .a(_0524_),
    .b(_0491_),
    .c(_0531_),
    .y(_0532_)
  );
  al_mux2l _4617_ (
    .a(\DFF_505.Q ),
    .b(_0532_),
    .s(_0015_),
    .y(\DFF_505.D )
  );
  al_mux2l _4618_ (
    .a(\DFF_506.Q ),
    .b(_0532_),
    .s(_0012_),
    .y(\DFF_506.D )
  );
  al_mux2l _4619_ (
    .a(\DFF_507.Q ),
    .b(_0532_),
    .s(_0013_),
    .y(\DFF_507.D )
  );
  al_and3 _4620_ (
    .a(\DFF_586.Q ),
    .b(\DFF_587.Q ),
    .c(_0346_),
    .y(_0533_)
  );
  al_ao21 _4621_ (
    .a(\DFF_586.Q ),
    .b(_0346_),
    .c(\DFF_587.Q ),
    .y(_0534_)
  );
  al_and3fft _4622_ (
    .a(_0449_),
    .b(_0533_),
    .c(_0534_),
    .y(\DFF_587.D )
  );
  al_and2 _4623_ (
    .a(\DFF_54.Q ),
    .b(\DFF_48.Q ),
    .y(_0535_)
  );
  al_and3ftt _4624_ (
    .a(\DFF_52.Q ),
    .b(\DFF_650.D ),
    .c(_0535_),
    .y(_0536_)
  );
  al_mux2l _4625_ (
    .a(\DFF_544.Q ),
    .b(_0536_),
    .s(_0454_),
    .y(\DFF_544.D )
  );
  al_mux2l _4626_ (
    .a(\DFF_545.Q ),
    .b(_0536_),
    .s(_0457_),
    .y(\DFF_545.D )
  );
  al_mux2l _4627_ (
    .a(\DFF_546.Q ),
    .b(_0536_),
    .s(_0458_),
    .y(\DFF_546.D )
  );
  al_mux2l _4628_ (
    .a(\DFF_547.Q ),
    .b(\DFF_660.D ),
    .s(_0454_),
    .y(\DFF_547.D )
  );
  al_mux2l _4629_ (
    .a(\DFF_548.Q ),
    .b(\DFF_660.D ),
    .s(_0457_),
    .y(\DFF_548.D )
  );
  al_mux2l _4630_ (
    .a(\DFF_549.Q ),
    .b(\DFF_660.D ),
    .s(_0458_),
    .y(\DFF_549.D )
  );
  al_mux2l _4631_ (
    .a(\DFF_550.Q ),
    .b(\DFF_662.D ),
    .s(_0454_),
    .y(\DFF_550.D )
  );
  al_mux2l _4632_ (
    .a(\DFF_551.Q ),
    .b(\DFF_662.D ),
    .s(_0457_),
    .y(\DFF_551.D )
  );
  al_mux2l _4633_ (
    .a(\DFF_552.Q ),
    .b(\DFF_662.D ),
    .s(_0458_),
    .y(\DFF_552.D )
  );
  al_and2 _4634_ (
    .a(\DFF_60.Q ),
    .b(\DFF_62.Q ),
    .y(_0537_)
  );
  al_nand3 _4635_ (
    .a(\DFF_50.Q ),
    .b(\DFF_52.Q ),
    .c(_0537_),
    .y(_0538_)
  );
  al_nand3 _4636_ (
    .a(\DFF_56.Q ),
    .b(\DFF_58.Q ),
    .c(_0535_),
    .y(_0539_)
  );
  al_or2 _4637_ (
    .a(_0538_),
    .b(_0539_),
    .y(_0540_)
  );
  al_mux2l _4638_ (
    .a(\DFF_553.Q ),
    .b(_0540_),
    .s(_0454_),
    .y(\DFF_553.D )
  );
  al_mux2l _4639_ (
    .a(\DFF_554.Q ),
    .b(_0540_),
    .s(_0457_),
    .y(\DFF_554.D )
  );
  al_mux2l _4640_ (
    .a(\DFF_555.Q ),
    .b(_0540_),
    .s(_0458_),
    .y(\DFF_555.D )
  );
  al_inv _4641_ (
    .a(_0035_),
    .y(_0541_)
  );
  al_and3 _4642_ (
    .a(\DFF_812.Q ),
    .b(\DFF_813.Q ),
    .c(_0293_),
    .y(_0542_)
  );
  al_aoi21 _4643_ (
    .a(\DFF_812.Q ),
    .b(_0293_),
    .c(\DFF_813.Q ),
    .y(_0543_)
  );
  al_nor3ftt _4644_ (
    .a(_0541_),
    .b(_0542_),
    .c(_0543_),
    .y(\DFF_813.D )
  );
  al_nand2ft _4645_ (
    .a(\DFF_838.Q ),
    .b(\DFF_1505.Q ),
    .y(_0544_)
  );
  al_aoi21ftf _4646_ (
    .a(\DFF_839.Q ),
    .b(\DFF_1506.Q ),
    .c(_0544_),
    .y(_0545_)
  );
  al_ao21ftf _4647_ (
    .a(\DFF_837.Q ),
    .b(\DFF_1504.Q ),
    .c(_0545_),
    .y(_0546_)
  );
  al_and2 _4648_ (
    .a(\DFF_815.Q ),
    .b(_0546_),
    .y(_0547_)
  );
  al_or2 _4649_ (
    .a(\DFF_815.Q ),
    .b(_0546_),
    .y(_0548_)
  );
  al_nand2ft _4650_ (
    .a(_0547_),
    .b(_0548_),
    .y(_0549_)
  );
  al_nand2ft _4651_ (
    .a(\DFF_832.Q ),
    .b(\DFF_1505.Q ),
    .y(_0550_)
  );
  al_aoi21ftf _4652_ (
    .a(\DFF_833.Q ),
    .b(\DFF_1506.Q ),
    .c(_0550_),
    .y(_0551_)
  );
  al_ao21ftf _4653_ (
    .a(\DFF_831.Q ),
    .b(\DFF_1504.Q ),
    .c(_0551_),
    .y(_0552_)
  );
  al_nand2 _4654_ (
    .a(_0045_),
    .b(_0552_),
    .y(_0553_)
  );
  al_or2 _4655_ (
    .a(_0045_),
    .b(_0552_),
    .y(_0554_)
  );
  al_nand2ft _4656_ (
    .a(\DFF_829.Q ),
    .b(\DFF_1505.Q ),
    .y(_0555_)
  );
  al_aoi21ftf _4657_ (
    .a(\DFF_830.Q ),
    .b(\DFF_1506.Q ),
    .c(_0555_),
    .y(_0556_)
  );
  al_ao21ftf _4658_ (
    .a(\DFF_828.Q ),
    .b(\DFF_1504.Q ),
    .c(_0556_),
    .y(_0557_)
  );
  al_and2 _4659_ (
    .a(\DFF_812.Q ),
    .b(_0557_),
    .y(_0558_)
  );
  al_or2 _4660_ (
    .a(\DFF_812.Q ),
    .b(_0557_),
    .y(_0559_)
  );
  al_nand2ft _4661_ (
    .a(_0558_),
    .b(_0559_),
    .y(_0560_)
  );
  al_and3 _4662_ (
    .a(_0553_),
    .b(_0554_),
    .c(_0560_),
    .y(_0561_)
  );
  al_nand2ft _4663_ (
    .a(\DFF_847.Q ),
    .b(\DFF_1505.Q ),
    .y(_0562_)
  );
  al_aoi21ftf _4664_ (
    .a(\DFF_848.Q ),
    .b(\DFF_1506.Q ),
    .c(_0562_),
    .y(_0563_)
  );
  al_aoi21ftf _4665_ (
    .a(\DFF_846.Q ),
    .b(\DFF_1504.Q ),
    .c(_0563_),
    .y(_0564_)
  );
  al_nand2 _4666_ (
    .a(\DFF_818.Q ),
    .b(_0564_),
    .y(_0565_)
  );
  al_or2 _4667_ (
    .a(\DFF_818.Q ),
    .b(_0564_),
    .y(_0566_)
  );
  al_nand2ft _4668_ (
    .a(\DFF_835.Q ),
    .b(\DFF_1505.Q ),
    .y(_0567_)
  );
  al_aoi21ftf _4669_ (
    .a(\DFF_836.Q ),
    .b(\DFF_1506.Q ),
    .c(_0567_),
    .y(_0568_)
  );
  al_ao21ftf _4670_ (
    .a(\DFF_834.Q ),
    .b(\DFF_1504.Q ),
    .c(_0568_),
    .y(_0569_)
  );
  al_nand2 _4671_ (
    .a(_0046_),
    .b(_0569_),
    .y(_0570_)
  );
  al_nand2ft _4672_ (
    .a(\DFF_826.Q ),
    .b(\DFF_1505.Q ),
    .y(_0571_)
  );
  al_aoi21ftf _4673_ (
    .a(\DFF_827.Q ),
    .b(\DFF_1506.Q ),
    .c(_0571_),
    .y(_0572_)
  );
  al_ao21ftf _4674_ (
    .a(\DFF_825.Q ),
    .b(\DFF_1504.Q ),
    .c(_0572_),
    .y(_0573_)
  );
  al_aoi21ftf _4675_ (
    .a(_0573_),
    .b(\DFF_811.Q ),
    .c(_0570_),
    .y(_0574_)
  );
  al_and3 _4676_ (
    .a(_0565_),
    .b(_0566_),
    .c(_0574_),
    .y(_0575_)
  );
  al_and3 _4677_ (
    .a(_0549_),
    .b(_0575_),
    .c(_0561_),
    .y(_0576_)
  );
  al_nand2ft _4678_ (
    .a(\DFF_841.Q ),
    .b(\DFF_1505.Q ),
    .y(_0577_)
  );
  al_aoi21ftf _4679_ (
    .a(\DFF_842.Q ),
    .b(\DFF_1506.Q ),
    .c(_0577_),
    .y(_0578_)
  );
  al_ao21ftf _4680_ (
    .a(\DFF_840.Q ),
    .b(\DFF_1504.Q ),
    .c(_0578_),
    .y(_0579_)
  );
  al_and2 _4681_ (
    .a(\DFF_816.Q ),
    .b(_0579_),
    .y(_0580_)
  );
  al_or2 _4682_ (
    .a(\DFF_816.Q ),
    .b(_0579_),
    .y(_0581_)
  );
  al_nand2ft _4683_ (
    .a(_0580_),
    .b(_0581_),
    .y(_0582_)
  );
  al_nand2ft _4684_ (
    .a(\DFF_844.Q ),
    .b(\DFF_1505.Q ),
    .y(_0583_)
  );
  al_aoi21ftf _4685_ (
    .a(\DFF_845.Q ),
    .b(\DFF_1506.Q ),
    .c(_0583_),
    .y(_0584_)
  );
  al_ao21ftf _4686_ (
    .a(\DFF_843.Q ),
    .b(\DFF_1504.Q ),
    .c(_0584_),
    .y(_0585_)
  );
  al_and2 _4687_ (
    .a(_0049_),
    .b(_0585_),
    .y(_0586_)
  );
  al_nor2 _4688_ (
    .a(_0049_),
    .b(_0585_),
    .y(_0587_)
  );
  al_nand2ft _4689_ (
    .a(\DFF_820.Q ),
    .b(\DFF_1505.Q ),
    .y(_0588_)
  );
  al_aoi21ftf _4690_ (
    .a(\DFF_821.Q ),
    .b(\DFF_1506.Q ),
    .c(_0588_),
    .y(_0589_)
  );
  al_ao21ftf _4691_ (
    .a(\DFF_819.Q ),
    .b(\DFF_1504.Q ),
    .c(_0589_),
    .y(_0590_)
  );
  al_nand2 _4692_ (
    .a(_0037_),
    .b(_0590_),
    .y(_0591_)
  );
  al_aoi21ftf _4693_ (
    .a(_0569_),
    .b(\DFF_814.Q ),
    .c(_0591_),
    .y(_0592_)
  );
  al_nand3fft _4694_ (
    .a(_0586_),
    .b(_0587_),
    .c(_0592_),
    .y(_0593_)
  );
  al_nand2ft _4695_ (
    .a(\DFF_823.Q ),
    .b(\DFF_1505.Q ),
    .y(_0594_)
  );
  al_aoi21ftf _4696_ (
    .a(\DFF_824.Q ),
    .b(\DFF_1506.Q ),
    .c(_0594_),
    .y(_0595_)
  );
  al_ao21ftf _4697_ (
    .a(\DFF_822.Q ),
    .b(\DFF_1504.Q ),
    .c(_0595_),
    .y(_0596_)
  );
  al_nor2 _4698_ (
    .a(_0042_),
    .b(_0596_),
    .y(_0597_)
  );
  al_and2 _4699_ (
    .a(_0042_),
    .b(_0596_),
    .y(_0598_)
  );
  al_nand2 _4700_ (
    .a(_0043_),
    .b(_0573_),
    .y(_0599_)
  );
  al_aoi21ftf _4701_ (
    .a(_0590_),
    .b(\DFF_809.Q ),
    .c(_0599_),
    .y(_0600_)
  );
  al_nand3fft _4702_ (
    .a(_0597_),
    .b(_0598_),
    .c(_0600_),
    .y(_0601_)
  );
  al_nor3ftt _4703_ (
    .a(_0582_),
    .b(_0593_),
    .c(_0601_),
    .y(_0602_)
  );
  al_nand2ft _4704_ (
    .a(\DFF_853.Q ),
    .b(\DFF_1505.Q ),
    .y(_0603_)
  );
  al_aoi21ftf _4705_ (
    .a(\DFF_854.Q ),
    .b(\DFF_1506.Q ),
    .c(_0603_),
    .y(_0604_)
  );
  al_aoi21ftf _4706_ (
    .a(\DFF_852.Q ),
    .b(\DFF_1504.Q ),
    .c(_0604_),
    .y(_0605_)
  );
  al_nand2ft _4707_ (
    .a(\DFF_850.Q ),
    .b(\DFF_1505.Q ),
    .y(_0606_)
  );
  al_nand2ft _4708_ (
    .a(\DFF_849.Q ),
    .b(\DFF_1504.Q ),
    .y(_0607_)
  );
  al_aoi21ftf _4709_ (
    .a(\DFF_851.Q ),
    .b(\DFF_1506.Q ),
    .c(_0607_),
    .y(_0608_)
  );
  al_nand3 _4710_ (
    .a(_0606_),
    .b(_0608_),
    .c(_0605_),
    .y(_0609_)
  );
  al_aoi21 _4711_ (
    .a(_0602_),
    .b(_0576_),
    .c(_0609_),
    .y(_0610_)
  );
  al_mux2l _4712_ (
    .a(\DFF_855.Q ),
    .b(_0610_),
    .s(_0039_),
    .y(\DFF_855.D )
  );
  al_mux2l _4713_ (
    .a(\DFF_856.Q ),
    .b(_0610_),
    .s(_0040_),
    .y(\DFF_856.D )
  );
  al_mux2l _4714_ (
    .a(\DFF_857.Q ),
    .b(_0610_),
    .s(_0041_),
    .y(\DFF_857.D )
  );
  al_and3 _4715_ (
    .a(\DFF_936.Q ),
    .b(\DFF_937.Q ),
    .c(_0346_),
    .y(_0611_)
  );
  al_ao21 _4716_ (
    .a(\DFF_936.Q ),
    .b(_0346_),
    .c(\DFF_937.Q ),
    .y(_0612_)
  );
  al_and3fft _4717_ (
    .a(_0449_),
    .b(_0611_),
    .c(_0612_),
    .y(\DFF_937.D )
  );
  al_and2 _4718_ (
    .a(\DFF_41.Q ),
    .b(\DFF_38.Q ),
    .y(_0613_)
  );
  al_and3ftt _4719_ (
    .a(\DFF_40.Q ),
    .b(\DFF_1000.D ),
    .c(_0613_),
    .y(_0614_)
  );
  al_mux2l _4720_ (
    .a(\DFF_894.Q ),
    .b(_0614_),
    .s(_0454_),
    .y(\DFF_894.D )
  );
  al_mux2l _4721_ (
    .a(\DFF_895.Q ),
    .b(_0614_),
    .s(_0457_),
    .y(\DFF_895.D )
  );
  al_mux2l _4722_ (
    .a(\DFF_896.Q ),
    .b(_0614_),
    .s(_0458_),
    .y(\DFF_896.D )
  );
  al_mux2l _4723_ (
    .a(\DFF_897.Q ),
    .b(\DFF_1010.D ),
    .s(_0454_),
    .y(\DFF_897.D )
  );
  al_mux2l _4724_ (
    .a(\DFF_898.Q ),
    .b(\DFF_1010.D ),
    .s(_0457_),
    .y(\DFF_898.D )
  );
  al_mux2l _4725_ (
    .a(\DFF_899.Q ),
    .b(\DFF_1010.D ),
    .s(_0458_),
    .y(\DFF_899.D )
  );
  al_mux2l _4726_ (
    .a(\DFF_900.Q ),
    .b(\DFF_1012.D ),
    .s(_0454_),
    .y(\DFF_900.D )
  );
  al_mux2l _4727_ (
    .a(\DFF_901.Q ),
    .b(\DFF_1012.D ),
    .s(_0457_),
    .y(\DFF_901.D )
  );
  al_mux2l _4728_ (
    .a(\DFF_902.Q ),
    .b(\DFF_1012.D ),
    .s(_0458_),
    .y(\DFF_902.D )
  );
  al_and2 _4729_ (
    .a(\DFF_44.Q ),
    .b(\DFF_45.Q ),
    .y(_0615_)
  );
  al_and3 _4730_ (
    .a(\DFF_39.Q ),
    .b(\DFF_40.Q ),
    .c(_0615_),
    .y(_0616_)
  );
  al_nand3 _4731_ (
    .a(\DFF_42.Q ),
    .b(\DFF_43.Q ),
    .c(_0613_),
    .y(_0617_)
  );
  al_and2ft _4732_ (
    .a(_0617_),
    .b(_0616_),
    .y(_0618_)
  );
  al_inv _4733_ (
    .a(_0618_),
    .y(_0619_)
  );
  al_mux2l _4734_ (
    .a(\DFF_903.Q ),
    .b(_0619_),
    .s(_0454_),
    .y(\DFF_903.D )
  );
  al_mux2l _4735_ (
    .a(\DFF_904.Q ),
    .b(_0619_),
    .s(_0457_),
    .y(\DFF_904.D )
  );
  al_mux2l _4736_ (
    .a(\DFF_905.Q ),
    .b(_0619_),
    .s(_0458_),
    .y(\DFF_905.D )
  );
  al_inv _4737_ (
    .a(_0062_),
    .y(_0620_)
  );
  al_and3 _4738_ (
    .a(\DFF_1162.Q ),
    .b(\DFF_1163.Q ),
    .c(_0309_),
    .y(_0621_)
  );
  al_aoi21 _4739_ (
    .a(\DFF_1162.Q ),
    .b(_0309_),
    .c(\DFF_1163.Q ),
    .y(_0622_)
  );
  al_nor3ftt _4740_ (
    .a(_0620_),
    .b(_0621_),
    .c(_0622_),
    .y(\DFF_1163.D )
  );
  al_nand2ft _4741_ (
    .a(\DFF_1191.Q ),
    .b(\DFF_1505.Q ),
    .y(_0623_)
  );
  al_aoi21ftf _4742_ (
    .a(\DFF_1192.Q ),
    .b(\DFF_1506.Q ),
    .c(_0623_),
    .y(_0624_)
  );
  al_ao21ftf _4743_ (
    .a(\DFF_1190.Q ),
    .b(\DFF_1504.Q ),
    .c(_0624_),
    .y(_0625_)
  );
  al_and2 _4744_ (
    .a(\DFF_1166.Q ),
    .b(_0625_),
    .y(_0626_)
  );
  al_aoi21ftf _4745_ (
    .a(\DFF_1190.Q ),
    .b(\DFF_1504.Q ),
    .c(_0624_),
    .y(_0627_)
  );
  al_nand2 _4746_ (
    .a(_0075_),
    .b(_0627_),
    .y(_0628_)
  );
  al_nand2ft _4747_ (
    .a(_0626_),
    .b(_0628_),
    .y(_0629_)
  );
  al_nand2ft _4748_ (
    .a(\DFF_1185.Q ),
    .b(\DFF_1505.Q ),
    .y(_0630_)
  );
  al_aoi21ftf _4749_ (
    .a(\DFF_1186.Q ),
    .b(\DFF_1506.Q ),
    .c(_0630_),
    .y(_0631_)
  );
  al_aoi21ftf _4750_ (
    .a(\DFF_1184.Q ),
    .b(\DFF_1504.Q ),
    .c(_0631_),
    .y(_0632_)
  );
  al_or2 _4751_ (
    .a(\DFF_1164.Q ),
    .b(_0632_),
    .y(_0633_)
  );
  al_nand2 _4752_ (
    .a(\DFF_1164.Q ),
    .b(_0632_),
    .y(_0634_)
  );
  al_nand2ft _4753_ (
    .a(\DFF_1194.Q ),
    .b(\DFF_1505.Q ),
    .y(_0635_)
  );
  al_aoi21ftf _4754_ (
    .a(\DFF_1195.Q ),
    .b(\DFF_1506.Q ),
    .c(_0635_),
    .y(_0636_)
  );
  al_ao21ftf _4755_ (
    .a(\DFF_1193.Q ),
    .b(\DFF_1504.Q ),
    .c(_0636_),
    .y(_0637_)
  );
  al_and2 _4756_ (
    .a(\DFF_1167.Q ),
    .b(_0637_),
    .y(_0638_)
  );
  al_or2 _4757_ (
    .a(\DFF_1167.Q ),
    .b(_0637_),
    .y(_0639_)
  );
  al_nand2ft _4758_ (
    .a(_0638_),
    .b(_0639_),
    .y(_0640_)
  );
  al_and3 _4759_ (
    .a(_0633_),
    .b(_0634_),
    .c(_0640_),
    .y(_0641_)
  );
  al_nand2ft _4760_ (
    .a(\DFF_1188.Q ),
    .b(\DFF_1505.Q ),
    .y(_0642_)
  );
  al_aoi21ftf _4761_ (
    .a(\DFF_1189.Q ),
    .b(\DFF_1506.Q ),
    .c(_0642_),
    .y(_0643_)
  );
  al_ao21ftf _4762_ (
    .a(\DFF_1187.Q ),
    .b(\DFF_1504.Q ),
    .c(_0643_),
    .y(_0644_)
  );
  al_nand2ft _4763_ (
    .a(\DFF_1197.Q ),
    .b(\DFF_1505.Q ),
    .y(_0645_)
  );
  al_aoi21ftf _4764_ (
    .a(\DFF_1198.Q ),
    .b(\DFF_1506.Q ),
    .c(_0645_),
    .y(_0646_)
  );
  al_ao21ftf _4765_ (
    .a(\DFF_1196.Q ),
    .b(\DFF_1504.Q ),
    .c(_0646_),
    .y(_0647_)
  );
  al_nand2 _4766_ (
    .a(_0074_),
    .b(_0644_),
    .y(_0648_)
  );
  al_aoi21ftf _4767_ (
    .a(_0647_),
    .b(\DFF_1168.Q ),
    .c(_0648_),
    .y(_0649_)
  );
  al_aoi21ftf _4768_ (
    .a(_0644_),
    .b(\DFF_1165.Q ),
    .c(_0649_),
    .y(_0650_)
  );
  al_and3 _4769_ (
    .a(_0629_),
    .b(_0650_),
    .c(_0641_),
    .y(_0651_)
  );
  al_nand2ft _4770_ (
    .a(\DFF_1179.Q ),
    .b(\DFF_1505.Q ),
    .y(_0652_)
  );
  al_aoi21ftf _4771_ (
    .a(\DFF_1180.Q ),
    .b(\DFF_1506.Q ),
    .c(_0652_),
    .y(_0653_)
  );
  al_ao21ftf _4772_ (
    .a(\DFF_1178.Q ),
    .b(\DFF_1504.Q ),
    .c(_0653_),
    .y(_0654_)
  );
  al_nand2 _4773_ (
    .a(_0071_),
    .b(_0654_),
    .y(_0655_)
  );
  al_or2 _4774_ (
    .a(_0071_),
    .b(_0654_),
    .y(_0656_)
  );
  al_nand2ft _4775_ (
    .a(\DFF_1182.Q ),
    .b(\DFF_1505.Q ),
    .y(_0657_)
  );
  al_aoi21ftf _4776_ (
    .a(\DFF_1183.Q ),
    .b(\DFF_1506.Q ),
    .c(_0657_),
    .y(_0658_)
  );
  al_ao21ftf _4777_ (
    .a(\DFF_1181.Q ),
    .b(\DFF_1504.Q ),
    .c(_0658_),
    .y(_0659_)
  );
  al_nand2 _4778_ (
    .a(\DFF_1163.Q ),
    .b(_0659_),
    .y(_0660_)
  );
  al_or2 _4779_ (
    .a(\DFF_1163.Q ),
    .b(_0659_),
    .y(_0661_)
  );
  al_and2 _4780_ (
    .a(_0077_),
    .b(_0647_),
    .y(_0662_)
  );
  al_aoi21 _4781_ (
    .a(_0660_),
    .b(_0661_),
    .c(_0662_),
    .y(_0663_)
  );
  al_and3 _4782_ (
    .a(_0655_),
    .b(_0656_),
    .c(_0663_),
    .y(_0664_)
  );
  al_nand2ft _4783_ (
    .a(\DFF_1170.Q ),
    .b(\DFF_1505.Q ),
    .y(_0665_)
  );
  al_aoi21ftf _4784_ (
    .a(\DFF_1171.Q ),
    .b(\DFF_1506.Q ),
    .c(_0665_),
    .y(_0666_)
  );
  al_ao21ftf _4785_ (
    .a(\DFF_1169.Q ),
    .b(\DFF_1504.Q ),
    .c(_0666_),
    .y(_0667_)
  );
  al_nand2 _4786_ (
    .a(_0064_),
    .b(_0667_),
    .y(_0668_)
  );
  al_nand2ft _4787_ (
    .a(\DFF_1177.Q ),
    .b(\DFF_1506.Q ),
    .y(_0669_)
  );
  al_aoi21ftf _4788_ (
    .a(\DFF_1175.Q ),
    .b(\DFF_1504.Q ),
    .c(_0669_),
    .y(_0670_)
  );
  al_ao21ftf _4789_ (
    .a(\DFF_1176.Q ),
    .b(\DFF_1505.Q ),
    .c(_0670_),
    .y(_0671_)
  );
  al_and2 _4790_ (
    .a(_0070_),
    .b(_0671_),
    .y(_0672_)
  );
  al_or2 _4791_ (
    .a(_0070_),
    .b(_0671_),
    .y(_0673_)
  );
  al_and3ftt _4792_ (
    .a(_0672_),
    .b(_0668_),
    .c(_0673_),
    .y(_0674_)
  );
  al_or2 _4793_ (
    .a(_0064_),
    .b(_0667_),
    .y(_0675_)
  );
  al_nand2ft _4794_ (
    .a(\DFF_1173.Q ),
    .b(\DFF_1505.Q ),
    .y(_0676_)
  );
  al_aoi21ftf _4795_ (
    .a(\DFF_1174.Q ),
    .b(\DFF_1506.Q ),
    .c(_0676_),
    .y(_0677_)
  );
  al_ao21ftf _4796_ (
    .a(\DFF_1172.Q ),
    .b(\DFF_1504.Q ),
    .c(_0677_),
    .y(_0678_)
  );
  al_and2 _4797_ (
    .a(_0069_),
    .b(_0678_),
    .y(_0679_)
  );
  al_or2 _4798_ (
    .a(_0069_),
    .b(_0678_),
    .y(_0680_)
  );
  al_and3ftt _4799_ (
    .a(_0679_),
    .b(_0675_),
    .c(_0680_),
    .y(_0681_)
  );
  al_and3 _4800_ (
    .a(_0674_),
    .b(_0681_),
    .c(_0664_),
    .y(_0682_)
  );
  al_nand2ft _4801_ (
    .a(\DFF_1203.Q ),
    .b(\DFF_1505.Q ),
    .y(_0683_)
  );
  al_nand2ft _4802_ (
    .a(\DFF_1202.Q ),
    .b(\DFF_1504.Q ),
    .y(_0684_)
  );
  al_and2ft _4803_ (
    .a(\DFF_1204.Q ),
    .b(\DFF_1506.Q ),
    .y(_0685_)
  );
  al_and3ftt _4804_ (
    .a(_0685_),
    .b(_0683_),
    .c(_0684_),
    .y(_0686_)
  );
  al_nand2ft _4805_ (
    .a(\DFF_1200.Q ),
    .b(\DFF_1505.Q ),
    .y(_0687_)
  );
  al_nand2ft _4806_ (
    .a(\DFF_1199.Q ),
    .b(\DFF_1504.Q ),
    .y(_0688_)
  );
  al_aoi21ftf _4807_ (
    .a(\DFF_1201.Q ),
    .b(\DFF_1506.Q ),
    .c(_0688_),
    .y(_0689_)
  );
  al_nand3 _4808_ (
    .a(_0687_),
    .b(_0689_),
    .c(_0686_),
    .y(_0690_)
  );
  al_aoi21 _4809_ (
    .a(_0651_),
    .b(_0682_),
    .c(_0690_),
    .y(_0691_)
  );
  al_mux2l _4810_ (
    .a(\DFF_1205.Q ),
    .b(_0691_),
    .s(_0066_),
    .y(\DFF_1205.D )
  );
  al_mux2l _4811_ (
    .a(\DFF_1206.Q ),
    .b(_0691_),
    .s(_0067_),
    .y(\DFF_1206.D )
  );
  al_mux2l _4812_ (
    .a(\DFF_1207.Q ),
    .b(_0691_),
    .s(_0068_),
    .y(\DFF_1207.D )
  );
  al_and3 _4813_ (
    .a(\DFF_1286.Q ),
    .b(\DFF_1287.Q ),
    .c(_0346_),
    .y(_0692_)
  );
  al_ao21 _4814_ (
    .a(\DFF_1286.Q ),
    .b(_0346_),
    .c(\DFF_1287.Q ),
    .y(_0693_)
  );
  al_and3fft _4815_ (
    .a(_0449_),
    .b(_0692_),
    .c(_0693_),
    .y(\DFF_1287.D )
  );
  al_and2 _4816_ (
    .a(\DFF_86.Q ),
    .b(\DFF_83.Q ),
    .y(_0694_)
  );
  al_and3ftt _4817_ (
    .a(\DFF_85.Q ),
    .b(\DFF_1350.D ),
    .c(_0694_),
    .y(_0695_)
  );
  al_mux2l _4818_ (
    .a(\DFF_1244.Q ),
    .b(_0695_),
    .s(_0454_),
    .y(\DFF_1244.D )
  );
  al_mux2l _4819_ (
    .a(\DFF_1245.Q ),
    .b(_0695_),
    .s(_0457_),
    .y(\DFF_1245.D )
  );
  al_mux2l _4820_ (
    .a(\DFF_1246.Q ),
    .b(_0695_),
    .s(_0458_),
    .y(\DFF_1246.D )
  );
  al_mux2l _4821_ (
    .a(\DFF_1247.Q ),
    .b(\DFF_1360.D ),
    .s(_0454_),
    .y(\DFF_1247.D )
  );
  al_mux2l _4822_ (
    .a(\DFF_1248.Q ),
    .b(\DFF_1360.D ),
    .s(_0457_),
    .y(\DFF_1248.D )
  );
  al_mux2l _4823_ (
    .a(\DFF_1249.Q ),
    .b(\DFF_1360.D ),
    .s(_0458_),
    .y(\DFF_1249.D )
  );
  al_mux2l _4824_ (
    .a(\DFF_1250.Q ),
    .b(\DFF_1362.D ),
    .s(_0454_),
    .y(\DFF_1250.D )
  );
  al_mux2l _4825_ (
    .a(\DFF_1251.Q ),
    .b(\DFF_1362.D ),
    .s(_0457_),
    .y(\DFF_1251.D )
  );
  al_mux2l _4826_ (
    .a(\DFF_1252.Q ),
    .b(\DFF_1362.D ),
    .s(_0458_),
    .y(\DFF_1252.D )
  );
  al_and2 _4827_ (
    .a(\DFF_89.Q ),
    .b(\DFF_90.Q ),
    .y(_0696_)
  );
  al_and3 _4828_ (
    .a(\DFF_84.Q ),
    .b(\DFF_85.Q ),
    .c(_0696_),
    .y(_0697_)
  );
  al_nand3 _4829_ (
    .a(\DFF_87.Q ),
    .b(\DFF_88.Q ),
    .c(_0694_),
    .y(_0698_)
  );
  al_and2ft _4830_ (
    .a(_0698_),
    .b(_0697_),
    .y(_0699_)
  );
  al_inv _4831_ (
    .a(_0699_),
    .y(_0700_)
  );
  al_mux2l _4832_ (
    .a(\DFF_1253.Q ),
    .b(_0700_),
    .s(_0454_),
    .y(\DFF_1253.D )
  );
  al_mux2l _4833_ (
    .a(\DFF_1254.Q ),
    .b(_0700_),
    .s(_0457_),
    .y(\DFF_1254.D )
  );
  al_mux2l _4834_ (
    .a(\DFF_1255.Q ),
    .b(_0700_),
    .s(_0458_),
    .y(\DFF_1255.D )
  );
  al_inv _4835_ (
    .a(_0088_),
    .y(_0701_)
  );
  al_and3 _4836_ (
    .a(\DFF_1512.Q ),
    .b(\DFF_1513.Q ),
    .c(_0324_),
    .y(_0702_)
  );
  al_aoi21 _4837_ (
    .a(\DFF_1512.Q ),
    .b(_0324_),
    .c(\DFF_1513.Q ),
    .y(_0703_)
  );
  al_nor3ftt _4838_ (
    .a(_0701_),
    .b(_0702_),
    .c(_0703_),
    .y(\DFF_1513.D )
  );
  al_nand2ft _4839_ (
    .a(\DFF_1531.Q ),
    .b(\DFF_1504.Q ),
    .y(_0704_)
  );
  al_nand2ft _4840_ (
    .a(\DFF_1532.Q ),
    .b(\DFF_1505.Q ),
    .y(_0705_)
  );
  al_aoi21ftf _4841_ (
    .a(\DFF_1533.Q ),
    .b(\DFF_1506.Q ),
    .c(_0705_),
    .y(_0706_)
  );
  al_ao21 _4842_ (
    .a(_0704_),
    .b(_0706_),
    .c(\DFF_1513.Q ),
    .y(_0707_)
  );
  al_nand3 _4843_ (
    .a(\DFF_1513.Q ),
    .b(_0704_),
    .c(_0706_),
    .y(_0708_)
  );
  al_nand2ft _4844_ (
    .a(\DFF_1541.Q ),
    .b(\DFF_1505.Q ),
    .y(_0709_)
  );
  al_aoi21ftf _4845_ (
    .a(\DFF_1542.Q ),
    .b(\DFF_1506.Q ),
    .c(_0709_),
    .y(_0710_)
  );
  al_ao21ftf _4846_ (
    .a(\DFF_1540.Q ),
    .b(\DFF_1504.Q ),
    .c(_0710_),
    .y(_0711_)
  );
  al_nand2ft _4847_ (
    .a(\DFF_1529.Q ),
    .b(\DFF_1505.Q ),
    .y(_0712_)
  );
  al_aoi21ftf _4848_ (
    .a(\DFF_1530.Q ),
    .b(\DFF_1506.Q ),
    .c(_0712_),
    .y(_0713_)
  );
  al_ao21ftf _4849_ (
    .a(\DFF_1528.Q ),
    .b(\DFF_1504.Q ),
    .c(_0713_),
    .y(_0714_)
  );
  al_nand2 _4850_ (
    .a(_0097_),
    .b(_0714_),
    .y(_0715_)
  );
  al_aoi21ftf _4851_ (
    .a(\DFF_1516.Q ),
    .b(_0711_),
    .c(_0715_),
    .y(_0716_)
  );
  al_and3 _4852_ (
    .a(_0707_),
    .b(_0708_),
    .c(_0716_),
    .y(_0717_)
  );
  al_nand2ft _4853_ (
    .a(\DFF_1535.Q ),
    .b(\DFF_1505.Q ),
    .y(_0718_)
  );
  al_aoi21ftf _4854_ (
    .a(\DFF_1536.Q ),
    .b(\DFF_1506.Q ),
    .c(_0718_),
    .y(_0719_)
  );
  al_ao21ftf _4855_ (
    .a(\DFF_1534.Q ),
    .b(\DFF_1504.Q ),
    .c(_0719_),
    .y(_0720_)
  );
  al_nand2ft _4856_ (
    .a(\DFF_1537.Q ),
    .b(\DFF_1504.Q ),
    .y(_0721_)
  );
  al_nand2ft _4857_ (
    .a(\DFF_1538.Q ),
    .b(\DFF_1505.Q ),
    .y(_0722_)
  );
  al_aoi21ftf _4858_ (
    .a(\DFF_1539.Q ),
    .b(\DFF_1506.Q ),
    .c(_0722_),
    .y(_0723_)
  );
  al_ao21 _4859_ (
    .a(_0721_),
    .b(_0723_),
    .c(\DFF_1515.Q ),
    .y(_0724_)
  );
  al_aoi21ttf _4860_ (
    .a(_0099_),
    .b(_0720_),
    .c(_0724_),
    .y(_0725_)
  );
  al_and3 _4861_ (
    .a(\DFF_1515.Q ),
    .b(_0721_),
    .c(_0723_),
    .y(_0726_)
  );
  al_oa21ftf _4862_ (
    .a(\DFF_1512.Q ),
    .b(_0714_),
    .c(_0726_),
    .y(_0727_)
  );
  al_and3 _4863_ (
    .a(_0725_),
    .b(_0727_),
    .c(_0717_),
    .y(_0728_)
  );
  al_nand2ft _4864_ (
    .a(\DFF_1544.Q ),
    .b(\DFF_1505.Q ),
    .y(_0729_)
  );
  al_aoi21ftf _4865_ (
    .a(\DFF_1545.Q ),
    .b(\DFF_1506.Q ),
    .c(_0729_),
    .y(_0730_)
  );
  al_ao21ftf _4866_ (
    .a(\DFF_1543.Q ),
    .b(\DFF_1504.Q ),
    .c(_0730_),
    .y(_0731_)
  );
  al_and2 _4867_ (
    .a(_0102_),
    .b(_0731_),
    .y(_0732_)
  );
  al_or2 _4868_ (
    .a(_0102_),
    .b(_0731_),
    .y(_0733_)
  );
  al_nand2ft _4869_ (
    .a(\DFF_1526.Q ),
    .b(\DFF_1505.Q ),
    .y(_0734_)
  );
  al_aoi21ftf _4870_ (
    .a(\DFF_1527.Q ),
    .b(\DFF_1506.Q ),
    .c(_0734_),
    .y(_0735_)
  );
  al_ao21ftf _4871_ (
    .a(\DFF_1525.Q ),
    .b(\DFF_1504.Q ),
    .c(_0735_),
    .y(_0736_)
  );
  al_and2ft _4872_ (
    .a(\DFF_1523.Q ),
    .b(\DFF_1505.Q ),
    .y(_0737_)
  );
  al_and2ft _4873_ (
    .a(\DFF_1522.Q ),
    .b(\DFF_1504.Q ),
    .y(_0738_)
  );
  al_nand2ft _4874_ (
    .a(\DFF_1524.Q ),
    .b(\DFF_1506.Q ),
    .y(_0739_)
  );
  al_nand3fft _4875_ (
    .a(_0737_),
    .b(_0738_),
    .c(_0739_),
    .y(_0740_)
  );
  al_nand2 _4876_ (
    .a(_0095_),
    .b(_0740_),
    .y(_0741_)
  );
  al_oa21 _4877_ (
    .a(_0096_),
    .b(_0736_),
    .c(_0741_),
    .y(_0742_)
  );
  al_and3ftt _4878_ (
    .a(_0732_),
    .b(_0733_),
    .c(_0742_),
    .y(_0743_)
  );
  al_and2ft _4879_ (
    .a(\DFF_1546.Q ),
    .b(\DFF_1504.Q ),
    .y(_0744_)
  );
  al_nand2ft _4880_ (
    .a(\DFF_1547.Q ),
    .b(\DFF_1505.Q ),
    .y(_0745_)
  );
  al_aoi21ftf _4881_ (
    .a(\DFF_1548.Q ),
    .b(\DFF_1506.Q ),
    .c(_0745_),
    .y(_0746_)
  );
  al_aoi21ftf _4882_ (
    .a(_0744_),
    .b(_0746_),
    .c(_0103_),
    .y(_0747_)
  );
  al_nor2 _4883_ (
    .a(_0095_),
    .b(_0740_),
    .y(_0748_)
  );
  al_nand3fft _4884_ (
    .a(_0103_),
    .b(_0744_),
    .c(_0746_),
    .y(_0749_)
  );
  al_nand2ft _4885_ (
    .a(\DFF_1520.Q ),
    .b(\DFF_1505.Q ),
    .y(_0750_)
  );
  al_nand2ft _4886_ (
    .a(\DFF_1519.Q ),
    .b(\DFF_1504.Q ),
    .y(_0751_)
  );
  al_and2ft _4887_ (
    .a(\DFF_1521.Q ),
    .b(\DFF_1506.Q ),
    .y(_0752_)
  );
  al_and3ftt _4888_ (
    .a(_0752_),
    .b(_0750_),
    .c(_0751_),
    .y(_0753_)
  );
  al_aoi21ftf _4889_ (
    .a(_0090_),
    .b(_0753_),
    .c(_0749_),
    .y(_0754_)
  );
  al_nand3fft _4890_ (
    .a(_0747_),
    .b(_0748_),
    .c(_0754_),
    .y(_0755_)
  );
  al_or2 _4891_ (
    .a(\DFF_1509.Q ),
    .b(_0753_),
    .y(_0756_)
  );
  al_aoi21ftf _4892_ (
    .a(_0711_),
    .b(\DFF_1516.Q ),
    .c(_0756_),
    .y(_0757_)
  );
  al_nand2 _4893_ (
    .a(_0096_),
    .b(_0736_),
    .y(_0758_)
  );
  al_or2 _4894_ (
    .a(_0099_),
    .b(_0720_),
    .y(_0759_)
  );
  al_nand3 _4895_ (
    .a(_0758_),
    .b(_0759_),
    .c(_0757_),
    .y(_0760_)
  );
  al_and3fft _4896_ (
    .a(_0755_),
    .b(_0760_),
    .c(_0743_),
    .y(_0761_)
  );
  al_nand2ft _4897_ (
    .a(\DFF_1553.Q ),
    .b(\DFF_1505.Q ),
    .y(_0762_)
  );
  al_aoi21ftf _4898_ (
    .a(\DFF_1554.Q ),
    .b(\DFF_1506.Q ),
    .c(_0762_),
    .y(_0763_)
  );
  al_aoi21ftf _4899_ (
    .a(\DFF_1552.Q ),
    .b(\DFF_1504.Q ),
    .c(_0763_),
    .y(_0764_)
  );
  al_nand2ft _4900_ (
    .a(\DFF_1550.Q ),
    .b(\DFF_1505.Q ),
    .y(_0765_)
  );
  al_nand2ft _4901_ (
    .a(\DFF_1549.Q ),
    .b(\DFF_1504.Q ),
    .y(_0766_)
  );
  al_aoi21ftf _4902_ (
    .a(\DFF_1551.Q ),
    .b(\DFF_1506.Q ),
    .c(_0766_),
    .y(_0767_)
  );
  al_nand3 _4903_ (
    .a(_0765_),
    .b(_0767_),
    .c(_0764_),
    .y(_0768_)
  );
  al_aoi21 _4904_ (
    .a(_0761_),
    .b(_0728_),
    .c(_0768_),
    .y(_0769_)
  );
  al_mux2l _4905_ (
    .a(\DFF_1555.Q ),
    .b(_0769_),
    .s(_0092_),
    .y(\DFF_1555.D )
  );
  al_mux2l _4906_ (
    .a(\DFF_1556.Q ),
    .b(_0769_),
    .s(_0093_),
    .y(\DFF_1556.D )
  );
  al_mux2l _4907_ (
    .a(\DFF_1557.Q ),
    .b(_0769_),
    .s(_0094_),
    .y(\DFF_1557.D )
  );
  al_oa21 _4908_ (
    .a(\DFF_14.Q ),
    .b(_0443_),
    .c(_0329_),
    .y(_0770_)
  );
  al_aoi21ttf _4909_ (
    .a(\DFF_14.Q ),
    .b(_0443_),
    .c(_0770_),
    .y(\DFF_14.D )
  );
  al_nand3 _4910_ (
    .a(\DFF_7.Q ),
    .b(\DFF_8.Q ),
    .c(_0333_),
    .y(_0771_)
  );
  al_nand2ft _4911_ (
    .a(\DFF_8.Q ),
    .b(_0440_),
    .y(_0772_)
  );
  al_and3 _4912_ (
    .a(_0771_),
    .b(_0772_),
    .c(_0261_),
    .y(\DFF_8.D )
  );
  al_aoi21 _4913_ (
    .a(\DFF_1600.Q ),
    .b(\DFF_1563.Q ),
    .c(g3234),
    .y(_0773_)
  );
  al_oa21 _4914_ (
    .a(\DFF_1600.Q ),
    .b(\DFF_1563.Q ),
    .c(_0773_),
    .y(\DFF_1600.D )
  );
  al_oa21 _4915_ (
    .a(\DFF_1610.Q ),
    .b(_0447_),
    .c(_0336_),
    .y(_0774_)
  );
  al_aoi21ttf _4916_ (
    .a(\DFF_1610.Q ),
    .b(_0447_),
    .c(_0774_),
    .y(\DFF_1610.D )
  );
  al_and2 _4917_ (
    .a(\DFF_1604.Q ),
    .b(_0444_),
    .y(_0775_)
  );
  al_or2 _4918_ (
    .a(\DFF_1604.Q ),
    .b(_0444_),
    .y(_0776_)
  );
  al_and3ftt _4919_ (
    .a(_0775_),
    .b(_0776_),
    .c(_0339_),
    .y(\DFF_1604.D )
  );
  al_nand3 _4920_ (
    .a(\DFF_399.Q ),
    .b(\DFF_402.Q ),
    .c(\DFF_1504.Q ),
    .y(_0777_)
  );
  al_ao21ftf _4921_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_107.Q ),
    .c(_0777_),
    .y(\DFF_107.D )
  );
  al_mux2h _4922_ (
    .a(\DFF_108.Q ),
    .b(\DFF_400.D ),
    .s(\DFF_1505.Q ),
    .y(\DFF_108.D )
  );
  al_mux2h _4923_ (
    .a(\DFF_109.Q ),
    .b(\DFF_400.D ),
    .s(\DFF_1506.Q ),
    .y(\DFF_109.D )
  );
  al_inv _4924_ (
    .a(_0449_),
    .y(_0778_)
  );
  al_nand2 _4925_ (
    .a(\DFF_238.Q ),
    .b(_0448_),
    .y(_0779_)
  );
  al_or2 _4926_ (
    .a(\DFF_238.Q ),
    .b(_0448_),
    .y(_0780_)
  );
  al_and3 _4927_ (
    .a(_0778_),
    .b(_0779_),
    .c(_0780_),
    .y(\DFF_238.D )
  );
  al_nand2ft _4928_ (
    .a(\DFF_297.Q ),
    .b(\DFF_1429.Q ),
    .y(_0781_)
  );
  al_aoi21ftf _4929_ (
    .a(\DFF_295.Q ),
    .b(\DFF_1427.Q ),
    .c(_0781_),
    .y(_0782_)
  );
  al_ao21ftf _4930_ (
    .a(\DFF_296.Q ),
    .b(\DFF_1428.Q ),
    .c(_0782_),
    .y(_0783_)
  );
  al_nand2ft _4931_ (
    .a(\DFF_167.Q ),
    .b(\DFF_1427.Q ),
    .y(_0784_)
  );
  al_nand2ft _4932_ (
    .a(\DFF_168.Q ),
    .b(\DFF_1428.Q ),
    .y(_0785_)
  );
  al_aoi21ftf _4933_ (
    .a(\DFF_169.Q ),
    .b(\DFF_1429.Q ),
    .c(_0785_),
    .y(_0786_)
  );
  al_and3 _4934_ (
    .a(\DFF_78.Q ),
    .b(_0784_),
    .c(_0786_),
    .y(_0787_)
  );
  al_aoi21 _4935_ (
    .a(_0784_),
    .b(_0786_),
    .c(\DFF_78.Q ),
    .y(_0788_)
  );
  al_or2 _4936_ (
    .a(_0787_),
    .b(_0788_),
    .y(_0789_)
  );
  al_nand2ft _4937_ (
    .a(\DFF_177.Q ),
    .b(\DFF_1428.Q ),
    .y(_0790_)
  );
  al_aoi21ftf _4938_ (
    .a(\DFF_178.Q ),
    .b(\DFF_1429.Q ),
    .c(_0790_),
    .y(_0791_)
  );
  al_aoi21ftf _4939_ (
    .a(\DFF_176.Q ),
    .b(\DFF_1427.Q ),
    .c(_0791_),
    .y(_0792_)
  );
  al_or2 _4940_ (
    .a(\DFF_304.D ),
    .b(_0792_),
    .y(_0793_)
  );
  al_and2 _4941_ (
    .a(\DFF_304.D ),
    .b(_0792_),
    .y(_0794_)
  );
  al_nand2ft _4942_ (
    .a(_0794_),
    .b(_0793_),
    .y(_0795_)
  );
  al_nand2ft _4943_ (
    .a(\DFF_179.Q ),
    .b(\DFF_1427.Q ),
    .y(_0796_)
  );
  al_nand2ft _4944_ (
    .a(\DFF_180.Q ),
    .b(\DFF_1428.Q ),
    .y(_0797_)
  );
  al_aoi21ftf _4945_ (
    .a(\DFF_181.Q ),
    .b(\DFF_1429.Q ),
    .c(_0797_),
    .y(_0798_)
  );
  al_ao21 _4946_ (
    .a(_0796_),
    .b(_0798_),
    .c(\DFF_302.D ),
    .y(_0799_)
  );
  al_and3 _4947_ (
    .a(\DFF_302.D ),
    .b(_0796_),
    .c(_0798_),
    .y(_0800_)
  );
  al_nand2ft _4948_ (
    .a(_0800_),
    .b(_0799_),
    .y(_0801_)
  );
  al_nand2ft _4949_ (
    .a(\DFF_174.Q ),
    .b(\DFF_1428.Q ),
    .y(_0802_)
  );
  al_aoi21ftf _4950_ (
    .a(\DFF_175.Q ),
    .b(\DFF_1429.Q ),
    .c(_0802_),
    .y(_0803_)
  );
  al_ao21ftf _4951_ (
    .a(\DFF_173.Q ),
    .b(\DFF_1427.Q ),
    .c(_0803_),
    .y(_0804_)
  );
  al_nor2 _4952_ (
    .a(\DFF_306.D ),
    .b(_0804_),
    .y(_0805_)
  );
  al_nand2 _4953_ (
    .a(\DFF_306.D ),
    .b(_0804_),
    .y(_0806_)
  );
  al_nand3ftt _4954_ (
    .a(_0805_),
    .b(_0806_),
    .c(_0801_),
    .y(_0807_)
  );
  al_and3fft _4955_ (
    .a(_0789_),
    .b(_0807_),
    .c(_0795_),
    .y(_0808_)
  );
  al_nand2ft _4956_ (
    .a(\DFF_165.Q ),
    .b(\DFF_1428.Q ),
    .y(_0809_)
  );
  al_aoi21ftf _4957_ (
    .a(\DFF_166.Q ),
    .b(\DFF_1429.Q ),
    .c(_0809_),
    .y(_0810_)
  );
  al_ao21ftf _4958_ (
    .a(\DFF_164.Q ),
    .b(\DFF_1427.Q ),
    .c(_0810_),
    .y(_0811_)
  );
  al_or2 _4959_ (
    .a(\DFF_80.Q ),
    .b(_0811_),
    .y(_0812_)
  );
  al_and2 _4960_ (
    .a(\DFF_80.Q ),
    .b(_0811_),
    .y(_0813_)
  );
  al_nand2ft _4961_ (
    .a(_0813_),
    .b(_0812_),
    .y(_0814_)
  );
  al_nand2ft _4962_ (
    .a(\DFF_192.Q ),
    .b(\DFF_1428.Q ),
    .y(_0815_)
  );
  al_aoi21ftf _4963_ (
    .a(\DFF_193.Q ),
    .b(\DFF_1429.Q ),
    .c(_0815_),
    .y(_0816_)
  );
  al_ao21ftf _4964_ (
    .a(\DFF_191.Q ),
    .b(\DFF_1427.Q ),
    .c(_0816_),
    .y(_0817_)
  );
  al_nand2ft _4965_ (
    .a(_0165_),
    .b(_0817_),
    .y(_0818_)
  );
  al_nand2ft _4966_ (
    .a(_0817_),
    .b(_0165_),
    .y(_0819_)
  );
  al_and2 _4967_ (
    .a(_0819_),
    .b(_0818_),
    .y(_0820_)
  );
  al_nand2ft _4968_ (
    .a(\DFF_188.Q ),
    .b(\DFF_1427.Q ),
    .y(_0821_)
  );
  al_aoi21ftf _4969_ (
    .a(\DFF_190.Q ),
    .b(\DFF_1429.Q ),
    .c(_0821_),
    .y(_0822_)
  );
  al_aoi21ftf _4970_ (
    .a(\DFF_189.Q ),
    .b(\DFF_1428.Q ),
    .c(_0822_),
    .y(_0823_)
  );
  al_and2ft _4971_ (
    .a(_0161_),
    .b(_0823_),
    .y(_0824_)
  );
  al_nand2ft _4972_ (
    .a(_0823_),
    .b(_0161_),
    .y(_0825_)
  );
  al_nand2ft _4973_ (
    .a(_0824_),
    .b(_0825_),
    .y(_0826_)
  );
  al_and3 _4974_ (
    .a(_0814_),
    .b(_0826_),
    .c(_0820_),
    .y(_0827_)
  );
  al_nand2ft _4975_ (
    .a(\DFF_186.Q ),
    .b(\DFF_1428.Q ),
    .y(_0828_)
  );
  al_aoi21ftf _4976_ (
    .a(\DFF_187.Q ),
    .b(\DFF_1429.Q ),
    .c(_0828_),
    .y(_0829_)
  );
  al_ao21ftf _4977_ (
    .a(\DFF_185.Q ),
    .b(\DFF_1427.Q ),
    .c(_0829_),
    .y(_0830_)
  );
  al_or2 _4978_ (
    .a(\DFF_66.Q ),
    .b(_0830_),
    .y(_0831_)
  );
  al_and2 _4979_ (
    .a(\DFF_66.Q ),
    .b(_0830_),
    .y(_0832_)
  );
  al_nand2ft _4980_ (
    .a(_0832_),
    .b(_0831_),
    .y(_0833_)
  );
  al_nand2ft _4981_ (
    .a(\DFF_183.Q ),
    .b(\DFF_1428.Q ),
    .y(_0834_)
  );
  al_aoi21ftf _4982_ (
    .a(\DFF_184.Q ),
    .b(\DFF_1429.Q ),
    .c(_0834_),
    .y(_0835_)
  );
  al_ao21ftf _4983_ (
    .a(\DFF_182.Q ),
    .b(\DFF_1427.Q ),
    .c(_0835_),
    .y(_0836_)
  );
  al_or2 _4984_ (
    .a(\DFF_68.Q ),
    .b(_0836_),
    .y(_0837_)
  );
  al_and2 _4985_ (
    .a(\DFF_68.Q ),
    .b(_0836_),
    .y(_0838_)
  );
  al_nand2ft _4986_ (
    .a(_0838_),
    .b(_0837_),
    .y(_0839_)
  );
  al_nand2ft _4987_ (
    .a(\DFF_171.Q ),
    .b(\DFF_1428.Q ),
    .y(_0840_)
  );
  al_aoi21ftf _4988_ (
    .a(\DFF_172.Q ),
    .b(\DFF_1429.Q ),
    .c(_0840_),
    .y(_0841_)
  );
  al_ao21ftf _4989_ (
    .a(\DFF_170.Q ),
    .b(\DFF_1427.Q ),
    .c(_0841_),
    .y(_0842_)
  );
  al_nor2 _4990_ (
    .a(\DFF_308.D ),
    .b(_0842_),
    .y(_0843_)
  );
  al_and2 _4991_ (
    .a(\DFF_308.D ),
    .b(_0842_),
    .y(_0844_)
  );
  al_nand2ft _4992_ (
    .a(\DFF_195.Q ),
    .b(\DFF_1428.Q ),
    .y(_0845_)
  );
  al_aoi21ftf _4993_ (
    .a(\DFF_196.Q ),
    .b(\DFF_1429.Q ),
    .c(_0845_),
    .y(_0846_)
  );
  al_ao21ftf _4994_ (
    .a(\DFF_194.Q ),
    .b(\DFF_1427.Q ),
    .c(_0846_),
    .y(_0847_)
  );
  al_nand2 _4995_ (
    .a(\DFF_1302.Q ),
    .b(_0847_),
    .y(_0848_)
  );
  al_or3 _4996_ (
    .a(_0848_),
    .b(_0843_),
    .c(_0844_),
    .y(_0849_)
  );
  al_nand3ftt _4997_ (
    .a(_0849_),
    .b(_0833_),
    .c(_0839_),
    .y(_0850_)
  );
  al_and3ftt _4998_ (
    .a(_0850_),
    .b(_0808_),
    .c(_0827_),
    .y(_0851_)
  );
  al_nand2ft _4999_ (
    .a(_0783_),
    .b(_0851_),
    .y(_0852_)
  );
  al_mux2h _5000_ (
    .a(\DFF_295.Q ),
    .b(_0852_),
    .s(_0156_),
    .y(\DFF_295.D )
  );
  al_mux2h _5001_ (
    .a(\DFF_296.Q ),
    .b(_0852_),
    .s(_0157_),
    .y(\DFF_296.D )
  );
  al_mux2h _5002_ (
    .a(\DFF_297.Q ),
    .b(_0852_),
    .s(_0158_),
    .y(\DFF_297.D )
  );
  al_nor3fft _5003_ (
    .a(\DFF_361.Q ),
    .b(_0183_),
    .c(_0180_),
    .y(_0853_)
  );
  al_mux2h _5004_ (
    .a(\DFF_429.Q ),
    .b(_0853_),
    .s(\DFF_1504.Q ),
    .y(\DFF_429.D )
  );
  al_mux2h _5005_ (
    .a(\DFF_430.Q ),
    .b(_0853_),
    .s(\DFF_1505.Q ),
    .y(\DFF_430.D )
  );
  al_mux2h _5006_ (
    .a(\DFF_431.Q ),
    .b(_0853_),
    .s(\DFF_1506.Q ),
    .y(\DFF_431.D )
  );
  al_oa21ftf _5007_ (
    .a(_0019_),
    .b(_0464_),
    .c(_0029_),
    .y(_0854_)
  );
  al_aoi21ftf _5008_ (
    .a(_0019_),
    .b(_0464_),
    .c(_0854_),
    .y(\DFF_464.D )
  );
  al_and3 _5009_ (
    .a(\DFF_586.Q ),
    .b(\DFF_1429.Q ),
    .c(_0393_),
    .y(_0855_)
  );
  al_and3 _5010_ (
    .a(\DFF_588.Q ),
    .b(\DFF_587.Q ),
    .c(_0855_),
    .y(_0856_)
  );
  al_ao21 _5011_ (
    .a(\DFF_587.Q ),
    .b(_0855_),
    .c(\DFF_588.Q ),
    .y(_0857_)
  );
  al_and3fft _5012_ (
    .a(_0449_),
    .b(_0856_),
    .c(_0857_),
    .y(\DFF_588.D )
  );
  al_oai21 _5013_ (
    .a(\DFF_316.Q ),
    .b(\DFF_328.Q ),
    .c(\DFF_1428.Q ),
    .y(_0858_)
  );
  al_nor2 _5014_ (
    .a(\DFF_666.Q ),
    .b(\DFF_678.Q ),
    .y(_0859_)
  );
  al_oa21 _5015_ (
    .a(\DFF_667.Q ),
    .b(\DFF_1428.Q ),
    .c(\DFF_666.Q ),
    .y(_0860_)
  );
  al_ao21 _5016_ (
    .a(_0858_),
    .b(_0860_),
    .c(_0859_),
    .y(\DFF_667.D )
  );
  al_nand2ft _5017_ (
    .a(\DFF_647.Q ),
    .b(\DFF_1429.Q ),
    .y(_0861_)
  );
  al_aoi21ftf _5018_ (
    .a(\DFF_645.Q ),
    .b(\DFF_1427.Q ),
    .c(_0861_),
    .y(_0862_)
  );
  al_ao21ftf _5019_ (
    .a(\DFF_646.Q ),
    .b(\DFF_1428.Q ),
    .c(_0862_),
    .y(_0863_)
  );
  al_nand2ft _5020_ (
    .a(\DFF_533.Q ),
    .b(\DFF_1428.Q ),
    .y(_0864_)
  );
  al_aoi21ftf _5021_ (
    .a(\DFF_534.Q ),
    .b(\DFF_1429.Q ),
    .c(_0864_),
    .y(_0865_)
  );
  al_ao21ftf _5022_ (
    .a(\DFF_532.Q ),
    .b(\DFF_1427.Q ),
    .c(_0865_),
    .y(_0866_)
  );
  al_nor2 _5023_ (
    .a(\DFF_50.Q ),
    .b(_0866_),
    .y(_0867_)
  );
  al_and2 _5024_ (
    .a(\DFF_50.Q ),
    .b(_0866_),
    .y(_0868_)
  );
  al_or2 _5025_ (
    .a(_0868_),
    .b(_0867_),
    .y(_0869_)
  );
  al_nand2ft _5026_ (
    .a(\DFF_518.Q ),
    .b(\DFF_1428.Q ),
    .y(_0870_)
  );
  al_aoi21ftf _5027_ (
    .a(\DFF_519.Q ),
    .b(\DFF_1429.Q ),
    .c(_0870_),
    .y(_0871_)
  );
  al_ao21ftf _5028_ (
    .a(\DFF_517.Q ),
    .b(\DFF_1427.Q ),
    .c(_0871_),
    .y(_0872_)
  );
  al_nor2 _5029_ (
    .a(\DFF_60.Q ),
    .b(_0872_),
    .y(_0873_)
  );
  al_and2 _5030_ (
    .a(\DFF_60.Q ),
    .b(_0872_),
    .y(_0874_)
  );
  al_or2 _5031_ (
    .a(_0874_),
    .b(_0873_),
    .y(_0875_)
  );
  al_nand2ft _5032_ (
    .a(\DFF_523.Q ),
    .b(\DFF_1427.Q ),
    .y(_0876_)
  );
  al_nand2ft _5033_ (
    .a(\DFF_524.Q ),
    .b(\DFF_1428.Q ),
    .y(_0877_)
  );
  al_aoi21ftf _5034_ (
    .a(\DFF_525.Q ),
    .b(\DFF_1429.Q ),
    .c(_0877_),
    .y(_0878_)
  );
  al_ao21 _5035_ (
    .a(_0876_),
    .b(_0878_),
    .c(\DFF_56.Q ),
    .y(_0879_)
  );
  al_and3 _5036_ (
    .a(\DFF_56.Q ),
    .b(_0876_),
    .c(_0878_),
    .y(_0880_)
  );
  al_nand2ft _5037_ (
    .a(_0880_),
    .b(_0879_),
    .y(_0881_)
  );
  al_and3ftt _5038_ (
    .a(_0881_),
    .b(_0869_),
    .c(_0875_),
    .y(_0882_)
  );
  al_nand2ft _5039_ (
    .a(\DFF_514.Q ),
    .b(\DFF_1427.Q ),
    .y(_0883_)
  );
  al_nand2ft _5040_ (
    .a(\DFF_515.Q ),
    .b(\DFF_1428.Q ),
    .y(_0884_)
  );
  al_aoi21ftf _5041_ (
    .a(\DFF_516.Q ),
    .b(\DFF_1429.Q ),
    .c(_0884_),
    .y(_0885_)
  );
  al_and3 _5042_ (
    .a(\DFF_662.D ),
    .b(_0883_),
    .c(_0885_),
    .y(_0886_)
  );
  al_ao21 _5043_ (
    .a(_0883_),
    .b(_0885_),
    .c(\DFF_662.D ),
    .y(_0887_)
  );
  al_nand2ft _5044_ (
    .a(_0886_),
    .b(_0887_),
    .y(_0888_)
  );
  al_nand2ft _5045_ (
    .a(\DFF_536.Q ),
    .b(\DFF_1428.Q ),
    .y(_0889_)
  );
  al_aoi21ftf _5046_ (
    .a(\DFF_537.Q ),
    .b(\DFF_1429.Q ),
    .c(_0889_),
    .y(_0890_)
  );
  al_ao21ftf _5047_ (
    .a(\DFF_535.Q ),
    .b(\DFF_1427.Q ),
    .c(_0890_),
    .y(_0891_)
  );
  al_or2 _5048_ (
    .a(\DFF_648.D ),
    .b(_0891_),
    .y(_0892_)
  );
  al_nand2 _5049_ (
    .a(\DFF_648.D ),
    .b(_0891_),
    .y(_0893_)
  );
  al_nand3 _5050_ (
    .a(_0893_),
    .b(_0892_),
    .c(_0888_),
    .y(_0894_)
  );
  al_nand2ft _5051_ (
    .a(\DFF_530.Q ),
    .b(\DFF_1428.Q ),
    .y(_0895_)
  );
  al_aoi21ftf _5052_ (
    .a(\DFF_531.Q ),
    .b(\DFF_1429.Q ),
    .c(_0895_),
    .y(_0896_)
  );
  al_ao21ftf _5053_ (
    .a(\DFF_529.Q ),
    .b(\DFF_1427.Q ),
    .c(_0896_),
    .y(_0897_)
  );
  al_nor2 _5054_ (
    .a(\DFF_52.Q ),
    .b(_0897_),
    .y(_0898_)
  );
  al_nand2 _5055_ (
    .a(\DFF_52.Q ),
    .b(_0897_),
    .y(_0899_)
  );
  al_nand2ft _5056_ (
    .a(\DFF_543.Q ),
    .b(\DFF_1429.Q ),
    .y(_0900_)
  );
  al_aoi21ftf _5057_ (
    .a(\DFF_541.Q ),
    .b(\DFF_1427.Q ),
    .c(_0900_),
    .y(_0901_)
  );
  al_ao21ftf _5058_ (
    .a(\DFF_542.Q ),
    .b(\DFF_1428.Q ),
    .c(_0901_),
    .y(_0902_)
  );
  al_nand2ft _5059_ (
    .a(\DFF_520.Q ),
    .b(\DFF_1427.Q ),
    .y(_0903_)
  );
  al_nand2ft _5060_ (
    .a(\DFF_521.Q ),
    .b(\DFF_1428.Q ),
    .y(_0904_)
  );
  al_aoi21ftf _5061_ (
    .a(\DFF_522.Q ),
    .b(\DFF_1429.Q ),
    .c(_0904_),
    .y(_0905_)
  );
  al_aoi21 _5062_ (
    .a(_0903_),
    .b(_0905_),
    .c(\DFF_58.Q ),
    .y(_0906_)
  );
  al_oa21ttf _5063_ (
    .a(_0195_),
    .b(_0902_),
    .c(_0906_),
    .y(_0907_)
  );
  al_oa21ftt _5064_ (
    .a(_0899_),
    .b(_0898_),
    .c(_0907_),
    .y(_0908_)
  );
  al_nand2ft _5065_ (
    .a(\DFF_538.Q ),
    .b(\DFF_1427.Q ),
    .y(_0909_)
  );
  al_nand2ft _5066_ (
    .a(\DFF_539.Q ),
    .b(\DFF_1428.Q ),
    .y(_0910_)
  );
  al_aoi21ftf _5067_ (
    .a(\DFF_540.Q ),
    .b(\DFF_1429.Q ),
    .c(_0910_),
    .y(_0911_)
  );
  al_ao21ttf _5068_ (
    .a(_0909_),
    .b(_0911_),
    .c(_0191_),
    .y(_0912_)
  );
  al_nand3ftt _5069_ (
    .a(_0189_),
    .b(_0188_),
    .c(_0190_),
    .y(_0913_)
  );
  al_nand3 _5070_ (
    .a(_0909_),
    .b(_0911_),
    .c(_0913_),
    .y(_0914_)
  );
  al_and3 _5071_ (
    .a(\DFF_58.Q ),
    .b(_0903_),
    .c(_0905_),
    .y(_0915_)
  );
  al_and3ftt _5072_ (
    .a(_0915_),
    .b(_0914_),
    .c(_0912_),
    .y(_0916_)
  );
  al_nand3ftt _5073_ (
    .a(_0193_),
    .b(_0192_),
    .c(_0194_),
    .y(_0917_)
  );
  al_and2ft _5074_ (
    .a(\DFF_526.Q ),
    .b(\DFF_1427.Q ),
    .y(_0918_)
  );
  al_nand2ft _5075_ (
    .a(\DFF_527.Q ),
    .b(\DFF_1428.Q ),
    .y(_0919_)
  );
  al_aoi21ftf _5076_ (
    .a(\DFF_528.Q ),
    .b(\DFF_1429.Q ),
    .c(_0919_),
    .y(_0920_)
  );
  al_ao21ftf _5077_ (
    .a(_0918_),
    .b(_0920_),
    .c(\DFF_654.D ),
    .y(_0921_)
  );
  al_ao21ftf _5078_ (
    .a(_0917_),
    .b(_0902_),
    .c(_0921_),
    .y(_0922_)
  );
  al_and3ftt _5079_ (
    .a(_0918_),
    .b(\DFF_54.Q ),
    .c(_0920_),
    .y(_0923_)
  );
  al_nand2ft _5080_ (
    .a(\DFF_545.Q ),
    .b(\DFF_1428.Q ),
    .y(_0924_)
  );
  al_aoi21ftf _5081_ (
    .a(\DFF_546.Q ),
    .b(\DFF_1429.Q ),
    .c(_0924_),
    .y(_0925_)
  );
  al_aoi21ftf _5082_ (
    .a(\DFF_544.Q ),
    .b(\DFF_1427.Q ),
    .c(_0925_),
    .y(_0926_)
  );
  al_nor3ftt _5083_ (
    .a(\DFF_1302.Q ),
    .b(_0923_),
    .c(_0926_),
    .y(_0927_)
  );
  al_and3ftt _5084_ (
    .a(_0922_),
    .b(_0927_),
    .c(_0916_),
    .y(_0928_)
  );
  al_and3ftt _5085_ (
    .a(_0894_),
    .b(_0908_),
    .c(_0928_),
    .y(_0929_)
  );
  al_nand3ftt _5086_ (
    .a(_0863_),
    .b(_0882_),
    .c(_0929_),
    .y(_0930_)
  );
  al_mux2h _5087_ (
    .a(\DFF_645.Q ),
    .b(_0930_),
    .s(_0156_),
    .y(\DFF_645.D )
  );
  al_mux2h _5088_ (
    .a(\DFF_646.Q ),
    .b(_0930_),
    .s(_0157_),
    .y(\DFF_646.D )
  );
  al_mux2h _5089_ (
    .a(\DFF_647.Q ),
    .b(_0930_),
    .s(_0158_),
    .y(\DFF_647.D )
  );
  al_nor3fft _5090_ (
    .a(\DFF_711.Q ),
    .b(_0207_),
    .c(_0054_),
    .y(_0931_)
  );
  al_mux2h _5091_ (
    .a(\DFF_779.Q ),
    .b(_0931_),
    .s(\DFF_1504.Q ),
    .y(\DFF_779.D )
  );
  al_mux2h _5092_ (
    .a(\DFF_780.Q ),
    .b(_0931_),
    .s(\DFF_1505.Q ),
    .y(\DFF_780.D )
  );
  al_mux2h _5093_ (
    .a(\DFF_781.Q ),
    .b(_0931_),
    .s(\DFF_1506.Q ),
    .y(\DFF_781.D )
  );
  al_nand3ftt _5094_ (
    .a(\DFF_433.Q ),
    .b(\DFF_1505.Q ),
    .c(\DFF_432.Q ),
    .y(_0932_)
  );
  al_oa21 _5095_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_792.Q ),
    .c(_0932_),
    .y(_0933_)
  );
  al_mux2l _5096_ (
    .a(\DFF_783.Q ),
    .b(_0933_),
    .s(\DFF_782.Q ),
    .y(\DFF_792.D )
  );
  al_oa21ftf _5097_ (
    .a(\DFF_750.Q ),
    .b(\DFF_1504.Q ),
    .c(\DFF_752.Q ),
    .y(_0934_)
  );
  al_and2ft _5098_ (
    .a(\DFF_749.Q ),
    .b(\DFF_752.Q ),
    .y(_0935_)
  );
  al_aoi21 _5099_ (
    .a(_0777_),
    .b(_0934_),
    .c(_0935_),
    .y(\DFF_750.D )
  );
  al_oa21ftf _5100_ (
    .a(_0046_),
    .b(_0542_),
    .c(_0035_),
    .y(_0936_)
  );
  al_aoi21ftf _5101_ (
    .a(_0046_),
    .b(_0542_),
    .c(_0936_),
    .y(\DFF_814.D )
  );
  al_and3 _5102_ (
    .a(\DFF_938.Q ),
    .b(\DFF_937.Q ),
    .c(_0394_),
    .y(_0937_)
  );
  al_ao21 _5103_ (
    .a(\DFF_937.Q ),
    .b(_0394_),
    .c(\DFF_938.Q ),
    .y(_0938_)
  );
  al_and3fft _5104_ (
    .a(_0449_),
    .b(_0937_),
    .c(_0938_),
    .y(\DFF_938.D )
  );
  al_nand2ft _5105_ (
    .a(\DFF_997.Q ),
    .b(\DFF_1429.Q ),
    .y(_0939_)
  );
  al_aoi21ftf _5106_ (
    .a(\DFF_995.Q ),
    .b(\DFF_1427.Q ),
    .c(_0939_),
    .y(_0940_)
  );
  al_ao21ftf _5107_ (
    .a(\DFF_996.Q ),
    .b(\DFF_1428.Q ),
    .c(_0940_),
    .y(_0941_)
  );
  al_nand2ft _5108_ (
    .a(\DFF_886.Q ),
    .b(\DFF_1428.Q ),
    .y(_0942_)
  );
  al_aoi21ftf _5109_ (
    .a(\DFF_887.Q ),
    .b(\DFF_1429.Q ),
    .c(_0942_),
    .y(_0943_)
  );
  al_aoi21ftf _5110_ (
    .a(\DFF_885.Q ),
    .b(\DFF_1427.Q ),
    .c(_0943_),
    .y(_0944_)
  );
  al_nor2 _5111_ (
    .a(\DFF_38.Q ),
    .b(_0944_),
    .y(_0945_)
  );
  al_and2 _5112_ (
    .a(\DFF_38.Q ),
    .b(_0944_),
    .y(_0946_)
  );
  al_nor2 _5113_ (
    .a(_0946_),
    .b(_0945_),
    .y(_0947_)
  );
  al_nand2ft _5114_ (
    .a(\DFF_874.Q ),
    .b(\DFF_1428.Q ),
    .y(_0948_)
  );
  al_aoi21ftf _5115_ (
    .a(\DFF_875.Q ),
    .b(\DFF_1429.Q ),
    .c(_0948_),
    .y(_0949_)
  );
  al_ao21ftf _5116_ (
    .a(\DFF_873.Q ),
    .b(\DFF_1427.Q ),
    .c(_0949_),
    .y(_0950_)
  );
  al_nand2 _5117_ (
    .a(\DFF_1006.D ),
    .b(_0950_),
    .y(_0951_)
  );
  al_nor2 _5118_ (
    .a(\DFF_1006.D ),
    .b(_0950_),
    .y(_0952_)
  );
  al_nand3ftt _5119_ (
    .a(_0212_),
    .b(_0211_),
    .c(_0213_),
    .y(_0953_)
  );
  al_and2ft _5120_ (
    .a(\DFF_889.Q ),
    .b(\DFF_1428.Q ),
    .y(_0954_)
  );
  al_and2ft _5121_ (
    .a(\DFF_888.Q ),
    .b(\DFF_1427.Q ),
    .y(_0955_)
  );
  al_nand2ft _5122_ (
    .a(\DFF_890.Q ),
    .b(\DFF_1429.Q ),
    .y(_0956_)
  );
  al_nand3fft _5123_ (
    .a(_0954_),
    .b(_0955_),
    .c(_0956_),
    .y(_0957_)
  );
  al_nand2ft _5124_ (
    .a(_0957_),
    .b(_0953_),
    .y(_0958_)
  );
  al_nand2ft _5125_ (
    .a(_0953_),
    .b(_0957_),
    .y(_0959_)
  );
  al_nand2ft _5126_ (
    .a(\DFF_867.Q ),
    .b(\DFF_1427.Q ),
    .y(_0960_)
  );
  al_nand2ft _5127_ (
    .a(\DFF_868.Q ),
    .b(\DFF_1428.Q ),
    .y(_0961_)
  );
  al_aoi21ftf _5128_ (
    .a(\DFF_869.Q ),
    .b(\DFF_1429.Q ),
    .c(_0961_),
    .y(_0962_)
  );
  al_ao21 _5129_ (
    .a(_0960_),
    .b(_0962_),
    .c(\DFF_1010.D ),
    .y(_0963_)
  );
  al_and3 _5130_ (
    .a(\DFF_1010.D ),
    .b(_0960_),
    .c(_0962_),
    .y(_0964_)
  );
  al_nand2ft _5131_ (
    .a(_0964_),
    .b(_0963_),
    .y(_0965_)
  );
  al_and3 _5132_ (
    .a(_0958_),
    .b(_0959_),
    .c(_0965_),
    .y(_0966_)
  );
  al_and3ftt _5133_ (
    .a(_0952_),
    .b(_0951_),
    .c(_0966_),
    .y(_0967_)
  );
  al_nand2ft _5134_ (
    .a(\DFF_864.Q ),
    .b(\DFF_1427.Q ),
    .y(_0968_)
  );
  al_nand2ft _5135_ (
    .a(\DFF_865.Q ),
    .b(\DFF_1428.Q ),
    .y(_0969_)
  );
  al_aoi21ftf _5136_ (
    .a(\DFF_866.Q ),
    .b(\DFF_1429.Q ),
    .c(_0969_),
    .y(_0970_)
  );
  al_and3 _5137_ (
    .a(\DFF_1012.D ),
    .b(_0968_),
    .c(_0970_),
    .y(_0971_)
  );
  al_ao21 _5138_ (
    .a(_0968_),
    .b(_0970_),
    .c(\DFF_1012.D ),
    .y(_0972_)
  );
  al_nand2ft _5139_ (
    .a(_0971_),
    .b(_0972_),
    .y(_0973_)
  );
  al_nand2ft _5140_ (
    .a(\DFF_892.Q ),
    .b(\DFF_1428.Q ),
    .y(_0974_)
  );
  al_aoi21ftf _5141_ (
    .a(\DFF_893.Q ),
    .b(\DFF_1429.Q ),
    .c(_0974_),
    .y(_0975_)
  );
  al_aoi21ftf _5142_ (
    .a(\DFF_891.Q ),
    .b(\DFF_1427.Q ),
    .c(_0975_),
    .y(_0976_)
  );
  al_or3 _5143_ (
    .a(_0215_),
    .b(_0217_),
    .c(_0976_),
    .y(_0977_)
  );
  al_oai21 _5144_ (
    .a(_0215_),
    .b(_0217_),
    .c(_0976_),
    .y(_0978_)
  );
  al_nand2ft _5145_ (
    .a(\DFF_882.Q ),
    .b(\DFF_1427.Q ),
    .y(_0979_)
  );
  al_nand2ft _5146_ (
    .a(\DFF_883.Q ),
    .b(\DFF_1428.Q ),
    .y(_0980_)
  );
  al_aoi21ftf _5147_ (
    .a(\DFF_884.Q ),
    .b(\DFF_1429.Q ),
    .c(_0980_),
    .y(_0981_)
  );
  al_and3 _5148_ (
    .a(\DFF_1000.D ),
    .b(_0979_),
    .c(_0981_),
    .y(_0982_)
  );
  al_ao21 _5149_ (
    .a(_0979_),
    .b(_0981_),
    .c(\DFF_1000.D ),
    .y(_0983_)
  );
  al_nand2ft _5150_ (
    .a(_0982_),
    .b(_0983_),
    .y(_0984_)
  );
  al_and3 _5151_ (
    .a(_0978_),
    .b(_0977_),
    .c(_0984_),
    .y(_0985_)
  );
  al_nand2ft _5152_ (
    .a(\DFF_877.Q ),
    .b(\DFF_1428.Q ),
    .y(_0986_)
  );
  al_aoi21ftf _5153_ (
    .a(\DFF_878.Q ),
    .b(\DFF_1429.Q ),
    .c(_0986_),
    .y(_0987_)
  );
  al_ao21ftf _5154_ (
    .a(\DFF_876.Q ),
    .b(\DFF_1427.Q ),
    .c(_0987_),
    .y(_0988_)
  );
  al_or2 _5155_ (
    .a(\DFF_41.Q ),
    .b(_0988_),
    .y(_0989_)
  );
  al_and2 _5156_ (
    .a(\DFF_41.Q ),
    .b(_0988_),
    .y(_0990_)
  );
  al_nand2ft _5157_ (
    .a(_0990_),
    .b(_0989_),
    .y(_0991_)
  );
  al_nand2ft _5158_ (
    .a(\DFF_879.Q ),
    .b(\DFF_1427.Q ),
    .y(_0992_)
  );
  al_nand2ft _5159_ (
    .a(\DFF_880.Q ),
    .b(\DFF_1428.Q ),
    .y(_0993_)
  );
  al_aoi21ftf _5160_ (
    .a(\DFF_881.Q ),
    .b(\DFF_1429.Q ),
    .c(_0993_),
    .y(_0994_)
  );
  al_and3 _5161_ (
    .a(\DFF_1002.D ),
    .b(_0992_),
    .c(_0994_),
    .y(_0995_)
  );
  al_ao21 _5162_ (
    .a(_0992_),
    .b(_0994_),
    .c(\DFF_1002.D ),
    .y(_0996_)
  );
  al_nand2ft _5163_ (
    .a(_0995_),
    .b(_0996_),
    .y(_0997_)
  );
  al_nand2ft _5164_ (
    .a(\DFF_871.Q ),
    .b(\DFF_1428.Q ),
    .y(_0998_)
  );
  al_aoi21ftf _5165_ (
    .a(\DFF_872.Q ),
    .b(\DFF_1429.Q ),
    .c(_0998_),
    .y(_0999_)
  );
  al_ao21ftf _5166_ (
    .a(\DFF_870.Q ),
    .b(\DFF_1427.Q ),
    .c(_0999_),
    .y(_1000_)
  );
  al_nor2 _5167_ (
    .a(\DFF_1008.D ),
    .b(_1000_),
    .y(_1001_)
  );
  al_nand2 _5168_ (
    .a(\DFF_1008.D ),
    .b(_1000_),
    .y(_1002_)
  );
  al_nand2ft _5169_ (
    .a(\DFF_895.Q ),
    .b(\DFF_1428.Q ),
    .y(_1003_)
  );
  al_aoi21ftf _5170_ (
    .a(\DFF_896.Q ),
    .b(\DFF_1429.Q ),
    .c(_1003_),
    .y(_1004_)
  );
  al_ao21ftf _5171_ (
    .a(\DFF_894.Q ),
    .b(\DFF_1427.Q ),
    .c(_1004_),
    .y(_1005_)
  );
  al_nand2 _5172_ (
    .a(\DFF_1302.Q ),
    .b(_1005_),
    .y(_1006_)
  );
  al_and3fft _5173_ (
    .a(_1006_),
    .b(_1001_),
    .c(_1002_),
    .y(_1007_)
  );
  al_and3 _5174_ (
    .a(_0997_),
    .b(_1007_),
    .c(_0991_),
    .y(_1008_)
  );
  al_and3 _5175_ (
    .a(_0973_),
    .b(_0985_),
    .c(_1008_),
    .y(_1009_)
  );
  al_and3 _5176_ (
    .a(_0947_),
    .b(_0967_),
    .c(_1009_),
    .y(_1010_)
  );
  al_nand2ft _5177_ (
    .a(_0941_),
    .b(_1010_),
    .y(_1011_)
  );
  al_mux2h _5178_ (
    .a(\DFF_995.Q ),
    .b(_1011_),
    .s(_0156_),
    .y(\DFF_995.D )
  );
  al_mux2h _5179_ (
    .a(\DFF_996.Q ),
    .b(_1011_),
    .s(_0157_),
    .y(\DFF_996.D )
  );
  al_mux2h _5180_ (
    .a(\DFF_997.Q ),
    .b(_1011_),
    .s(_0158_),
    .y(\DFF_997.D )
  );
  al_nor3fft _5181_ (
    .a(\DFF_1061.Q ),
    .b(_0230_),
    .c(_0081_),
    .y(_1012_)
  );
  al_mux2h _5182_ (
    .a(\DFF_1129.Q ),
    .b(_1012_),
    .s(\DFF_1504.Q ),
    .y(\DFF_1129.D )
  );
  al_mux2h _5183_ (
    .a(\DFF_1130.Q ),
    .b(_1012_),
    .s(\DFF_1505.Q ),
    .y(\DFF_1130.D )
  );
  al_mux2h _5184_ (
    .a(\DFF_1131.Q ),
    .b(_1012_),
    .s(\DFF_1506.Q ),
    .y(\DFF_1131.D )
  );
  al_oa21ftf _5185_ (
    .a(_0073_),
    .b(_0621_),
    .c(_0062_),
    .y(_1013_)
  );
  al_aoi21ftf _5186_ (
    .a(_0073_),
    .b(_0621_),
    .c(_1013_),
    .y(\DFF_1164.D )
  );
  al_and3 _5187_ (
    .a(\DFF_1288.Q ),
    .b(\DFF_1287.Q ),
    .c(_0417_),
    .y(_1014_)
  );
  al_ao21 _5188_ (
    .a(\DFF_1287.Q ),
    .b(_0417_),
    .c(\DFF_1288.Q ),
    .y(_1015_)
  );
  al_and3fft _5189_ (
    .a(_0449_),
    .b(_1014_),
    .c(_1015_),
    .y(\DFF_1288.D )
  );
  al_nand2ft _5190_ (
    .a(\DFF_1347.Q ),
    .b(\DFF_1429.Q ),
    .y(_1016_)
  );
  al_aoi21ftf _5191_ (
    .a(\DFF_1345.Q ),
    .b(\DFF_1427.Q ),
    .c(_1016_),
    .y(_1017_)
  );
  al_ao21ftf _5192_ (
    .a(\DFF_1346.Q ),
    .b(\DFF_1428.Q ),
    .c(_1017_),
    .y(_1018_)
  );
  al_nand2ft _5193_ (
    .a(\DFF_1224.Q ),
    .b(\DFF_1428.Q ),
    .y(_1019_)
  );
  al_aoi21ftf _5194_ (
    .a(\DFF_1225.Q ),
    .b(\DFF_1429.Q ),
    .c(_1019_),
    .y(_1020_)
  );
  al_ao21ftf _5195_ (
    .a(\DFF_1223.Q ),
    .b(\DFF_1427.Q ),
    .c(_1020_),
    .y(_1021_)
  );
  al_nand2 _5196_ (
    .a(\DFF_1356.D ),
    .b(_1021_),
    .y(_1022_)
  );
  al_nor2 _5197_ (
    .a(\DFF_1356.D ),
    .b(_1021_),
    .y(_1023_)
  );
  al_or2ft _5198_ (
    .a(_1022_),
    .b(_1023_),
    .y(_1024_)
  );
  al_and2ft _5199_ (
    .a(\DFF_1239.Q ),
    .b(\DFF_1428.Q ),
    .y(_1025_)
  );
  al_and2ft _5200_ (
    .a(\DFF_1238.Q ),
    .b(\DFF_1427.Q ),
    .y(_1026_)
  );
  al_nand2ft _5201_ (
    .a(\DFF_1240.Q ),
    .b(\DFF_1429.Q ),
    .y(_1027_)
  );
  al_nand3fft _5202_ (
    .a(_1025_),
    .b(_1026_),
    .c(_1027_),
    .y(_1028_)
  );
  al_and2ft _5203_ (
    .a(_1028_),
    .b(_0236_),
    .y(_1029_)
  );
  al_or2ft _5204_ (
    .a(_1028_),
    .b(_0236_),
    .y(_1030_)
  );
  al_nand2ft _5205_ (
    .a(\DFF_1217.Q ),
    .b(\DFF_1427.Q ),
    .y(_1031_)
  );
  al_nand2ft _5206_ (
    .a(\DFF_1218.Q ),
    .b(\DFF_1428.Q ),
    .y(_1032_)
  );
  al_aoi21ftf _5207_ (
    .a(\DFF_1219.Q ),
    .b(\DFF_1429.Q ),
    .c(_1032_),
    .y(_1033_)
  );
  al_ao21 _5208_ (
    .a(_1031_),
    .b(_1033_),
    .c(\DFF_1360.D ),
    .y(_1034_)
  );
  al_and3 _5209_ (
    .a(\DFF_1360.D ),
    .b(_1031_),
    .c(_1033_),
    .y(_1035_)
  );
  al_nand2ft _5210_ (
    .a(_1035_),
    .b(_1034_),
    .y(_1036_)
  );
  al_and3ftt _5211_ (
    .a(_1029_),
    .b(_1030_),
    .c(_1036_),
    .y(_1037_)
  );
  al_nand2ft _5212_ (
    .a(\DFF_1236.Q ),
    .b(\DFF_1428.Q ),
    .y(_1038_)
  );
  al_aoi21ftf _5213_ (
    .a(\DFF_1237.Q ),
    .b(\DFF_1429.Q ),
    .c(_1038_),
    .y(_1039_)
  );
  al_ao21ftf _5214_ (
    .a(\DFF_1235.Q ),
    .b(\DFF_1427.Q ),
    .c(_1039_),
    .y(_1040_)
  );
  al_nand2 _5215_ (
    .a(\DFF_1348.D ),
    .b(_1040_),
    .y(_1041_)
  );
  al_or2 _5216_ (
    .a(\DFF_1348.D ),
    .b(_1040_),
    .y(_1042_)
  );
  al_and2 _5217_ (
    .a(_1041_),
    .b(_1042_),
    .y(_1043_)
  );
  al_nand3ftt _5218_ (
    .a(_1024_),
    .b(_1037_),
    .c(_1043_),
    .y(_1044_)
  );
  al_nand2ft _5219_ (
    .a(\DFF_1215.Q ),
    .b(\DFF_1428.Q ),
    .y(_1045_)
  );
  al_aoi21ftf _5220_ (
    .a(\DFF_1216.Q ),
    .b(\DFF_1429.Q ),
    .c(_1045_),
    .y(_1046_)
  );
  al_ao21ftf _5221_ (
    .a(\DFF_1214.Q ),
    .b(\DFF_1427.Q ),
    .c(_1046_),
    .y(_1047_)
  );
  al_or2 _5222_ (
    .a(\DFF_90.Q ),
    .b(_1047_),
    .y(_1048_)
  );
  al_and2 _5223_ (
    .a(\DFF_90.Q ),
    .b(_1047_),
    .y(_1049_)
  );
  al_nand2ft _5224_ (
    .a(_1049_),
    .b(_1048_),
    .y(_1050_)
  );
  al_nand2ft _5225_ (
    .a(\DFF_1242.Q ),
    .b(\DFF_1428.Q ),
    .y(_1051_)
  );
  al_aoi21ftf _5226_ (
    .a(\DFF_1243.Q ),
    .b(\DFF_1429.Q ),
    .c(_1051_),
    .y(_1052_)
  );
  al_aoi21ftf _5227_ (
    .a(\DFF_1241.Q ),
    .b(\DFF_1427.Q ),
    .c(_1052_),
    .y(_1053_)
  );
  al_nor2 _5228_ (
    .a(_0240_),
    .b(_1053_),
    .y(_1054_)
  );
  al_nand2 _5229_ (
    .a(_0240_),
    .b(_1053_),
    .y(_1055_)
  );
  al_and2ft _5230_ (
    .a(_1054_),
    .b(_1055_),
    .y(_1056_)
  );
  al_nand2ft _5231_ (
    .a(\DFF_1233.Q ),
    .b(\DFF_1428.Q ),
    .y(_1057_)
  );
  al_aoi21ftf _5232_ (
    .a(\DFF_1234.Q ),
    .b(\DFF_1429.Q ),
    .c(_1057_),
    .y(_1058_)
  );
  al_aoi21ftf _5233_ (
    .a(\DFF_1232.Q ),
    .b(\DFF_1427.Q ),
    .c(_1058_),
    .y(_1059_)
  );
  al_nand2 _5234_ (
    .a(\DFF_1350.D ),
    .b(_1059_),
    .y(_1060_)
  );
  al_ao21ftf _5235_ (
    .a(\DFF_1232.Q ),
    .b(\DFF_1427.Q ),
    .c(_1058_),
    .y(_1061_)
  );
  al_and2 _5236_ (
    .a(\DFF_84.Q ),
    .b(_1061_),
    .y(_1062_)
  );
  al_nand2ft _5237_ (
    .a(_1062_),
    .b(_1060_),
    .y(_1063_)
  );
  al_and3 _5238_ (
    .a(_1050_),
    .b(_1063_),
    .c(_1056_),
    .y(_1064_)
  );
  al_nand2ft _5239_ (
    .a(\DFF_1227.Q ),
    .b(\DFF_1428.Q ),
    .y(_1065_)
  );
  al_aoi21ftf _5240_ (
    .a(\DFF_1228.Q ),
    .b(\DFF_1429.Q ),
    .c(_1065_),
    .y(_1066_)
  );
  al_ao21ftf _5241_ (
    .a(\DFF_1226.Q ),
    .b(\DFF_1427.Q ),
    .c(_1066_),
    .y(_1067_)
  );
  al_nor2 _5242_ (
    .a(\DFF_86.Q ),
    .b(_1067_),
    .y(_1068_)
  );
  al_and2 _5243_ (
    .a(\DFF_86.Q ),
    .b(_1067_),
    .y(_1069_)
  );
  al_or2 _5244_ (
    .a(_1069_),
    .b(_1068_),
    .y(_1070_)
  );
  al_nand2ft _5245_ (
    .a(\DFF_1230.Q ),
    .b(\DFF_1428.Q ),
    .y(_1071_)
  );
  al_aoi21ftf _5246_ (
    .a(\DFF_1231.Q ),
    .b(\DFF_1429.Q ),
    .c(_1071_),
    .y(_1072_)
  );
  al_ao21ftf _5247_ (
    .a(\DFF_1229.Q ),
    .b(\DFF_1427.Q ),
    .c(_1072_),
    .y(_1073_)
  );
  al_or2 _5248_ (
    .a(\DFF_85.Q ),
    .b(_1073_),
    .y(_1074_)
  );
  al_and2 _5249_ (
    .a(\DFF_85.Q ),
    .b(_1073_),
    .y(_1075_)
  );
  al_nand2ft _5250_ (
    .a(_1075_),
    .b(_1074_),
    .y(_1076_)
  );
  al_nand2ft _5251_ (
    .a(\DFF_1221.Q ),
    .b(\DFF_1428.Q ),
    .y(_1077_)
  );
  al_aoi21ftf _5252_ (
    .a(\DFF_1222.Q ),
    .b(\DFF_1429.Q ),
    .c(_1077_),
    .y(_1078_)
  );
  al_ao21ftf _5253_ (
    .a(\DFF_1220.Q ),
    .b(\DFF_1427.Q ),
    .c(_1078_),
    .y(_1079_)
  );
  al_nor2 _5254_ (
    .a(\DFF_1358.D ),
    .b(_1079_),
    .y(_1080_)
  );
  al_nand2 _5255_ (
    .a(\DFF_1358.D ),
    .b(_1079_),
    .y(_1081_)
  );
  al_nand2ft _5256_ (
    .a(\DFF_1245.Q ),
    .b(\DFF_1428.Q ),
    .y(_1082_)
  );
  al_aoi21ftf _5257_ (
    .a(\DFF_1246.Q ),
    .b(\DFF_1429.Q ),
    .c(_1082_),
    .y(_1083_)
  );
  al_ao21ftf _5258_ (
    .a(\DFF_1244.Q ),
    .b(\DFF_1427.Q ),
    .c(_1083_),
    .y(_1084_)
  );
  al_and2 _5259_ (
    .a(\DFF_1302.Q ),
    .b(_1084_),
    .y(_1085_)
  );
  al_or3fft _5260_ (
    .a(_1081_),
    .b(_1085_),
    .c(_1080_),
    .y(_1086_)
  );
  al_and3ftt _5261_ (
    .a(_1086_),
    .b(_1070_),
    .c(_1076_),
    .y(_1087_)
  );
  al_and3ftt _5262_ (
    .a(_1044_),
    .b(_1064_),
    .c(_1087_),
    .y(_1088_)
  );
  al_nand2ft _5263_ (
    .a(_1018_),
    .b(_1088_),
    .y(_1089_)
  );
  al_mux2h _5264_ (
    .a(\DFF_1345.Q ),
    .b(_1089_),
    .s(_0156_),
    .y(\DFF_1345.D )
  );
  al_mux2h _5265_ (
    .a(\DFF_1346.Q ),
    .b(_1089_),
    .s(_0157_),
    .y(\DFF_1346.D )
  );
  al_mux2h _5266_ (
    .a(\DFF_1347.Q ),
    .b(_1089_),
    .s(_0158_),
    .y(\DFF_1347.D )
  );
  al_and3 _5267_ (
    .a(\DFF_1411.Q ),
    .b(_0107_),
    .c(_0252_),
    .y(_1090_)
  );
  al_mux2h _5268_ (
    .a(\DFF_1479.Q ),
    .b(_1090_),
    .s(\DFF_1504.Q ),
    .y(\DFF_1479.D )
  );
  al_mux2h _5269_ (
    .a(\DFF_1480.Q ),
    .b(_1090_),
    .s(\DFF_1505.Q ),
    .y(\DFF_1480.D )
  );
  al_mux2h _5270_ (
    .a(\DFF_1481.Q ),
    .b(_1090_),
    .s(\DFF_1506.Q ),
    .y(\DFF_1481.D )
  );
  al_oa21ftf _5271_ (
    .a(_0099_),
    .b(_0702_),
    .c(_0088_),
    .y(_1091_)
  );
  al_aoi21ftf _5272_ (
    .a(_0099_),
    .b(_0702_),
    .c(_1091_),
    .y(\DFF_1514.D )
  );
  al_nor3fft _5273_ (
    .a(\DFF_8.Q ),
    .b(\DFF_9.Q ),
    .c(_0440_),
    .y(_1092_)
  );
  al_oai21ftf _5274_ (
    .a(\DFF_8.Q ),
    .b(_0440_),
    .c(\DFF_9.Q ),
    .y(_1093_)
  );
  al_and3ftt _5275_ (
    .a(_1092_),
    .b(_1093_),
    .c(_0261_),
    .y(\DFF_9.D )
  );
  al_aoi21 _5276_ (
    .a(\DFF_1600.Q ),
    .b(\DFF_1563.Q ),
    .c(\DFF_1601.Q ),
    .y(_1094_)
  );
  al_nor2 _5277_ (
    .a(_1094_),
    .b(_0340_),
    .y(_1095_)
  );
  al_ao21ttf _5278_ (
    .a(\DFF_1563.Q ),
    .b(_0006_),
    .c(_1095_),
    .y(_1096_)
  );
  al_nand2ft _5279_ (
    .a(g3234),
    .b(_1096_),
    .y(\DFF_1601.D )
  );
  al_ao21 _5280_ (
    .a(\DFF_1604.Q ),
    .b(_0444_),
    .c(\DFF_1605.Q ),
    .y(_1097_)
  );
  al_inv _5281_ (
    .a(\DFF_1605.Q ),
    .y(_1098_)
  );
  al_nand3fft _5282_ (
    .a(_0176_),
    .b(_1098_),
    .c(_0444_),
    .y(_1099_)
  );
  al_and3 _5283_ (
    .a(_1099_),
    .b(_1097_),
    .c(_0339_),
    .y(\DFF_1605.D )
  );
  al_and3 _5284_ (
    .a(\DFF_239.Q ),
    .b(\DFF_238.Q ),
    .c(_0448_),
    .y(_1100_)
  );
  al_aoi21 _5285_ (
    .a(\DFF_238.Q ),
    .b(_0448_),
    .c(\DFF_239.Q ),
    .y(_1101_)
  );
  al_nor3ftt _5286_ (
    .a(_0778_),
    .b(_1100_),
    .c(_1101_),
    .y(\DFF_239.D )
  );
  al_inv _5287_ (
    .a(\DFF_1302.Q ),
    .y(_1102_)
  );
  al_and2 _5288_ (
    .a(\DFF_274.Q ),
    .b(\DFF_1427.Q ),
    .y(_1103_)
  );
  al_aoi21 _5289_ (
    .a(\DFF_276.Q ),
    .b(\DFF_1429.Q ),
    .c(_1103_),
    .y(_1104_)
  );
  al_aoi21ftf _5290_ (
    .a(_0246_),
    .b(\DFF_275.Q ),
    .c(_1104_),
    .y(_1105_)
  );
  al_nand2ft _5291_ (
    .a(\DFF_205.Q ),
    .b(\DFF_1429.Q ),
    .y(_1106_)
  );
  al_aoi21ftf _5292_ (
    .a(\DFF_204.Q ),
    .b(\DFF_1428.Q ),
    .c(_1106_),
    .y(_1107_)
  );
  al_ao21ftf _5293_ (
    .a(\DFF_203.Q ),
    .b(\DFF_1427.Q ),
    .c(_1107_),
    .y(_1108_)
  );
  al_or3fft _5294_ (
    .a(\DFF_1302.Q ),
    .b(_1108_),
    .c(_0462_),
    .y(_1109_)
  );
  al_ao21ftf _5295_ (
    .a(_1105_),
    .b(_1102_),
    .c(_1109_),
    .y(_1110_)
  );
  al_mux2h _5296_ (
    .a(\DFF_274.Q ),
    .b(_1110_),
    .s(\DFF_1427.Q ),
    .y(\DFF_274.D )
  );
  al_mux2h _5297_ (
    .a(\DFF_275.Q ),
    .b(_1110_),
    .s(\DFF_1428.Q ),
    .y(\DFF_275.D )
  );
  al_mux2h _5298_ (
    .a(\DFF_276.Q ),
    .b(_1110_),
    .s(\DFF_1429.Q ),
    .y(\DFF_276.D )
  );
  al_nand2ft _5299_ (
    .a(\DFF_282.Q ),
    .b(\DFF_1429.Q ),
    .y(_1111_)
  );
  al_aoi21ftf _5300_ (
    .a(\DFF_280.Q ),
    .b(\DFF_1427.Q ),
    .c(_1111_),
    .y(_1112_)
  );
  al_ao21ftf _5301_ (
    .a(\DFF_281.Q ),
    .b(\DFF_1428.Q ),
    .c(_1112_),
    .y(_1113_)
  );
  al_oai21ftt _5302_ (
    .a(_1108_),
    .b(_0462_),
    .c(_1105_),
    .y(_1114_)
  );
  al_ao21ftf _5303_ (
    .a(_1105_),
    .b(_0174_),
    .c(_1114_),
    .y(_1115_)
  );
  al_oai21ftt _5304_ (
    .a(_1108_),
    .b(_0462_),
    .c(_0174_),
    .y(_1116_)
  );
  al_and3 _5305_ (
    .a(\DFF_1302.Q ),
    .b(_1116_),
    .c(_1115_),
    .y(_1117_)
  );
  al_and3 _5306_ (
    .a(_0174_),
    .b(_1113_),
    .c(_1117_),
    .y(_1118_)
  );
  al_ao21 _5307_ (
    .a(_1113_),
    .b(_1117_),
    .c(_0174_),
    .y(_1119_)
  );
  al_nand2ft _5308_ (
    .a(_1118_),
    .b(_1119_),
    .y(_1120_)
  );
  al_mux2h _5309_ (
    .a(\DFF_277.Q ),
    .b(_1120_),
    .s(\DFF_1427.Q ),
    .y(\DFF_277.D )
  );
  al_mux2h _5310_ (
    .a(\DFF_278.Q ),
    .b(_1120_),
    .s(\DFF_1428.Q ),
    .y(\DFF_278.D )
  );
  al_mux2h _5311_ (
    .a(\DFF_279.Q ),
    .b(_1120_),
    .s(\DFF_1429.Q ),
    .y(\DFF_279.D )
  );
  al_and3 _5312_ (
    .a(\DFF_464.Q ),
    .b(\DFF_465.Q ),
    .c(_0464_),
    .y(_1121_)
  );
  al_aoi21 _5313_ (
    .a(\DFF_464.Q ),
    .b(_0464_),
    .c(\DFF_465.Q ),
    .y(_1122_)
  );
  al_nor3ftt _5314_ (
    .a(_0463_),
    .b(_1121_),
    .c(_1122_),
    .y(\DFF_465.D )
  );
  al_and3 _5315_ (
    .a(\DFF_589.Q ),
    .b(\DFF_588.Q ),
    .c(_0533_),
    .y(_1123_)
  );
  al_aoi21 _5316_ (
    .a(\DFF_588.Q ),
    .b(_0533_),
    .c(\DFF_589.Q ),
    .y(_1124_)
  );
  al_nor3ftt _5317_ (
    .a(_0778_),
    .b(_1123_),
    .c(_1124_),
    .y(\DFF_589.D )
  );
  al_nand2ft _5318_ (
    .a(\DFF_555.Q ),
    .b(\DFF_1429.Q ),
    .y(_1125_)
  );
  al_aoi21ftf _5319_ (
    .a(\DFF_554.Q ),
    .b(\DFF_1428.Q ),
    .c(_1125_),
    .y(_1126_)
  );
  al_ao21ftf _5320_ (
    .a(\DFF_553.Q ),
    .b(\DFF_1427.Q ),
    .c(_1126_),
    .y(_1127_)
  );
  al_nand3fft _5321_ (
    .a(_0538_),
    .b(_0539_),
    .c(_1127_),
    .y(_1128_)
  );
  al_and2 _5322_ (
    .a(\DFF_625.Q ),
    .b(\DFF_1428.Q ),
    .y(_1129_)
  );
  al_and2 _5323_ (
    .a(\DFF_624.Q ),
    .b(\DFF_1427.Q ),
    .y(_1130_)
  );
  al_aoi21 _5324_ (
    .a(\DFF_626.Q ),
    .b(\DFF_1429.Q ),
    .c(_1130_),
    .y(_1131_)
  );
  al_and3ftt _5325_ (
    .a(_1129_),
    .b(_1102_),
    .c(_1131_),
    .y(_1132_)
  );
  al_aoi21 _5326_ (
    .a(\DFF_1302.Q ),
    .b(_1128_),
    .c(_1132_),
    .y(_1133_)
  );
  al_mux2h _5327_ (
    .a(\DFF_624.Q ),
    .b(_1133_),
    .s(\DFF_1427.Q ),
    .y(\DFF_624.D )
  );
  al_mux2h _5328_ (
    .a(\DFF_625.Q ),
    .b(_1133_),
    .s(\DFF_1428.Q ),
    .y(\DFF_625.D )
  );
  al_mux2h _5329_ (
    .a(\DFF_626.Q ),
    .b(_1133_),
    .s(\DFF_1429.Q ),
    .y(\DFF_626.D )
  );
  al_nand2ft _5330_ (
    .a(\DFF_632.Q ),
    .b(\DFF_1429.Q ),
    .y(_1134_)
  );
  al_aoi21ftf _5331_ (
    .a(\DFF_630.Q ),
    .b(\DFF_1427.Q ),
    .c(_1134_),
    .y(_1135_)
  );
  al_ao21ftf _5332_ (
    .a(\DFF_631.Q ),
    .b(\DFF_1428.Q ),
    .c(_1135_),
    .y(_1136_)
  );
  al_and2ft _5333_ (
    .a(_1129_),
    .b(_1131_),
    .y(_1137_)
  );
  al_mux2h _5334_ (
    .a(_0203_),
    .b(_1128_),
    .s(_1137_),
    .y(_1138_)
  );
  al_nand2 _5335_ (
    .a(_0203_),
    .b(_1128_),
    .y(_1139_)
  );
  al_and3 _5336_ (
    .a(\DFF_1302.Q ),
    .b(_1139_),
    .c(_1138_),
    .y(_1140_)
  );
  al_and3 _5337_ (
    .a(_0203_),
    .b(_1136_),
    .c(_1140_),
    .y(_1141_)
  );
  al_ao21 _5338_ (
    .a(_1136_),
    .b(_1140_),
    .c(_0203_),
    .y(_1142_)
  );
  al_nand2ft _5339_ (
    .a(_1141_),
    .b(_1142_),
    .y(_1143_)
  );
  al_mux2h _5340_ (
    .a(\DFF_627.Q ),
    .b(_1143_),
    .s(\DFF_1427.Q ),
    .y(\DFF_627.D )
  );
  al_mux2h _5341_ (
    .a(\DFF_628.Q ),
    .b(_1143_),
    .s(\DFF_1428.Q ),
    .y(\DFF_628.D )
  );
  al_mux2h _5342_ (
    .a(\DFF_629.Q ),
    .b(_1143_),
    .s(\DFF_1429.Q ),
    .y(\DFF_629.D )
  );
  al_and3 _5343_ (
    .a(\DFF_814.Q ),
    .b(\DFF_815.Q ),
    .c(_0542_),
    .y(_1144_)
  );
  al_aoi21 _5344_ (
    .a(\DFF_814.Q ),
    .b(_0542_),
    .c(\DFF_815.Q ),
    .y(_1145_)
  );
  al_nor3ftt _5345_ (
    .a(_0541_),
    .b(_1144_),
    .c(_1145_),
    .y(\DFF_815.D )
  );
  al_and3 _5346_ (
    .a(\DFF_939.Q ),
    .b(\DFF_938.Q ),
    .c(_0611_),
    .y(_1146_)
  );
  al_aoi21 _5347_ (
    .a(\DFF_938.Q ),
    .b(_0611_),
    .c(\DFF_939.Q ),
    .y(_1147_)
  );
  al_nor3ftt _5348_ (
    .a(_0778_),
    .b(_1146_),
    .c(_1147_),
    .y(\DFF_939.D )
  );
  al_nand2ft _5349_ (
    .a(\DFF_905.Q ),
    .b(\DFF_1429.Q ),
    .y(_1148_)
  );
  al_aoi21ftf _5350_ (
    .a(\DFF_904.Q ),
    .b(\DFF_1428.Q ),
    .c(_1148_),
    .y(_1149_)
  );
  al_ao21ftf _5351_ (
    .a(\DFF_903.Q ),
    .b(\DFF_1427.Q ),
    .c(_1149_),
    .y(_1150_)
  );
  al_nand3ftt _5352_ (
    .a(_0617_),
    .b(_0616_),
    .c(_1150_),
    .y(_1151_)
  );
  al_and2 _5353_ (
    .a(\DFF_975.Q ),
    .b(\DFF_1428.Q ),
    .y(_1152_)
  );
  al_and2 _5354_ (
    .a(\DFF_974.Q ),
    .b(\DFF_1427.Q ),
    .y(_1153_)
  );
  al_aoi21 _5355_ (
    .a(\DFF_976.Q ),
    .b(\DFF_1429.Q ),
    .c(_1153_),
    .y(_1154_)
  );
  al_and3ftt _5356_ (
    .a(_1152_),
    .b(_1102_),
    .c(_1154_),
    .y(_1155_)
  );
  al_aoi21 _5357_ (
    .a(\DFF_1302.Q ),
    .b(_1151_),
    .c(_1155_),
    .y(_1156_)
  );
  al_mux2h _5358_ (
    .a(\DFF_974.Q ),
    .b(_1156_),
    .s(\DFF_1427.Q ),
    .y(\DFF_974.D )
  );
  al_mux2h _5359_ (
    .a(\DFF_975.Q ),
    .b(_1156_),
    .s(\DFF_1428.Q ),
    .y(\DFF_975.D )
  );
  al_mux2h _5360_ (
    .a(\DFF_976.Q ),
    .b(_1156_),
    .s(\DFF_1429.Q ),
    .y(\DFF_976.D )
  );
  al_nand2ft _5361_ (
    .a(\DFF_982.Q ),
    .b(\DFF_1429.Q ),
    .y(_1157_)
  );
  al_aoi21ftf _5362_ (
    .a(\DFF_980.Q ),
    .b(\DFF_1427.Q ),
    .c(_1157_),
    .y(_1158_)
  );
  al_ao21ftf _5363_ (
    .a(\DFF_981.Q ),
    .b(\DFF_1428.Q ),
    .c(_1158_),
    .y(_1159_)
  );
  al_and2ft _5364_ (
    .a(_1152_),
    .b(_1154_),
    .y(_1160_)
  );
  al_mux2h _5365_ (
    .a(_0226_),
    .b(_1151_),
    .s(_1160_),
    .y(_1161_)
  );
  al_nand2 _5366_ (
    .a(_0226_),
    .b(_1151_),
    .y(_1162_)
  );
  al_and3 _5367_ (
    .a(\DFF_1302.Q ),
    .b(_1162_),
    .c(_1161_),
    .y(_1163_)
  );
  al_and3 _5368_ (
    .a(_0226_),
    .b(_1159_),
    .c(_1163_),
    .y(_1164_)
  );
  al_ao21 _5369_ (
    .a(_1159_),
    .b(_1163_),
    .c(_0226_),
    .y(_1165_)
  );
  al_nand2ft _5370_ (
    .a(_1164_),
    .b(_1165_),
    .y(_1166_)
  );
  al_mux2h _5371_ (
    .a(\DFF_977.Q ),
    .b(_1166_),
    .s(\DFF_1427.Q ),
    .y(\DFF_977.D )
  );
  al_mux2h _5372_ (
    .a(\DFF_978.Q ),
    .b(_1166_),
    .s(\DFF_1428.Q ),
    .y(\DFF_978.D )
  );
  al_mux2h _5373_ (
    .a(\DFF_979.Q ),
    .b(_1166_),
    .s(\DFF_1429.Q ),
    .y(\DFF_979.D )
  );
  al_and3 _5374_ (
    .a(\DFF_1164.Q ),
    .b(\DFF_1165.Q ),
    .c(_0621_),
    .y(_1167_)
  );
  al_aoi21 _5375_ (
    .a(\DFF_1164.Q ),
    .b(_0621_),
    .c(\DFF_1165.Q ),
    .y(_1168_)
  );
  al_nor3ftt _5376_ (
    .a(_0620_),
    .b(_1167_),
    .c(_1168_),
    .y(\DFF_1165.D )
  );
  al_and3 _5377_ (
    .a(\DFF_1289.Q ),
    .b(\DFF_1288.Q ),
    .c(_0692_),
    .y(_1169_)
  );
  al_aoi21 _5378_ (
    .a(\DFF_1288.Q ),
    .b(_0692_),
    .c(\DFF_1289.Q ),
    .y(_1170_)
  );
  al_nor3ftt _5379_ (
    .a(_0778_),
    .b(_1169_),
    .c(_1170_),
    .y(\DFF_1289.D )
  );
  al_nand2ft _5380_ (
    .a(\DFF_1255.Q ),
    .b(\DFF_1429.Q ),
    .y(_1171_)
  );
  al_aoi21ftf _5381_ (
    .a(\DFF_1254.Q ),
    .b(\DFF_1428.Q ),
    .c(_1171_),
    .y(_1172_)
  );
  al_ao21ftf _5382_ (
    .a(\DFF_1253.Q ),
    .b(\DFF_1427.Q ),
    .c(_1172_),
    .y(_1173_)
  );
  al_nand3ftt _5383_ (
    .a(_0698_),
    .b(_0697_),
    .c(_1173_),
    .y(_1174_)
  );
  al_nand2 _5384_ (
    .a(\DFF_1324.Q ),
    .b(\DFF_1427.Q ),
    .y(_1175_)
  );
  al_aoi21ttf _5385_ (
    .a(\DFF_1326.Q ),
    .b(\DFF_1429.Q ),
    .c(_1175_),
    .y(_1176_)
  );
  al_aoi21ftf _5386_ (
    .a(_0246_),
    .b(\DFF_1325.Q ),
    .c(_1176_),
    .y(_1177_)
  );
  al_nand2 _5387_ (
    .a(_1102_),
    .b(_1177_),
    .y(_1178_)
  );
  al_aoi21ttf _5388_ (
    .a(\DFF_1302.Q ),
    .b(_1174_),
    .c(_1178_),
    .y(_1179_)
  );
  al_mux2h _5389_ (
    .a(\DFF_1324.Q ),
    .b(_1179_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1324.D )
  );
  al_mux2h _5390_ (
    .a(\DFF_1325.Q ),
    .b(_1179_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1325.D )
  );
  al_mux2h _5391_ (
    .a(\DFF_1326.Q ),
    .b(_1179_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1326.D )
  );
  al_nand2ft _5392_ (
    .a(\DFF_1330.Q ),
    .b(\DFF_1427.Q ),
    .y(_1180_)
  );
  al_aoi21ftf _5393_ (
    .a(\DFF_1332.Q ),
    .b(\DFF_1429.Q ),
    .c(_1180_),
    .y(_1181_)
  );
  al_aoi21ftf _5394_ (
    .a(\DFF_1331.Q ),
    .b(\DFF_1428.Q ),
    .c(_1181_),
    .y(_1182_)
  );
  al_ao21 _5395_ (
    .a(_1173_),
    .b(_0699_),
    .c(_0249_),
    .y(_1183_)
  );
  al_nand3 _5396_ (
    .a(_1173_),
    .b(_1177_),
    .c(_0699_),
    .y(_1184_)
  );
  al_oai21ftf _5397_ (
    .a(_0249_),
    .b(_1177_),
    .c(_1102_),
    .y(_1185_)
  );
  al_and3ftt _5398_ (
    .a(_1185_),
    .b(_1183_),
    .c(_1184_),
    .y(_1186_)
  );
  al_aoi21ftf _5399_ (
    .a(_1182_),
    .b(_1186_),
    .c(_0249_),
    .y(_1187_)
  );
  al_nand3fft _5400_ (
    .a(_0249_),
    .b(_1182_),
    .c(_1186_),
    .y(_1188_)
  );
  al_or2ft _5401_ (
    .a(_1188_),
    .b(_1187_),
    .y(_1189_)
  );
  al_mux2h _5402_ (
    .a(\DFF_1327.Q ),
    .b(_1189_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1327.D )
  );
  al_mux2h _5403_ (
    .a(\DFF_1328.Q ),
    .b(_1189_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1328.D )
  );
  al_mux2h _5404_ (
    .a(\DFF_1329.Q ),
    .b(_1189_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1329.D )
  );
  al_and3 _5405_ (
    .a(\DFF_1514.Q ),
    .b(\DFF_1515.Q ),
    .c(_0702_),
    .y(_1190_)
  );
  al_aoi21 _5406_ (
    .a(\DFF_1514.Q ),
    .b(_0702_),
    .c(\DFF_1515.Q ),
    .y(_1191_)
  );
  al_nor3ftt _5407_ (
    .a(_0701_),
    .b(_1190_),
    .c(_1191_),
    .y(\DFF_1515.D )
  );
  al_oa21 _5408_ (
    .a(\DFF_10.Q ),
    .b(_1092_),
    .c(_0261_),
    .y(_1192_)
  );
  al_aoi21ttf _5409_ (
    .a(\DFF_10.Q ),
    .b(_1092_),
    .c(_1192_),
    .y(\DFF_10.D )
  );
  al_nand2 _5410_ (
    .a(\DFF_1606.Q ),
    .b(_1099_),
    .y(_1193_)
  );
  al_nand3fft _5411_ (
    .a(\DFF_1606.Q ),
    .b(_1098_),
    .c(_0775_),
    .y(_1194_)
  );
  al_aoi21ttf _5412_ (
    .a(_1193_),
    .b(_1194_),
    .c(_0339_),
    .y(\DFF_1606.D )
  );
  al_inv _5413_ (
    .a(\DFF_240.Q ),
    .y(_1195_)
  );
  al_oa21ftf _5414_ (
    .a(_1195_),
    .b(_1100_),
    .c(_0449_),
    .y(_1196_)
  );
  al_aoi21ftf _5415_ (
    .a(_1195_),
    .b(_1100_),
    .c(_1196_),
    .y(\DFF_240.D )
  );
  al_inv _5416_ (
    .a(\DFF_1427.Q ),
    .y(_1197_)
  );
  al_and2ft _5417_ (
    .a(_0267_),
    .b(_0270_),
    .y(_1198_)
  );
  al_ao21ftt _5418_ (
    .a(_0273_),
    .b(_1198_),
    .c(_0393_),
    .y(_1199_)
  );
  al_nand3fft _5419_ (
    .a(_1197_),
    .b(_0274_),
    .c(_1199_),
    .y(_1200_)
  );
  al_inv _5420_ (
    .a(g3229),
    .y(_1201_)
  );
  al_nand2ft _5421_ (
    .a(\DFF_262.Q ),
    .b(\DFF_1427.Q ),
    .y(_1202_)
  );
  al_aoi21ftf _5422_ (
    .a(\DFF_264.Q ),
    .b(\DFF_1429.Q ),
    .c(_1202_),
    .y(_1203_)
  );
  al_aoi21ftf _5423_ (
    .a(\DFF_263.Q ),
    .b(\DFF_1428.Q ),
    .c(_1203_),
    .y(_1204_)
  );
  al_nand2ft _5424_ (
    .a(\DFF_254.Q ),
    .b(\DFF_1428.Q ),
    .y(_1205_)
  );
  al_aoi21ftf _5425_ (
    .a(\DFF_255.Q ),
    .b(\DFF_1429.Q ),
    .c(_1205_),
    .y(_1206_)
  );
  al_aoi21ftf _5426_ (
    .a(\DFF_253.Q ),
    .b(\DFF_1427.Q ),
    .c(_1206_),
    .y(_1207_)
  );
  al_nand2ft _5427_ (
    .a(\DFF_260.Q ),
    .b(\DFF_1428.Q ),
    .y(_1208_)
  );
  al_aoi21ftf _5428_ (
    .a(\DFF_261.Q ),
    .b(\DFF_1429.Q ),
    .c(_1208_),
    .y(_1209_)
  );
  al_aoi21ftf _5429_ (
    .a(\DFF_259.Q ),
    .b(\DFF_1427.Q ),
    .c(_1209_),
    .y(_1210_)
  );
  al_and2ft _5430_ (
    .a(\DFF_256.Q ),
    .b(\DFF_1427.Q ),
    .y(_1211_)
  );
  al_aoi21ftt _5431_ (
    .a(\DFF_258.Q ),
    .b(\DFF_1429.Q ),
    .c(_1211_),
    .y(_1212_)
  );
  al_ao21ftf _5432_ (
    .a(\DFF_257.Q ),
    .b(\DFF_1428.Q ),
    .c(_1212_),
    .y(_1213_)
  );
  al_nand2 _5433_ (
    .a(_1210_),
    .b(_1213_),
    .y(_1214_)
  );
  al_aoi21ftf _5434_ (
    .a(_1207_),
    .b(_1204_),
    .c(_1214_),
    .y(_1215_)
  );
  al_oai21ftt _5435_ (
    .a(_1204_),
    .b(_1213_),
    .c(_1210_),
    .y(_1216_)
  );
  al_aoi21ftf _5436_ (
    .a(_1207_),
    .b(_1216_),
    .c(_1204_),
    .y(_1217_)
  );
  al_mux2l _5437_ (
    .a(_1215_),
    .b(_1217_),
    .s(_1201_),
    .y(_1218_)
  );
  al_mux2l _5438_ (
    .a(\DFF_253.Q ),
    .b(_1218_),
    .s(_1200_),
    .y(\DFF_253.D )
  );
  al_nand3fft _5439_ (
    .a(_0246_),
    .b(_0274_),
    .c(_1199_),
    .y(_1219_)
  );
  al_mux2l _5440_ (
    .a(\DFF_254.Q ),
    .b(_1218_),
    .s(_1219_),
    .y(\DFF_254.D )
  );
  al_nand3fft _5441_ (
    .a(_0344_),
    .b(_0274_),
    .c(_1199_),
    .y(_1220_)
  );
  al_mux2l _5442_ (
    .a(\DFF_255.Q ),
    .b(_1218_),
    .s(_1220_),
    .y(\DFF_255.D )
  );
  al_or2 _5443_ (
    .a(_1201_),
    .b(_1207_),
    .y(_1221_)
  );
  al_and2 _5444_ (
    .a(_1201_),
    .b(_1207_),
    .y(_1222_)
  );
  al_nand2ft _5445_ (
    .a(_1222_),
    .b(_1221_),
    .y(_1223_)
  );
  al_aoi21ftf _5446_ (
    .a(_1210_),
    .b(_1223_),
    .c(_1214_),
    .y(_1224_)
  );
  al_mux2l _5447_ (
    .a(\DFF_256.Q ),
    .b(_1224_),
    .s(_1200_),
    .y(\DFF_256.D )
  );
  al_mux2l _5448_ (
    .a(\DFF_257.Q ),
    .b(_1224_),
    .s(_1219_),
    .y(\DFF_257.D )
  );
  al_mux2l _5449_ (
    .a(\DFF_258.Q ),
    .b(_1224_),
    .s(_1220_),
    .y(\DFF_258.D )
  );
  al_or2ft _5450_ (
    .a(_1204_),
    .b(_1213_),
    .y(_1225_)
  );
  al_and3fft _5451_ (
    .a(_1213_),
    .b(_1222_),
    .c(_1221_),
    .y(_1226_)
  );
  al_ao21 _5452_ (
    .a(_1225_),
    .b(_1223_),
    .c(_1226_),
    .y(_1227_)
  );
  al_mux2l _5453_ (
    .a(\DFF_259.Q ),
    .b(_1227_),
    .s(_1200_),
    .y(\DFF_259.D )
  );
  al_mux2l _5454_ (
    .a(\DFF_260.Q ),
    .b(_1227_),
    .s(_1219_),
    .y(\DFF_260.D )
  );
  al_mux2l _5455_ (
    .a(\DFF_261.Q ),
    .b(_1227_),
    .s(_1220_),
    .y(\DFF_261.D )
  );
  al_nand2 _5456_ (
    .a(_1210_),
    .b(_1226_),
    .y(_1228_)
  );
  al_mux2l _5457_ (
    .a(\DFF_262.Q ),
    .b(_1228_),
    .s(_1200_),
    .y(\DFF_262.D )
  );
  al_mux2l _5458_ (
    .a(\DFF_263.Q ),
    .b(_1228_),
    .s(_1219_),
    .y(\DFF_263.D )
  );
  al_mux2l _5459_ (
    .a(\DFF_264.Q ),
    .b(_1228_),
    .s(_1220_),
    .y(\DFF_264.D )
  );
  al_nand2 _5460_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_433.D ),
    .y(_1229_)
  );
  al_nand2ft _5461_ (
    .a(\DFF_406.Q ),
    .b(\DFF_1505.Q ),
    .y(_1230_)
  );
  al_aoi21ftf _5462_ (
    .a(\DFF_407.Q ),
    .b(\DFF_1506.Q ),
    .c(_1230_),
    .y(_1231_)
  );
  al_aoi21ftf _5463_ (
    .a(\DFF_405.Q ),
    .b(\DFF_1504.Q ),
    .c(_1231_),
    .y(_1232_)
  );
  al_nand2ft _5464_ (
    .a(\DFF_409.Q ),
    .b(\DFF_1505.Q ),
    .y(_1233_)
  );
  al_aoi21ftf _5465_ (
    .a(\DFF_410.Q ),
    .b(\DFF_1506.Q ),
    .c(_1233_),
    .y(_1234_)
  );
  al_aoi21ftf _5466_ (
    .a(\DFF_408.Q ),
    .b(\DFF_1504.Q ),
    .c(_1234_),
    .y(_1235_)
  );
  al_and2ft _5467_ (
    .a(_1232_),
    .b(_1235_),
    .y(_1236_)
  );
  al_nand2ft _5468_ (
    .a(\DFF_412.Q ),
    .b(\DFF_1505.Q ),
    .y(_1237_)
  );
  al_aoi21ftf _5469_ (
    .a(\DFF_413.Q ),
    .b(\DFF_1506.Q ),
    .c(_1237_),
    .y(_1238_)
  );
  al_aoi21ftf _5470_ (
    .a(\DFF_411.Q ),
    .b(\DFF_1504.Q ),
    .c(_1238_),
    .y(_1239_)
  );
  al_or2 _5471_ (
    .a(_1232_),
    .b(_1239_),
    .y(_1240_)
  );
  al_nand2ft _5472_ (
    .a(\DFF_415.Q ),
    .b(\DFF_1505.Q ),
    .y(_1241_)
  );
  al_aoi21ftf _5473_ (
    .a(\DFF_416.Q ),
    .b(\DFF_1506.Q ),
    .c(_1241_),
    .y(_1242_)
  );
  al_aoi21ftf _5474_ (
    .a(\DFF_414.Q ),
    .b(\DFF_1504.Q ),
    .c(_1242_),
    .y(_1243_)
  );
  al_and3 _5475_ (
    .a(g3229),
    .b(_1243_),
    .c(_1240_),
    .y(_1244_)
  );
  al_nand2ft _5476_ (
    .a(_1235_),
    .b(_1239_),
    .y(_1245_)
  );
  al_nand2ft _5477_ (
    .a(_1232_),
    .b(_1243_),
    .y(_1246_)
  );
  al_nand3 _5478_ (
    .a(_1201_),
    .b(_1246_),
    .c(_1245_),
    .y(_1247_)
  );
  al_ao21ftf _5479_ (
    .a(_1236_),
    .b(_1244_),
    .c(_1247_),
    .y(_1248_)
  );
  al_mux2l _5480_ (
    .a(\DFF_405.Q ),
    .b(_1248_),
    .s(_1229_),
    .y(\DFF_405.D )
  );
  al_nand2 _5481_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_433.D ),
    .y(_1249_)
  );
  al_mux2l _5482_ (
    .a(\DFF_406.Q ),
    .b(_1248_),
    .s(_1249_),
    .y(\DFF_406.D )
  );
  al_nand2 _5483_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_433.D ),
    .y(_1250_)
  );
  al_mux2l _5484_ (
    .a(\DFF_407.Q ),
    .b(_1248_),
    .s(_1250_),
    .y(\DFF_407.D )
  );
  al_nor2 _5485_ (
    .a(g3229),
    .b(_1232_),
    .y(_1251_)
  );
  al_nand2 _5486_ (
    .a(g3229),
    .b(_1232_),
    .y(_1252_)
  );
  al_or2ft _5487_ (
    .a(_1252_),
    .b(_1251_),
    .y(_1253_)
  );
  al_mux2l _5488_ (
    .a(_1235_),
    .b(_1253_),
    .s(_1239_),
    .y(_1254_)
  );
  al_mux2l _5489_ (
    .a(\DFF_408.Q ),
    .b(_1254_),
    .s(_1229_),
    .y(\DFF_408.D )
  );
  al_mux2l _5490_ (
    .a(\DFF_409.Q ),
    .b(_1254_),
    .s(_1249_),
    .y(\DFF_409.D )
  );
  al_mux2l _5491_ (
    .a(\DFF_410.Q ),
    .b(_1254_),
    .s(_1250_),
    .y(\DFF_410.D )
  );
  al_nand2 _5492_ (
    .a(_1235_),
    .b(_1243_),
    .y(_1255_)
  );
  al_mux2l _5493_ (
    .a(_1235_),
    .b(_1255_),
    .s(_1253_),
    .y(_1256_)
  );
  al_mux2l _5494_ (
    .a(\DFF_411.Q ),
    .b(_1256_),
    .s(_1229_),
    .y(\DFF_411.D )
  );
  al_mux2l _5495_ (
    .a(\DFF_412.Q ),
    .b(_1256_),
    .s(_1249_),
    .y(\DFF_412.D )
  );
  al_mux2l _5496_ (
    .a(\DFF_413.Q ),
    .b(_1256_),
    .s(_1250_),
    .y(\DFF_413.D )
  );
  al_nand2 _5497_ (
    .a(_1235_),
    .b(_1239_),
    .y(_1257_)
  );
  al_oai21ftf _5498_ (
    .a(_1252_),
    .b(_1251_),
    .c(_1257_),
    .y(_1258_)
  );
  al_mux2l _5499_ (
    .a(\DFF_414.Q ),
    .b(_1258_),
    .s(_1229_),
    .y(\DFF_414.D )
  );
  al_mux2l _5500_ (
    .a(\DFF_415.Q ),
    .b(_1258_),
    .s(_1249_),
    .y(\DFF_415.D )
  );
  al_mux2l _5501_ (
    .a(\DFF_416.Q ),
    .b(_1258_),
    .s(_1250_),
    .y(\DFF_416.D )
  );
  al_oa21ftf _5502_ (
    .a(_0021_),
    .b(_1121_),
    .c(_0029_),
    .y(_1259_)
  );
  al_aoi21ftf _5503_ (
    .a(_0021_),
    .b(_1121_),
    .c(_1259_),
    .y(\DFF_466.D )
  );
  al_and3 _5504_ (
    .a(\DFF_589.Q ),
    .b(\DFF_590.Q ),
    .c(_0856_),
    .y(_1260_)
  );
  al_aoi21 _5505_ (
    .a(\DFF_589.Q ),
    .b(_0856_),
    .c(\DFF_590.Q ),
    .y(_1261_)
  );
  al_nor3ftt _5506_ (
    .a(_0778_),
    .b(_1260_),
    .c(_1261_),
    .y(\DFF_590.D )
  );
  al_nand2ft _5507_ (
    .a(_0393_),
    .b(_0289_),
    .y(_1262_)
  );
  al_nand3fft _5508_ (
    .a(_1197_),
    .b(_0288_),
    .c(_1262_),
    .y(_1263_)
  );
  al_nand2ft _5509_ (
    .a(\DFF_612.Q ),
    .b(\DFF_1427.Q ),
    .y(_1264_)
  );
  al_aoi21ftf _5510_ (
    .a(\DFF_614.Q ),
    .b(\DFF_1429.Q ),
    .c(_1264_),
    .y(_1265_)
  );
  al_aoi21ftf _5511_ (
    .a(\DFF_613.Q ),
    .b(\DFF_1428.Q ),
    .c(_1265_),
    .y(_1266_)
  );
  al_nand2ft _5512_ (
    .a(\DFF_604.Q ),
    .b(\DFF_1428.Q ),
    .y(_1267_)
  );
  al_aoi21ftf _5513_ (
    .a(\DFF_605.Q ),
    .b(\DFF_1429.Q ),
    .c(_1267_),
    .y(_1268_)
  );
  al_aoi21ftf _5514_ (
    .a(\DFF_603.Q ),
    .b(\DFF_1427.Q ),
    .c(_1268_),
    .y(_1269_)
  );
  al_nand2ft _5515_ (
    .a(\DFF_610.Q ),
    .b(\DFF_1428.Q ),
    .y(_1270_)
  );
  al_aoi21ftf _5516_ (
    .a(\DFF_611.Q ),
    .b(\DFF_1429.Q ),
    .c(_1270_),
    .y(_1271_)
  );
  al_aoi21ftf _5517_ (
    .a(\DFF_609.Q ),
    .b(\DFF_1427.Q ),
    .c(_1271_),
    .y(_1272_)
  );
  al_and2ft _5518_ (
    .a(\DFF_606.Q ),
    .b(\DFF_1427.Q ),
    .y(_1273_)
  );
  al_aoi21ftt _5519_ (
    .a(\DFF_608.Q ),
    .b(\DFF_1429.Q ),
    .c(_1273_),
    .y(_1274_)
  );
  al_ao21ftf _5520_ (
    .a(\DFF_607.Q ),
    .b(\DFF_1428.Q ),
    .c(_1274_),
    .y(_1275_)
  );
  al_nand2 _5521_ (
    .a(_1272_),
    .b(_1275_),
    .y(_1276_)
  );
  al_aoi21ftf _5522_ (
    .a(_1269_),
    .b(_1266_),
    .c(_1276_),
    .y(_1277_)
  );
  al_oai21ftt _5523_ (
    .a(_1266_),
    .b(_1275_),
    .c(_1272_),
    .y(_1278_)
  );
  al_aoi21ftf _5524_ (
    .a(_1269_),
    .b(_1278_),
    .c(_1266_),
    .y(_1279_)
  );
  al_mux2l _5525_ (
    .a(_1277_),
    .b(_1279_),
    .s(_1201_),
    .y(_1280_)
  );
  al_mux2l _5526_ (
    .a(\DFF_603.Q ),
    .b(_1280_),
    .s(_1263_),
    .y(\DFF_603.D )
  );
  al_nand3fft _5527_ (
    .a(_0246_),
    .b(_0288_),
    .c(_1262_),
    .y(_1281_)
  );
  al_mux2l _5528_ (
    .a(\DFF_604.Q ),
    .b(_1280_),
    .s(_1281_),
    .y(\DFF_604.D )
  );
  al_nand3fft _5529_ (
    .a(_0344_),
    .b(_0288_),
    .c(_1262_),
    .y(_1282_)
  );
  al_mux2l _5530_ (
    .a(\DFF_605.Q ),
    .b(_1280_),
    .s(_1282_),
    .y(\DFF_605.D )
  );
  al_or2 _5531_ (
    .a(_1201_),
    .b(_1269_),
    .y(_1283_)
  );
  al_and2 _5532_ (
    .a(_1201_),
    .b(_1269_),
    .y(_1284_)
  );
  al_nand2ft _5533_ (
    .a(_1284_),
    .b(_1283_),
    .y(_1285_)
  );
  al_aoi21ftf _5534_ (
    .a(_1272_),
    .b(_1285_),
    .c(_1276_),
    .y(_1286_)
  );
  al_mux2l _5535_ (
    .a(\DFF_606.Q ),
    .b(_1286_),
    .s(_1263_),
    .y(\DFF_606.D )
  );
  al_mux2l _5536_ (
    .a(\DFF_607.Q ),
    .b(_1286_),
    .s(_1281_),
    .y(\DFF_607.D )
  );
  al_mux2l _5537_ (
    .a(\DFF_608.Q ),
    .b(_1286_),
    .s(_1282_),
    .y(\DFF_608.D )
  );
  al_or2ft _5538_ (
    .a(_1266_),
    .b(_1275_),
    .y(_1287_)
  );
  al_and3fft _5539_ (
    .a(_1275_),
    .b(_1284_),
    .c(_1283_),
    .y(_1288_)
  );
  al_ao21 _5540_ (
    .a(_1287_),
    .b(_1285_),
    .c(_1288_),
    .y(_1289_)
  );
  al_mux2l _5541_ (
    .a(\DFF_609.Q ),
    .b(_1289_),
    .s(_1263_),
    .y(\DFF_609.D )
  );
  al_mux2l _5542_ (
    .a(\DFF_610.Q ),
    .b(_1289_),
    .s(_1281_),
    .y(\DFF_610.D )
  );
  al_mux2l _5543_ (
    .a(\DFF_611.Q ),
    .b(_1289_),
    .s(_1282_),
    .y(\DFF_611.D )
  );
  al_nand2 _5544_ (
    .a(_1272_),
    .b(_1288_),
    .y(_1290_)
  );
  al_mux2l _5545_ (
    .a(\DFF_612.Q ),
    .b(_1290_),
    .s(_1263_),
    .y(\DFF_612.D )
  );
  al_mux2l _5546_ (
    .a(\DFF_613.Q ),
    .b(_1290_),
    .s(_1281_),
    .y(\DFF_613.D )
  );
  al_mux2l _5547_ (
    .a(\DFF_614.Q ),
    .b(_1290_),
    .s(_1282_),
    .y(\DFF_614.D )
  );
  al_nand2 _5548_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_783.D ),
    .y(_1291_)
  );
  al_nand2ft _5549_ (
    .a(\DFF_756.Q ),
    .b(\DFF_1505.Q ),
    .y(_1292_)
  );
  al_aoi21ftf _5550_ (
    .a(\DFF_757.Q ),
    .b(\DFF_1506.Q ),
    .c(_1292_),
    .y(_1293_)
  );
  al_aoi21ftf _5551_ (
    .a(\DFF_755.Q ),
    .b(\DFF_1504.Q ),
    .c(_1293_),
    .y(_1294_)
  );
  al_nand2ft _5552_ (
    .a(\DFF_758.Q ),
    .b(\DFF_1504.Q ),
    .y(_1295_)
  );
  al_aoi21ftf _5553_ (
    .a(\DFF_760.Q ),
    .b(\DFF_1506.Q ),
    .c(_1295_),
    .y(_1296_)
  );
  al_aoi21ftf _5554_ (
    .a(\DFF_759.Q ),
    .b(\DFF_1505.Q ),
    .c(_1296_),
    .y(_1297_)
  );
  al_and2ft _5555_ (
    .a(_1294_),
    .b(_1297_),
    .y(_1298_)
  );
  al_nand2ft _5556_ (
    .a(\DFF_762.Q ),
    .b(\DFF_1505.Q ),
    .y(_1299_)
  );
  al_aoi21ftf _5557_ (
    .a(\DFF_763.Q ),
    .b(\DFF_1506.Q ),
    .c(_1299_),
    .y(_1300_)
  );
  al_aoi21ftf _5558_ (
    .a(\DFF_761.Q ),
    .b(\DFF_1504.Q ),
    .c(_1300_),
    .y(_1301_)
  );
  al_nor2 _5559_ (
    .a(_1294_),
    .b(_1301_),
    .y(_1302_)
  );
  al_nand2ft _5560_ (
    .a(\DFF_765.Q ),
    .b(\DFF_1505.Q ),
    .y(_1303_)
  );
  al_aoi21ftf _5561_ (
    .a(\DFF_766.Q ),
    .b(\DFF_1506.Q ),
    .c(_1303_),
    .y(_1304_)
  );
  al_aoi21ftf _5562_ (
    .a(\DFF_764.Q ),
    .b(\DFF_1504.Q ),
    .c(_1304_),
    .y(_1305_)
  );
  al_and3fft _5563_ (
    .a(_1201_),
    .b(_1302_),
    .c(_1305_),
    .y(_1306_)
  );
  al_nand2ft _5564_ (
    .a(_1297_),
    .b(_1301_),
    .y(_1307_)
  );
  al_nand2ft _5565_ (
    .a(_1294_),
    .b(_1305_),
    .y(_1308_)
  );
  al_nand3 _5566_ (
    .a(_1201_),
    .b(_1308_),
    .c(_1307_),
    .y(_1309_)
  );
  al_ao21ftf _5567_ (
    .a(_1298_),
    .b(_1306_),
    .c(_1309_),
    .y(_1310_)
  );
  al_mux2l _5568_ (
    .a(\DFF_755.Q ),
    .b(_1310_),
    .s(_1291_),
    .y(\DFF_755.D )
  );
  al_nand2 _5569_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_783.D ),
    .y(_1311_)
  );
  al_mux2l _5570_ (
    .a(\DFF_756.Q ),
    .b(_1310_),
    .s(_1311_),
    .y(\DFF_756.D )
  );
  al_nand2 _5571_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_783.D ),
    .y(_1312_)
  );
  al_mux2l _5572_ (
    .a(\DFF_757.Q ),
    .b(_1310_),
    .s(_1312_),
    .y(\DFF_757.D )
  );
  al_or2 _5573_ (
    .a(_1201_),
    .b(_1294_),
    .y(_1313_)
  );
  al_nand2 _5574_ (
    .a(_1201_),
    .b(_1294_),
    .y(_1314_)
  );
  al_nand2 _5575_ (
    .a(_1314_),
    .b(_1313_),
    .y(_1315_)
  );
  al_aoi21ftf _5576_ (
    .a(_1301_),
    .b(_1315_),
    .c(_1307_),
    .y(_1316_)
  );
  al_mux2l _5577_ (
    .a(\DFF_758.Q ),
    .b(_1316_),
    .s(_1291_),
    .y(\DFF_758.D )
  );
  al_mux2l _5578_ (
    .a(\DFF_759.Q ),
    .b(_1316_),
    .s(_1311_),
    .y(\DFF_759.D )
  );
  al_mux2l _5579_ (
    .a(\DFF_760.Q ),
    .b(_1316_),
    .s(_1312_),
    .y(\DFF_760.D )
  );
  al_and2 _5580_ (
    .a(_1297_),
    .b(_1305_),
    .y(_1317_)
  );
  al_nand3 _5581_ (
    .a(_1297_),
    .b(_1314_),
    .c(_1313_),
    .y(_1318_)
  );
  al_ao21ftf _5582_ (
    .a(_1317_),
    .b(_1315_),
    .c(_1318_),
    .y(_1319_)
  );
  al_mux2l _5583_ (
    .a(\DFF_761.Q ),
    .b(_1319_),
    .s(_1291_),
    .y(\DFF_761.D )
  );
  al_mux2l _5584_ (
    .a(\DFF_762.Q ),
    .b(_1319_),
    .s(_1311_),
    .y(\DFF_762.D )
  );
  al_mux2l _5585_ (
    .a(\DFF_763.Q ),
    .b(_1319_),
    .s(_1312_),
    .y(\DFF_763.D )
  );
  al_nand2 _5586_ (
    .a(_1301_),
    .b(_1297_),
    .y(_1320_)
  );
  al_or3fft _5587_ (
    .a(_1314_),
    .b(_1313_),
    .c(_1320_),
    .y(_1321_)
  );
  al_mux2l _5588_ (
    .a(\DFF_764.Q ),
    .b(_1321_),
    .s(_1291_),
    .y(\DFF_764.D )
  );
  al_mux2l _5589_ (
    .a(\DFF_765.Q ),
    .b(_1321_),
    .s(_1311_),
    .y(\DFF_765.D )
  );
  al_mux2l _5590_ (
    .a(\DFF_766.Q ),
    .b(_1321_),
    .s(_1312_),
    .y(\DFF_766.D )
  );
  al_oa21ftf _5591_ (
    .a(_0048_),
    .b(_1144_),
    .c(_0035_),
    .y(_1322_)
  );
  al_aoi21ftf _5592_ (
    .a(_0048_),
    .b(_1144_),
    .c(_1322_),
    .y(\DFF_816.D )
  );
  al_and3 _5593_ (
    .a(\DFF_939.Q ),
    .b(\DFF_940.Q ),
    .c(_0937_),
    .y(_1323_)
  );
  al_aoi21 _5594_ (
    .a(\DFF_939.Q ),
    .b(_0937_),
    .c(\DFF_940.Q ),
    .y(_1324_)
  );
  al_nor3ftt _5595_ (
    .a(_0778_),
    .b(_1323_),
    .c(_1324_),
    .y(\DFF_940.D )
  );
  al_or2 _5596_ (
    .a(_0393_),
    .b(_0307_),
    .y(_1325_)
  );
  al_nand3fft _5597_ (
    .a(_1197_),
    .b(_0305_),
    .c(_1325_),
    .y(_1326_)
  );
  al_nand2ft _5598_ (
    .a(\DFF_962.Q ),
    .b(\DFF_1427.Q ),
    .y(_1327_)
  );
  al_aoi21ftf _5599_ (
    .a(\DFF_964.Q ),
    .b(\DFF_1429.Q ),
    .c(_1327_),
    .y(_1328_)
  );
  al_aoi21ftf _5600_ (
    .a(\DFF_963.Q ),
    .b(\DFF_1428.Q ),
    .c(_1328_),
    .y(_1329_)
  );
  al_nand2ft _5601_ (
    .a(\DFF_954.Q ),
    .b(\DFF_1428.Q ),
    .y(_1330_)
  );
  al_aoi21ftf _5602_ (
    .a(\DFF_955.Q ),
    .b(\DFF_1429.Q ),
    .c(_1330_),
    .y(_1331_)
  );
  al_aoi21ftf _5603_ (
    .a(\DFF_953.Q ),
    .b(\DFF_1427.Q ),
    .c(_1331_),
    .y(_1332_)
  );
  al_nand2ft _5604_ (
    .a(\DFF_960.Q ),
    .b(\DFF_1428.Q ),
    .y(_1333_)
  );
  al_aoi21ftf _5605_ (
    .a(\DFF_961.Q ),
    .b(\DFF_1429.Q ),
    .c(_1333_),
    .y(_1334_)
  );
  al_aoi21ftf _5606_ (
    .a(\DFF_959.Q ),
    .b(\DFF_1427.Q ),
    .c(_1334_),
    .y(_1335_)
  );
  al_and2ft _5607_ (
    .a(\DFF_956.Q ),
    .b(\DFF_1427.Q ),
    .y(_1336_)
  );
  al_aoi21ftt _5608_ (
    .a(\DFF_958.Q ),
    .b(\DFF_1429.Q ),
    .c(_1336_),
    .y(_1337_)
  );
  al_ao21ftf _5609_ (
    .a(\DFF_957.Q ),
    .b(\DFF_1428.Q ),
    .c(_1337_),
    .y(_1338_)
  );
  al_nand2 _5610_ (
    .a(_1335_),
    .b(_1338_),
    .y(_1339_)
  );
  al_aoi21ftf _5611_ (
    .a(_1332_),
    .b(_1329_),
    .c(_1339_),
    .y(_1340_)
  );
  al_oai21ftt _5612_ (
    .a(_1329_),
    .b(_1338_),
    .c(_1335_),
    .y(_1341_)
  );
  al_aoi21ftf _5613_ (
    .a(_1332_),
    .b(_1341_),
    .c(_1329_),
    .y(_1342_)
  );
  al_mux2l _5614_ (
    .a(_1340_),
    .b(_1342_),
    .s(_1201_),
    .y(_1343_)
  );
  al_mux2l _5615_ (
    .a(\DFF_953.Q ),
    .b(_1343_),
    .s(_1326_),
    .y(\DFF_953.D )
  );
  al_nand3fft _5616_ (
    .a(_0246_),
    .b(_0305_),
    .c(_1325_),
    .y(_1344_)
  );
  al_mux2l _5617_ (
    .a(\DFF_954.Q ),
    .b(_1343_),
    .s(_1344_),
    .y(\DFF_954.D )
  );
  al_nand3fft _5618_ (
    .a(_0344_),
    .b(_0305_),
    .c(_1325_),
    .y(_1345_)
  );
  al_mux2l _5619_ (
    .a(\DFF_955.Q ),
    .b(_1343_),
    .s(_1345_),
    .y(\DFF_955.D )
  );
  al_or2 _5620_ (
    .a(_1201_),
    .b(_1332_),
    .y(_1346_)
  );
  al_and2 _5621_ (
    .a(_1201_),
    .b(_1332_),
    .y(_1347_)
  );
  al_nand2ft _5622_ (
    .a(_1347_),
    .b(_1346_),
    .y(_1348_)
  );
  al_aoi21ftf _5623_ (
    .a(_1335_),
    .b(_1348_),
    .c(_1339_),
    .y(_1349_)
  );
  al_mux2l _5624_ (
    .a(\DFF_956.Q ),
    .b(_1349_),
    .s(_1326_),
    .y(\DFF_956.D )
  );
  al_mux2l _5625_ (
    .a(\DFF_957.Q ),
    .b(_1349_),
    .s(_1344_),
    .y(\DFF_957.D )
  );
  al_mux2l _5626_ (
    .a(\DFF_958.Q ),
    .b(_1349_),
    .s(_1345_),
    .y(\DFF_958.D )
  );
  al_or2ft _5627_ (
    .a(_1329_),
    .b(_1338_),
    .y(_1350_)
  );
  al_and3fft _5628_ (
    .a(_1338_),
    .b(_1347_),
    .c(_1346_),
    .y(_1351_)
  );
  al_ao21 _5629_ (
    .a(_1350_),
    .b(_1348_),
    .c(_1351_),
    .y(_1352_)
  );
  al_mux2l _5630_ (
    .a(\DFF_959.Q ),
    .b(_1352_),
    .s(_1326_),
    .y(\DFF_959.D )
  );
  al_mux2l _5631_ (
    .a(\DFF_960.Q ),
    .b(_1352_),
    .s(_1344_),
    .y(\DFF_960.D )
  );
  al_mux2l _5632_ (
    .a(\DFF_961.Q ),
    .b(_1352_),
    .s(_1345_),
    .y(\DFF_961.D )
  );
  al_nand2 _5633_ (
    .a(_1335_),
    .b(_1351_),
    .y(_1353_)
  );
  al_mux2l _5634_ (
    .a(\DFF_962.Q ),
    .b(_1353_),
    .s(_1326_),
    .y(\DFF_962.D )
  );
  al_mux2l _5635_ (
    .a(\DFF_963.Q ),
    .b(_1353_),
    .s(_1344_),
    .y(\DFF_963.D )
  );
  al_mux2l _5636_ (
    .a(\DFF_964.Q ),
    .b(_1353_),
    .s(_1345_),
    .y(\DFF_964.D )
  );
  al_nand2 _5637_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_1133.D ),
    .y(_1354_)
  );
  al_nand2ft _5638_ (
    .a(\DFF_1115.Q ),
    .b(\DFF_1505.Q ),
    .y(_1355_)
  );
  al_aoi21ftf _5639_ (
    .a(\DFF_1116.Q ),
    .b(\DFF_1506.Q ),
    .c(_1355_),
    .y(_1356_)
  );
  al_aoi21ftf _5640_ (
    .a(\DFF_1114.Q ),
    .b(\DFF_1504.Q ),
    .c(_1356_),
    .y(_1357_)
  );
  al_nand2ft _5641_ (
    .a(\DFF_1106.Q ),
    .b(\DFF_1505.Q ),
    .y(_1358_)
  );
  al_aoi21ftf _5642_ (
    .a(\DFF_1107.Q ),
    .b(\DFF_1506.Q ),
    .c(_1358_),
    .y(_1359_)
  );
  al_aoi21ftf _5643_ (
    .a(\DFF_1105.Q ),
    .b(\DFF_1504.Q ),
    .c(_1359_),
    .y(_1360_)
  );
  al_nand2ft _5644_ (
    .a(\DFF_1109.Q ),
    .b(\DFF_1505.Q ),
    .y(_1361_)
  );
  al_ao21ftf _5645_ (
    .a(\DFF_1110.Q ),
    .b(\DFF_1506.Q ),
    .c(_1361_),
    .y(_1362_)
  );
  al_aoi21ftt _5646_ (
    .a(\DFF_1108.Q ),
    .b(\DFF_1504.Q ),
    .c(_1362_),
    .y(_1363_)
  );
  al_oa21ftt _5647_ (
    .a(_1363_),
    .b(_1360_),
    .c(_1357_),
    .y(_1364_)
  );
  al_nand2ft _5648_ (
    .a(\DFF_1112.Q ),
    .b(\DFF_1505.Q ),
    .y(_1365_)
  );
  al_aoi21ftf _5649_ (
    .a(\DFF_1113.Q ),
    .b(\DFF_1506.Q ),
    .c(_1365_),
    .y(_1366_)
  );
  al_aoi21ftf _5650_ (
    .a(\DFF_1111.Q ),
    .b(\DFF_1504.Q ),
    .c(_1366_),
    .y(_1367_)
  );
  al_oai21ttf _5651_ (
    .a(_1360_),
    .b(_1367_),
    .c(_1201_),
    .y(_1368_)
  );
  al_nand2ft _5652_ (
    .a(_1360_),
    .b(_1357_),
    .y(_1369_)
  );
  al_nand2ft _5653_ (
    .a(_1363_),
    .b(_1367_),
    .y(_1370_)
  );
  al_nand3 _5654_ (
    .a(_1201_),
    .b(_1369_),
    .c(_1370_),
    .y(_1371_)
  );
  al_ao21ftf _5655_ (
    .a(_1368_),
    .b(_1364_),
    .c(_1371_),
    .y(_1372_)
  );
  al_mux2l _5656_ (
    .a(\DFF_1105.Q ),
    .b(_1372_),
    .s(_1354_),
    .y(\DFF_1105.D )
  );
  al_nand2 _5657_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_1133.D ),
    .y(_1373_)
  );
  al_mux2l _5658_ (
    .a(\DFF_1106.Q ),
    .b(_1372_),
    .s(_1373_),
    .y(\DFF_1106.D )
  );
  al_nand2 _5659_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_1133.D ),
    .y(_1374_)
  );
  al_mux2l _5660_ (
    .a(\DFF_1107.Q ),
    .b(_1372_),
    .s(_1374_),
    .y(\DFF_1107.D )
  );
  al_inv _5661_ (
    .a(_1367_),
    .y(_1375_)
  );
  al_nor2 _5662_ (
    .a(g3229),
    .b(_1360_),
    .y(_1376_)
  );
  al_nand2 _5663_ (
    .a(g3229),
    .b(_1360_),
    .y(_1377_)
  );
  al_or2ft _5664_ (
    .a(_1377_),
    .b(_1376_),
    .y(_1378_)
  );
  al_mux2h _5665_ (
    .a(_1363_),
    .b(_1378_),
    .s(_1375_),
    .y(_1379_)
  );
  al_mux2l _5666_ (
    .a(\DFF_1108.Q ),
    .b(_1379_),
    .s(_1354_),
    .y(\DFF_1108.D )
  );
  al_mux2l _5667_ (
    .a(\DFF_1109.Q ),
    .b(_1379_),
    .s(_1373_),
    .y(\DFF_1109.D )
  );
  al_mux2l _5668_ (
    .a(\DFF_1110.Q ),
    .b(_1379_),
    .s(_1374_),
    .y(\DFF_1110.D )
  );
  al_nand2 _5669_ (
    .a(_1357_),
    .b(_1363_),
    .y(_1380_)
  );
  al_mux2l _5670_ (
    .a(_1363_),
    .b(_1380_),
    .s(_1378_),
    .y(_1381_)
  );
  al_mux2l _5671_ (
    .a(\DFF_1111.Q ),
    .b(_1381_),
    .s(_1354_),
    .y(\DFF_1111.D )
  );
  al_mux2l _5672_ (
    .a(\DFF_1112.Q ),
    .b(_1381_),
    .s(_1373_),
    .y(\DFF_1112.D )
  );
  al_mux2l _5673_ (
    .a(\DFF_1113.Q ),
    .b(_1381_),
    .s(_1374_),
    .y(\DFF_1113.D )
  );
  al_and2 _5674_ (
    .a(_1367_),
    .b(_1363_),
    .y(_1382_)
  );
  al_oai21ftt _5675_ (
    .a(_1377_),
    .b(_1376_),
    .c(_1382_),
    .y(_1383_)
  );
  al_mux2l _5676_ (
    .a(\DFF_1114.Q ),
    .b(_1383_),
    .s(_1354_),
    .y(\DFF_1114.D )
  );
  al_mux2l _5677_ (
    .a(\DFF_1115.Q ),
    .b(_1383_),
    .s(_1373_),
    .y(\DFF_1115.D )
  );
  al_mux2l _5678_ (
    .a(\DFF_1116.Q ),
    .b(_1383_),
    .s(_1374_),
    .y(\DFF_1116.D )
  );
  al_oa21ftf _5679_ (
    .a(_0075_),
    .b(_1167_),
    .c(_0062_),
    .y(_1384_)
  );
  al_aoi21ftf _5680_ (
    .a(_0075_),
    .b(_1167_),
    .c(_1384_),
    .y(\DFF_1166.D )
  );
  al_and3 _5681_ (
    .a(\DFF_1289.Q ),
    .b(\DFF_1290.Q ),
    .c(_1014_),
    .y(_1385_)
  );
  al_aoi21 _5682_ (
    .a(\DFF_1289.Q ),
    .b(_1014_),
    .c(\DFF_1290.Q ),
    .y(_1386_)
  );
  al_nor3ftt _5683_ (
    .a(_0778_),
    .b(_1385_),
    .c(_1386_),
    .y(\DFF_1290.D )
  );
  al_and2ft _5684_ (
    .a(_0314_),
    .b(_0317_),
    .y(_1387_)
  );
  al_ao21ftt _5685_ (
    .a(_0320_),
    .b(_1387_),
    .c(_0393_),
    .y(_1388_)
  );
  al_nand3fft _5686_ (
    .a(_1197_),
    .b(_0321_),
    .c(_1388_),
    .y(_1389_)
  );
  al_nand2ft _5687_ (
    .a(\DFF_1312.Q ),
    .b(\DFF_1427.Q ),
    .y(_1390_)
  );
  al_aoi21ftf _5688_ (
    .a(\DFF_1314.Q ),
    .b(\DFF_1429.Q ),
    .c(_1390_),
    .y(_1391_)
  );
  al_aoi21ftf _5689_ (
    .a(\DFF_1313.Q ),
    .b(\DFF_1428.Q ),
    .c(_1391_),
    .y(_1392_)
  );
  al_nand2ft _5690_ (
    .a(\DFF_1304.Q ),
    .b(\DFF_1428.Q ),
    .y(_1393_)
  );
  al_aoi21ftf _5691_ (
    .a(\DFF_1305.Q ),
    .b(\DFF_1429.Q ),
    .c(_1393_),
    .y(_1394_)
  );
  al_aoi21ftf _5692_ (
    .a(\DFF_1303.Q ),
    .b(\DFF_1427.Q ),
    .c(_1394_),
    .y(_1395_)
  );
  al_nand2ft _5693_ (
    .a(\DFF_1310.Q ),
    .b(\DFF_1428.Q ),
    .y(_1396_)
  );
  al_aoi21ftf _5694_ (
    .a(\DFF_1311.Q ),
    .b(\DFF_1429.Q ),
    .c(_1396_),
    .y(_1397_)
  );
  al_aoi21ftf _5695_ (
    .a(\DFF_1309.Q ),
    .b(\DFF_1427.Q ),
    .c(_1397_),
    .y(_1398_)
  );
  al_and2ft _5696_ (
    .a(\DFF_1306.Q ),
    .b(\DFF_1427.Q ),
    .y(_1399_)
  );
  al_aoi21ftt _5697_ (
    .a(\DFF_1308.Q ),
    .b(\DFF_1429.Q ),
    .c(_1399_),
    .y(_1400_)
  );
  al_ao21ftf _5698_ (
    .a(\DFF_1307.Q ),
    .b(\DFF_1428.Q ),
    .c(_1400_),
    .y(_1401_)
  );
  al_nand2 _5699_ (
    .a(_1398_),
    .b(_1401_),
    .y(_1402_)
  );
  al_aoi21ftf _5700_ (
    .a(_1395_),
    .b(_1392_),
    .c(_1402_),
    .y(_1403_)
  );
  al_oai21ftt _5701_ (
    .a(_1392_),
    .b(_1401_),
    .c(_1398_),
    .y(_1404_)
  );
  al_aoi21ftf _5702_ (
    .a(_1395_),
    .b(_1404_),
    .c(_1392_),
    .y(_1405_)
  );
  al_mux2l _5703_ (
    .a(_1403_),
    .b(_1405_),
    .s(_1201_),
    .y(_1406_)
  );
  al_mux2l _5704_ (
    .a(\DFF_1303.Q ),
    .b(_1406_),
    .s(_1389_),
    .y(\DFF_1303.D )
  );
  al_nand3fft _5705_ (
    .a(_0246_),
    .b(_0321_),
    .c(_1388_),
    .y(_1407_)
  );
  al_mux2l _5706_ (
    .a(\DFF_1304.Q ),
    .b(_1406_),
    .s(_1407_),
    .y(\DFF_1304.D )
  );
  al_nand3fft _5707_ (
    .a(_0344_),
    .b(_0321_),
    .c(_1388_),
    .y(_1408_)
  );
  al_mux2l _5708_ (
    .a(\DFF_1305.Q ),
    .b(_1406_),
    .s(_1408_),
    .y(\DFF_1305.D )
  );
  al_or2 _5709_ (
    .a(_1201_),
    .b(_1395_),
    .y(_1409_)
  );
  al_and2 _5710_ (
    .a(_1201_),
    .b(_1395_),
    .y(_1410_)
  );
  al_nand2ft _5711_ (
    .a(_1410_),
    .b(_1409_),
    .y(_1411_)
  );
  al_aoi21ftf _5712_ (
    .a(_1398_),
    .b(_1411_),
    .c(_1402_),
    .y(_1412_)
  );
  al_mux2l _5713_ (
    .a(\DFF_1306.Q ),
    .b(_1412_),
    .s(_1389_),
    .y(\DFF_1306.D )
  );
  al_mux2l _5714_ (
    .a(\DFF_1307.Q ),
    .b(_1412_),
    .s(_1407_),
    .y(\DFF_1307.D )
  );
  al_mux2l _5715_ (
    .a(\DFF_1308.Q ),
    .b(_1412_),
    .s(_1408_),
    .y(\DFF_1308.D )
  );
  al_or2ft _5716_ (
    .a(_1392_),
    .b(_1401_),
    .y(_1413_)
  );
  al_and3fft _5717_ (
    .a(_1401_),
    .b(_1410_),
    .c(_1409_),
    .y(_1414_)
  );
  al_ao21 _5718_ (
    .a(_1413_),
    .b(_1411_),
    .c(_1414_),
    .y(_1415_)
  );
  al_mux2l _5719_ (
    .a(\DFF_1309.Q ),
    .b(_1415_),
    .s(_1389_),
    .y(\DFF_1309.D )
  );
  al_mux2l _5720_ (
    .a(\DFF_1310.Q ),
    .b(_1415_),
    .s(_1407_),
    .y(\DFF_1310.D )
  );
  al_mux2l _5721_ (
    .a(\DFF_1311.Q ),
    .b(_1415_),
    .s(_1408_),
    .y(\DFF_1311.D )
  );
  al_nand2 _5722_ (
    .a(_1398_),
    .b(_1414_),
    .y(_1416_)
  );
  al_mux2l _5723_ (
    .a(\DFF_1312.Q ),
    .b(_1416_),
    .s(_1389_),
    .y(\DFF_1312.D )
  );
  al_mux2l _5724_ (
    .a(\DFF_1313.Q ),
    .b(_1416_),
    .s(_1407_),
    .y(\DFF_1313.D )
  );
  al_mux2l _5725_ (
    .a(\DFF_1314.Q ),
    .b(_1416_),
    .s(_1408_),
    .y(\DFF_1314.D )
  );
  al_nand2 _5726_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_1483.D ),
    .y(_1417_)
  );
  al_nand2ft _5727_ (
    .a(\DFF_1456.Q ),
    .b(\DFF_1505.Q ),
    .y(_1418_)
  );
  al_aoi21ftf _5728_ (
    .a(\DFF_1457.Q ),
    .b(\DFF_1506.Q ),
    .c(_1418_),
    .y(_1419_)
  );
  al_aoi21ftf _5729_ (
    .a(\DFF_1455.Q ),
    .b(\DFF_1504.Q ),
    .c(_1419_),
    .y(_1420_)
  );
  al_nand2ft _5730_ (
    .a(\DFF_1459.Q ),
    .b(\DFF_1505.Q ),
    .y(_1421_)
  );
  al_aoi21ftf _5731_ (
    .a(\DFF_1460.Q ),
    .b(\DFF_1506.Q ),
    .c(_1421_),
    .y(_1422_)
  );
  al_aoi21ftf _5732_ (
    .a(\DFF_1458.Q ),
    .b(\DFF_1504.Q ),
    .c(_1422_),
    .y(_1423_)
  );
  al_and2ft _5733_ (
    .a(_1420_),
    .b(_1423_),
    .y(_1424_)
  );
  al_nand2ft _5734_ (
    .a(\DFF_1462.Q ),
    .b(\DFF_1505.Q ),
    .y(_1425_)
  );
  al_aoi21ftf _5735_ (
    .a(\DFF_1463.Q ),
    .b(\DFF_1506.Q ),
    .c(_1425_),
    .y(_1426_)
  );
  al_ao21ftf _5736_ (
    .a(\DFF_1461.Q ),
    .b(\DFF_1504.Q ),
    .c(_1426_),
    .y(_1427_)
  );
  al_nand2ft _5737_ (
    .a(_1420_),
    .b(_1427_),
    .y(_1428_)
  );
  al_nand2ft _5738_ (
    .a(\DFF_1465.Q ),
    .b(\DFF_1505.Q ),
    .y(_1429_)
  );
  al_aoi21ftf _5739_ (
    .a(\DFF_1466.Q ),
    .b(\DFF_1506.Q ),
    .c(_1429_),
    .y(_1430_)
  );
  al_ao21ftf _5740_ (
    .a(\DFF_1464.Q ),
    .b(\DFF_1504.Q ),
    .c(_1430_),
    .y(_1431_)
  );
  al_and3ftt _5741_ (
    .a(_1431_),
    .b(g3229),
    .c(_1428_),
    .y(_1432_)
  );
  al_or2 _5742_ (
    .a(_1427_),
    .b(_1423_),
    .y(_1433_)
  );
  al_or2 _5743_ (
    .a(_1431_),
    .b(_1420_),
    .y(_1434_)
  );
  al_nand3 _5744_ (
    .a(_1201_),
    .b(_1434_),
    .c(_1433_),
    .y(_1435_)
  );
  al_ao21ftf _5745_ (
    .a(_1424_),
    .b(_1432_),
    .c(_1435_),
    .y(_1436_)
  );
  al_mux2l _5746_ (
    .a(\DFF_1455.Q ),
    .b(_1436_),
    .s(_1417_),
    .y(\DFF_1455.D )
  );
  al_nand2 _5747_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_1483.D ),
    .y(_1437_)
  );
  al_mux2l _5748_ (
    .a(\DFF_1456.Q ),
    .b(_1436_),
    .s(_1437_),
    .y(\DFF_1456.D )
  );
  al_nand2 _5749_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_1483.D ),
    .y(_1438_)
  );
  al_mux2l _5750_ (
    .a(\DFF_1457.Q ),
    .b(_1436_),
    .s(_1438_),
    .y(\DFF_1457.D )
  );
  al_or2 _5751_ (
    .a(_1201_),
    .b(_1420_),
    .y(_1439_)
  );
  al_nand2 _5752_ (
    .a(_1201_),
    .b(_1420_),
    .y(_1440_)
  );
  al_nand2 _5753_ (
    .a(_1440_),
    .b(_1439_),
    .y(_1441_)
  );
  al_aoi21ttf _5754_ (
    .a(_1427_),
    .b(_1441_),
    .c(_1433_),
    .y(_1442_)
  );
  al_mux2l _5755_ (
    .a(\DFF_1458.Q ),
    .b(_1442_),
    .s(_1417_),
    .y(\DFF_1458.D )
  );
  al_mux2l _5756_ (
    .a(\DFF_1459.Q ),
    .b(_1442_),
    .s(_1437_),
    .y(\DFF_1459.D )
  );
  al_mux2l _5757_ (
    .a(\DFF_1460.Q ),
    .b(_1442_),
    .s(_1438_),
    .y(\DFF_1460.D )
  );
  al_nand2ft _5758_ (
    .a(_1431_),
    .b(_1423_),
    .y(_1443_)
  );
  al_mux2l _5759_ (
    .a(_1443_),
    .b(_1423_),
    .s(_1441_),
    .y(_1444_)
  );
  al_mux2l _5760_ (
    .a(\DFF_1461.Q ),
    .b(_1444_),
    .s(_1417_),
    .y(\DFF_1461.D )
  );
  al_mux2l _5761_ (
    .a(\DFF_1462.Q ),
    .b(_1444_),
    .s(_1437_),
    .y(\DFF_1462.D )
  );
  al_mux2l _5762_ (
    .a(\DFF_1463.Q ),
    .b(_1444_),
    .s(_1438_),
    .y(\DFF_1463.D )
  );
  al_nand2ft _5763_ (
    .a(_1427_),
    .b(_1423_),
    .y(_1445_)
  );
  al_or3fft _5764_ (
    .a(_1440_),
    .b(_1439_),
    .c(_1445_),
    .y(_1446_)
  );
  al_mux2l _5765_ (
    .a(\DFF_1464.Q ),
    .b(_1446_),
    .s(_1417_),
    .y(\DFF_1464.D )
  );
  al_mux2l _5766_ (
    .a(\DFF_1465.Q ),
    .b(_1446_),
    .s(_1437_),
    .y(\DFF_1465.D )
  );
  al_mux2l _5767_ (
    .a(\DFF_1466.Q ),
    .b(_1446_),
    .s(_1438_),
    .y(\DFF_1466.D )
  );
  al_oa21ftf _5768_ (
    .a(_0101_),
    .b(_1190_),
    .c(_0088_),
    .y(_1447_)
  );
  al_aoi21ftf _5769_ (
    .a(_0101_),
    .b(_1190_),
    .c(_1447_),
    .y(\DFF_1516.D )
  );
  al_inv _5770_ (
    .a(\DFF_146.Q ),
    .y(_1448_)
  );
  al_and2ft _5771_ (
    .a(g3230),
    .b(g3233),
    .y(_1449_)
  );
  al_inv _5772_ (
    .a(_1449_),
    .y(\DFF_150.D )
  );
  al_and3fft _5773_ (
    .a(\DFF_159.Q ),
    .b(\DFF_157.Q ),
    .c(\DFF_158.Q ),
    .y(_1450_)
  );
  al_or3 _5774_ (
    .a(\DFF_131.Q ),
    .b(\DFF_152.Q ),
    .c(\DFF_150.Q ),
    .y(_1451_)
  );
  al_and3fft _5775_ (
    .a(\DFF_151.Q ),
    .b(_1451_),
    .c(\DFF_156.Q ),
    .y(_1452_)
  );
  al_nand2 _5776_ (
    .a(_1450_),
    .b(_1452_),
    .y(_1453_)
  );
  al_oa21ftf _5777_ (
    .a(_1448_),
    .b(_1453_),
    .c(\DFF_150.D ),
    .y(\DFF_146.D )
  );
  al_inv _5778_ (
    .a(\DFF_146.D ),
    .y(\DFF_131.D )
  );
  al_and3 _5779_ (
    .a(\DFF_241.Q ),
    .b(\DFF_240.Q ),
    .c(_1100_),
    .y(_1454_)
  );
  al_aoi21 _5780_ (
    .a(\DFF_240.Q ),
    .b(_1100_),
    .c(\DFF_241.Q ),
    .y(_1455_)
  );
  al_nor3ftt _5781_ (
    .a(_0778_),
    .b(_1454_),
    .c(_1455_),
    .y(\DFF_241.D )
  );
  al_and3fft _5782_ (
    .a(_0174_),
    .b(_0462_),
    .c(_1108_),
    .y(_1456_)
  );
  al_and3fft _5783_ (
    .a(_1456_),
    .b(_1115_),
    .c(\DFF_1302.Q ),
    .y(_1457_)
  );
  al_ao21 _5784_ (
    .a(\DFF_1427.Q ),
    .b(_1457_),
    .c(\DFF_280.Q ),
    .y(_1458_)
  );
  al_and2ft _5785_ (
    .a(_1113_),
    .b(_1117_),
    .y(_1459_)
  );
  al_aoi21ftf _5786_ (
    .a(_1197_),
    .b(_1459_),
    .c(_1458_),
    .y(\DFF_280.D )
  );
  al_ao21 _5787_ (
    .a(\DFF_1428.Q ),
    .b(_1457_),
    .c(\DFF_281.Q ),
    .y(_1460_)
  );
  al_aoi21ftf _5788_ (
    .a(_0246_),
    .b(_1459_),
    .c(_1460_),
    .y(\DFF_281.D )
  );
  al_ao21 _5789_ (
    .a(\DFF_1429.Q ),
    .b(_1457_),
    .c(\DFF_282.Q ),
    .y(_1461_)
  );
  al_aoi21ftf _5790_ (
    .a(_0344_),
    .b(_1459_),
    .c(_1461_),
    .y(\DFF_282.D )
  );
  al_nand3fft _5791_ (
    .a(_0021_),
    .b(_0022_),
    .c(_1121_),
    .y(_1462_)
  );
  al_ao21 _5792_ (
    .a(\DFF_466.Q ),
    .b(_1121_),
    .c(\DFF_467.Q ),
    .y(_1463_)
  );
  al_and3 _5793_ (
    .a(_0463_),
    .b(_1462_),
    .c(_1463_),
    .y(\DFF_467.D )
  );
  al_nand3 _5794_ (
    .a(\DFF_591.Q ),
    .b(\DFF_590.Q ),
    .c(_1123_),
    .y(_1464_)
  );
  al_ao21 _5795_ (
    .a(\DFF_590.Q ),
    .b(_1123_),
    .c(\DFF_591.Q ),
    .y(_1465_)
  );
  al_and3 _5796_ (
    .a(_0778_),
    .b(_1464_),
    .c(_1465_),
    .y(\DFF_591.D )
  );
  al_and2ft _5797_ (
    .a(_1136_),
    .b(_1140_),
    .y(_1466_)
  );
  al_and3fft _5798_ (
    .a(_0203_),
    .b(_0540_),
    .c(_1127_),
    .y(_1467_)
  );
  al_and3fft _5799_ (
    .a(_1467_),
    .b(_1138_),
    .c(\DFF_1302.Q ),
    .y(_1468_)
  );
  al_ao21 _5800_ (
    .a(\DFF_1427.Q ),
    .b(_1468_),
    .c(\DFF_630.Q ),
    .y(_1469_)
  );
  al_aoi21ttf _5801_ (
    .a(\DFF_1427.Q ),
    .b(_1466_),
    .c(_1469_),
    .y(\DFF_630.D )
  );
  al_ao21 _5802_ (
    .a(\DFF_1428.Q ),
    .b(_1468_),
    .c(\DFF_631.Q ),
    .y(_1470_)
  );
  al_aoi21ttf _5803_ (
    .a(\DFF_1428.Q ),
    .b(_1466_),
    .c(_1470_),
    .y(\DFF_631.D )
  );
  al_ao21 _5804_ (
    .a(\DFF_1429.Q ),
    .b(_1468_),
    .c(\DFF_632.Q ),
    .y(_1471_)
  );
  al_aoi21ttf _5805_ (
    .a(\DFF_1429.Q ),
    .b(_1466_),
    .c(_1471_),
    .y(\DFF_632.D )
  );
  al_and3 _5806_ (
    .a(\DFF_816.Q ),
    .b(\DFF_817.Q ),
    .c(_1144_),
    .y(_1472_)
  );
  al_aoi21 _5807_ (
    .a(\DFF_816.Q ),
    .b(_1144_),
    .c(\DFF_817.Q ),
    .y(_1473_)
  );
  al_nor3ftt _5808_ (
    .a(_0541_),
    .b(_1472_),
    .c(_1473_),
    .y(\DFF_817.D )
  );
  al_nand3 _5809_ (
    .a(\DFF_941.Q ),
    .b(\DFF_940.Q ),
    .c(_1146_),
    .y(_1474_)
  );
  al_ao21 _5810_ (
    .a(\DFF_940.Q ),
    .b(_1146_),
    .c(\DFF_941.Q ),
    .y(_1475_)
  );
  al_and3 _5811_ (
    .a(_0778_),
    .b(_1474_),
    .c(_1475_),
    .y(\DFF_941.D )
  );
  al_and2ft _5812_ (
    .a(_1159_),
    .b(_1163_),
    .y(_1476_)
  );
  al_and3ftt _5813_ (
    .a(_0226_),
    .b(_1150_),
    .c(_0618_),
    .y(_1477_)
  );
  al_and3fft _5814_ (
    .a(_1477_),
    .b(_1161_),
    .c(\DFF_1302.Q ),
    .y(_1478_)
  );
  al_ao21 _5815_ (
    .a(\DFF_1427.Q ),
    .b(_1478_),
    .c(\DFF_980.Q ),
    .y(_1479_)
  );
  al_aoi21ttf _5816_ (
    .a(\DFF_1427.Q ),
    .b(_1476_),
    .c(_1479_),
    .y(\DFF_980.D )
  );
  al_ao21 _5817_ (
    .a(\DFF_1428.Q ),
    .b(_1478_),
    .c(\DFF_981.Q ),
    .y(_1480_)
  );
  al_aoi21ttf _5818_ (
    .a(\DFF_1428.Q ),
    .b(_1476_),
    .c(_1480_),
    .y(\DFF_981.D )
  );
  al_ao21 _5819_ (
    .a(\DFF_1429.Q ),
    .b(_1478_),
    .c(\DFF_982.Q ),
    .y(_1481_)
  );
  al_aoi21ttf _5820_ (
    .a(\DFF_1429.Q ),
    .b(_1476_),
    .c(_1481_),
    .y(\DFF_982.D )
  );
  al_nand3fft _5821_ (
    .a(_0075_),
    .b(_0076_),
    .c(_1167_),
    .y(_1482_)
  );
  al_ao21 _5822_ (
    .a(\DFF_1166.Q ),
    .b(_1167_),
    .c(\DFF_1167.Q ),
    .y(_1483_)
  );
  al_and3 _5823_ (
    .a(_0620_),
    .b(_1482_),
    .c(_1483_),
    .y(\DFF_1167.D )
  );
  al_nand3 _5824_ (
    .a(\DFF_1291.Q ),
    .b(\DFF_1290.Q ),
    .c(_1169_),
    .y(_1484_)
  );
  al_ao21 _5825_ (
    .a(\DFF_1290.Q ),
    .b(_1169_),
    .c(\DFF_1291.Q ),
    .y(_1485_)
  );
  al_and3 _5826_ (
    .a(_0778_),
    .b(_1484_),
    .c(_1485_),
    .y(\DFF_1291.D )
  );
  al_or3ftt _5827_ (
    .a(_1177_),
    .b(_0249_),
    .c(_1174_),
    .y(_1486_)
  );
  al_nand3ftt _5828_ (
    .a(_1177_),
    .b(_0249_),
    .c(_1174_),
    .y(_1487_)
  );
  al_aoi21 _5829_ (
    .a(_1487_),
    .b(_1486_),
    .c(_1102_),
    .y(_1488_)
  );
  al_ao21 _5830_ (
    .a(\DFF_1427.Q ),
    .b(_1488_),
    .c(\DFF_1330.Q ),
    .y(_1489_)
  );
  al_and2 _5831_ (
    .a(_1182_),
    .b(_1186_),
    .y(_1490_)
  );
  al_aoi21ftf _5832_ (
    .a(_1197_),
    .b(_1490_),
    .c(_1489_),
    .y(\DFF_1330.D )
  );
  al_ao21 _5833_ (
    .a(\DFF_1428.Q ),
    .b(_1488_),
    .c(\DFF_1331.Q ),
    .y(_1491_)
  );
  al_aoi21ftf _5834_ (
    .a(_0246_),
    .b(_1490_),
    .c(_1491_),
    .y(\DFF_1331.D )
  );
  al_ao21 _5835_ (
    .a(\DFF_1429.Q ),
    .b(_1488_),
    .c(\DFF_1332.Q ),
    .y(_1492_)
  );
  al_aoi21ftf _5836_ (
    .a(_0344_),
    .b(_1490_),
    .c(_1492_),
    .y(\DFF_1332.D )
  );
  al_nand3fft _5837_ (
    .a(_0101_),
    .b(_0102_),
    .c(_1190_),
    .y(_1493_)
  );
  al_ao21 _5838_ (
    .a(\DFF_1516.Q ),
    .b(_1190_),
    .c(\DFF_1517.Q ),
    .y(_1494_)
  );
  al_and3 _5839_ (
    .a(_0701_),
    .b(_1493_),
    .c(_1494_),
    .y(\DFF_1517.D )
  );
  al_inv _5840_ (
    .a(\DFF_144.Q ),
    .y(_1495_)
  );
  al_oa21ftf _5841_ (
    .a(_1495_),
    .b(_1453_),
    .c(\DFF_150.D ),
    .y(\DFF_144.D )
  );
  al_inv _5842_ (
    .a(\DFF_144.D ),
    .y(\DFF_151.D )
  );
  al_and2 _5843_ (
    .a(\DFF_242.Q ),
    .b(_1454_),
    .y(_1496_)
  );
  al_or2 _5844_ (
    .a(\DFF_242.Q ),
    .b(_1454_),
    .y(_1497_)
  );
  al_nor3fft _5845_ (
    .a(_0778_),
    .b(_1497_),
    .c(_1496_),
    .y(\DFF_242.D )
  );
  al_inv _5846_ (
    .a(_1243_),
    .y(_1498_)
  );
  al_nand2 _5847_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_338.Q ),
    .y(_1499_)
  );
  al_aoi21ttf _5848_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_340.Q ),
    .c(_1499_),
    .y(_1500_)
  );
  al_aoi21ftf _5849_ (
    .a(_0025_),
    .b(\DFF_336.Q ),
    .c(_1500_),
    .y(_1501_)
  );
  al_nand2 _5850_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_344.Q ),
    .y(_1502_)
  );
  al_nand2 _5851_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_342.Q ),
    .y(_1503_)
  );
  al_and2 _5852_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_346.Q ),
    .y(_1504_)
  );
  al_and3ftt _5853_ (
    .a(_1504_),
    .b(_1502_),
    .c(_1503_),
    .y(_1505_)
  );
  al_and2ft _5854_ (
    .a(_1505_),
    .b(_1501_),
    .y(_1506_)
  );
  al_nand3ftt _5855_ (
    .a(_1235_),
    .b(_1232_),
    .c(_1506_),
    .y(_1507_)
  );
  al_nand2 _5856_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_332.Q ),
    .y(_1508_)
  );
  al_aoi21ttf _5857_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_334.Q ),
    .c(_1508_),
    .y(_1509_)
  );
  al_aoi21ftf _5858_ (
    .a(_0025_),
    .b(\DFF_330.Q ),
    .c(_1509_),
    .y(_1510_)
  );
  al_and2ft _5859_ (
    .a(_1505_),
    .b(_1235_),
    .y(_1511_)
  );
  al_and3ftt _5860_ (
    .a(_1501_),
    .b(_1510_),
    .c(_1511_),
    .y(_1512_)
  );
  al_aoi21ftf _5861_ (
    .a(_1246_),
    .b(_1512_),
    .c(_1507_),
    .y(_1513_)
  );
  al_or3 _5862_ (
    .a(_1505_),
    .b(_1510_),
    .c(_1501_),
    .y(_1514_)
  );
  al_aoi21ftf _5863_ (
    .a(_1514_),
    .b(_1498_),
    .c(_1513_),
    .y(_1515_)
  );
  al_nand2 _5864_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_350.Q ),
    .y(_1516_)
  );
  al_aoi21ttf _5865_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_352.Q ),
    .c(_1516_),
    .y(_1517_)
  );
  al_aoi21ftf _5866_ (
    .a(_0025_),
    .b(\DFF_348.Q ),
    .c(_1517_),
    .y(_1518_)
  );
  al_nor2 _5867_ (
    .a(_1232_),
    .b(_1518_),
    .y(_1519_)
  );
  al_nor2 _5868_ (
    .a(_1501_),
    .b(_1518_),
    .y(_1520_)
  );
  al_ao21ftf _5869_ (
    .a(_1510_),
    .b(_1520_),
    .c(_1232_),
    .y(_1521_)
  );
  al_nand3fft _5870_ (
    .a(_1257_),
    .b(_1519_),
    .c(_1521_),
    .y(_1522_)
  );
  al_nor3ftt _5871_ (
    .a(_1505_),
    .b(_1232_),
    .c(_1235_),
    .y(_1523_)
  );
  al_oa21ftf _5872_ (
    .a(_1501_),
    .b(_1245_),
    .c(_1523_),
    .y(_1524_)
  );
  al_aoi21ftf _5873_ (
    .a(_1240_),
    .b(_1520_),
    .c(_1524_),
    .y(_1525_)
  );
  al_nand3ftt _5874_ (
    .a(_1239_),
    .b(_1232_),
    .c(_1501_),
    .y(_1526_)
  );
  al_and3 _5875_ (
    .a(_1505_),
    .b(_1232_),
    .c(_1243_),
    .y(_1527_)
  );
  al_aoi21ttf _5876_ (
    .a(_1235_),
    .b(_1527_),
    .c(_1526_),
    .y(_1528_)
  );
  al_mux2h _5877_ (
    .a(_1528_),
    .b(_1525_),
    .s(_1510_),
    .y(_1529_)
  );
  al_and3 _5878_ (
    .a(_1522_),
    .b(_1515_),
    .c(_1529_),
    .y(_1530_)
  );
  al_and3 _5879_ (
    .a(_1232_),
    .b(_1243_),
    .c(_1518_),
    .y(_1531_)
  );
  al_oa21ftf _5880_ (
    .a(_1501_),
    .b(_1240_),
    .c(_1531_),
    .y(_1532_)
  );
  al_nand3ftt _5881_ (
    .a(_1232_),
    .b(_1243_),
    .c(_1506_),
    .y(_1533_)
  );
  al_aoi21ftf _5882_ (
    .a(_1245_),
    .b(_1520_),
    .c(_1533_),
    .y(_1534_)
  );
  al_ao21 _5883_ (
    .a(_1532_),
    .b(_1534_),
    .c(_1510_),
    .y(_1535_)
  );
  al_oai21ftf _5884_ (
    .a(_1235_),
    .b(_1510_),
    .c(_1501_),
    .y(_1536_)
  );
  al_ao21 _5885_ (
    .a(_1510_),
    .b(_1257_),
    .c(_1536_),
    .y(_1537_)
  );
  al_mux2l _5886_ (
    .a(_1243_),
    .b(_1245_),
    .s(_1510_),
    .y(_1538_)
  );
  al_ao21ttf _5887_ (
    .a(_1538_),
    .b(_1537_),
    .c(_1505_),
    .y(_1539_)
  );
  al_inv _5888_ (
    .a(_1232_),
    .y(_1540_)
  );
  al_and3fft _5889_ (
    .a(_1239_),
    .b(_1514_),
    .c(_1232_),
    .y(_1541_)
  );
  al_ao21ftt _5890_ (
    .a(_1540_),
    .b(_1512_),
    .c(_1541_),
    .y(_1542_)
  );
  al_nand3 _5891_ (
    .a(_1510_),
    .b(_1501_),
    .c(_1236_),
    .y(_1543_)
  );
  al_ao21ftf _5892_ (
    .a(_1240_),
    .b(_1506_),
    .c(_1543_),
    .y(_1544_)
  );
  al_and2ft _5893_ (
    .a(_1243_),
    .b(_1510_),
    .y(_1545_)
  );
  al_and3ftt _5894_ (
    .a(_1239_),
    .b(_1232_),
    .c(_1518_),
    .y(_1546_)
  );
  al_aoi21 _5895_ (
    .a(_1545_),
    .b(_1519_),
    .c(_1546_),
    .y(_1547_)
  );
  al_nor3ftt _5896_ (
    .a(_1547_),
    .b(_1544_),
    .c(_1542_),
    .y(_1548_)
  );
  al_and3 _5897_ (
    .a(_1539_),
    .b(_1535_),
    .c(_1548_),
    .y(_1549_)
  );
  al_aoi21ttf _5898_ (
    .a(_0357_),
    .b(_0367_),
    .c(_0008_),
    .y(_1550_)
  );
  al_and2 _5899_ (
    .a(_1550_),
    .b(_1549_),
    .y(_1551_)
  );
  al_ao21ftf _5900_ (
    .a(_0357_),
    .b(_1530_),
    .c(_1551_),
    .y(_1552_)
  );
  al_ao21ftf _5901_ (
    .a(_0033_),
    .b(_0009_),
    .c(_1552_),
    .y(_1553_)
  );
  al_mux2h _5902_ (
    .a(\DFF_426.Q ),
    .b(_1553_),
    .s(\DFF_1504.Q ),
    .y(\DFF_426.D )
  );
  al_mux2h _5903_ (
    .a(\DFF_427.Q ),
    .b(_1553_),
    .s(\DFF_1505.Q ),
    .y(\DFF_427.D )
  );
  al_mux2h _5904_ (
    .a(\DFF_428.Q ),
    .b(_1553_),
    .s(\DFF_1506.Q ),
    .y(\DFF_428.D )
  );
  al_nor2 _5905_ (
    .a(_0028_),
    .b(_0008_),
    .y(_1554_)
  );
  al_aoi21ftf _5906_ (
    .a(_0367_),
    .b(_1549_),
    .c(_1530_),
    .y(_1555_)
  );
  al_ao21 _5907_ (
    .a(_1550_),
    .b(_1555_),
    .c(_1554_),
    .y(_1556_)
  );
  al_mux2h _5908_ (
    .a(\DFF_423.Q ),
    .b(_1556_),
    .s(\DFF_1504.Q ),
    .y(\DFF_423.D )
  );
  al_mux2h _5909_ (
    .a(\DFF_424.Q ),
    .b(_1556_),
    .s(\DFF_1505.Q ),
    .y(\DFF_424.D )
  );
  al_mux2h _5910_ (
    .a(\DFF_425.Q ),
    .b(_1556_),
    .s(\DFF_1506.Q ),
    .y(\DFF_425.D )
  );
  al_aoi21 _5911_ (
    .a(_0023_),
    .b(_1462_),
    .c(_0029_),
    .y(_1557_)
  );
  al_aoi21ftf _5912_ (
    .a(_1462_),
    .b(\DFF_468.Q ),
    .c(_1557_),
    .y(\DFF_468.D )
  );
  al_and3 _5913_ (
    .a(\DFF_591.Q ),
    .b(\DFF_592.Q ),
    .c(_1260_),
    .y(_1558_)
  );
  al_aoi21 _5914_ (
    .a(\DFF_591.Q ),
    .b(_1260_),
    .c(\DFF_592.Q ),
    .y(_1559_)
  );
  al_nor3ftt _5915_ (
    .a(_0778_),
    .b(_1558_),
    .c(_1559_),
    .y(\DFF_592.D )
  );
  al_nor2ft _5916_ (
    .a(_0059_),
    .b(_0008_),
    .y(_1560_)
  );
  al_aoi21ttf _5917_ (
    .a(_0380_),
    .b(_0390_),
    .c(_0008_),
    .y(_1561_)
  );
  al_nand2 _5918_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_694.Q ),
    .y(_1562_)
  );
  al_nand2 _5919_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_692.Q ),
    .y(_1563_)
  );
  al_and2 _5920_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_696.Q ),
    .y(_1564_)
  );
  al_and3ftt _5921_ (
    .a(_1564_),
    .b(_1562_),
    .c(_1563_),
    .y(_1565_)
  );
  al_nand2 _5922_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_688.Q ),
    .y(_1566_)
  );
  al_aoi21ttf _5923_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_690.Q ),
    .c(_1566_),
    .y(_1567_)
  );
  al_aoi21ftf _5924_ (
    .a(_0025_),
    .b(\DFF_686.Q ),
    .c(_1567_),
    .y(_1568_)
  );
  al_and2ft _5925_ (
    .a(_1565_),
    .b(_1568_),
    .y(_1569_)
  );
  al_and3ftt _5926_ (
    .a(_1297_),
    .b(_1294_),
    .c(_1569_),
    .y(_1570_)
  );
  al_nand2 _5927_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_682.Q ),
    .y(_1571_)
  );
  al_aoi21ttf _5928_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_684.Q ),
    .c(_1571_),
    .y(_1572_)
  );
  al_aoi21ftf _5929_ (
    .a(_0025_),
    .b(\DFF_680.Q ),
    .c(_1572_),
    .y(_1573_)
  );
  al_and2ft _5930_ (
    .a(_1565_),
    .b(_1573_),
    .y(_1574_)
  );
  al_nand3ftt _5931_ (
    .a(_1568_),
    .b(_1297_),
    .c(_1574_),
    .y(_1575_)
  );
  al_oa21ttf _5932_ (
    .a(_1308_),
    .b(_1575_),
    .c(_1570_),
    .y(_1576_)
  );
  al_inv _5933_ (
    .a(_1565_),
    .y(_1577_)
  );
  al_and3fft _5934_ (
    .a(_1573_),
    .b(_1568_),
    .c(_1577_),
    .y(_1578_)
  );
  al_ao21ftf _5935_ (
    .a(_1305_),
    .b(_1578_),
    .c(_1576_),
    .y(_1579_)
  );
  al_nand2 _5936_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_700.Q ),
    .y(_1580_)
  );
  al_aoi21ttf _5937_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_702.Q ),
    .c(_1580_),
    .y(_1581_)
  );
  al_ao21ftf _5938_ (
    .a(_0025_),
    .b(\DFF_698.Q ),
    .c(_1581_),
    .y(_1582_)
  );
  al_and2ft _5939_ (
    .a(_1294_),
    .b(_1582_),
    .y(_1583_)
  );
  al_nand3fft _5940_ (
    .a(_1573_),
    .b(_1568_),
    .c(_1582_),
    .y(_1584_)
  );
  al_nand2 _5941_ (
    .a(_1294_),
    .b(_1584_),
    .y(_1585_)
  );
  al_nand3fft _5942_ (
    .a(_1320_),
    .b(_1583_),
    .c(_1585_),
    .y(_1586_)
  );
  al_nor3ftt _5943_ (
    .a(_1565_),
    .b(_1294_),
    .c(_1297_),
    .y(_1587_)
  );
  al_oai21ftt _5944_ (
    .a(_1301_),
    .b(_1297_),
    .c(_1568_),
    .y(_1588_)
  );
  al_ao21 _5945_ (
    .a(_1582_),
    .b(_1302_),
    .c(_1568_),
    .y(_1589_)
  );
  al_ao21 _5946_ (
    .a(_1588_),
    .b(_1589_),
    .c(_1587_),
    .y(_1590_)
  );
  al_nand3ftt _5947_ (
    .a(_1301_),
    .b(_1294_),
    .c(_1568_),
    .y(_1591_)
  );
  al_and3 _5948_ (
    .a(_1565_),
    .b(_1294_),
    .c(_1305_),
    .y(_1592_)
  );
  al_ao21ttf _5949_ (
    .a(_1297_),
    .b(_1592_),
    .c(_1591_),
    .y(_1593_)
  );
  al_mux2h _5950_ (
    .a(_1593_),
    .b(_1590_),
    .s(_1573_),
    .y(_1594_)
  );
  al_and3fft _5951_ (
    .a(_1579_),
    .b(_1594_),
    .c(_1586_),
    .y(_1595_)
  );
  al_or3ftt _5952_ (
    .a(_1305_),
    .b(_1294_),
    .c(_1573_),
    .y(_1596_)
  );
  al_oa21ftt _5953_ (
    .a(_1596_),
    .b(_1302_),
    .c(_1569_),
    .y(_1597_)
  );
  al_nand3fft _5954_ (
    .a(_1294_),
    .b(_1301_),
    .c(_1568_),
    .y(_1598_)
  );
  al_nand3ftt _5955_ (
    .a(_1582_),
    .b(_1294_),
    .c(_1305_),
    .y(_1599_)
  );
  al_aoi21 _5956_ (
    .a(_1598_),
    .b(_1599_),
    .c(_1573_),
    .y(_1600_)
  );
  al_nand3 _5957_ (
    .a(_1573_),
    .b(_1568_),
    .c(_1298_),
    .y(_1601_)
  );
  al_and3ftt _5958_ (
    .a(_1305_),
    .b(_1573_),
    .c(_1583_),
    .y(_1602_)
  );
  al_aoi21ftf _5959_ (
    .a(_0025_),
    .b(\DFF_698.Q ),
    .c(_1581_),
    .y(_1603_)
  );
  al_nand3ftt _5960_ (
    .a(_1301_),
    .b(_1294_),
    .c(_1603_),
    .y(_1604_)
  );
  al_nor3fft _5961_ (
    .a(_1604_),
    .b(_1601_),
    .c(_1602_),
    .y(_1605_)
  );
  al_nand3fft _5962_ (
    .a(_1597_),
    .b(_1600_),
    .c(_1605_),
    .y(_1606_)
  );
  al_and2ft _5963_ (
    .a(_1305_),
    .b(_1573_),
    .y(_1607_)
  );
  al_mux2h _5964_ (
    .a(_1297_),
    .b(_1320_),
    .s(_1573_),
    .y(_1608_)
  );
  al_oai21ftf _5965_ (
    .a(_1588_),
    .b(_1608_),
    .c(_1607_),
    .y(_1609_)
  );
  al_and2 _5966_ (
    .a(_1565_),
    .b(_1609_),
    .y(_1610_)
  );
  al_and3fft _5967_ (
    .a(_1297_),
    .b(_1584_),
    .c(_1301_),
    .y(_1611_)
  );
  al_ao21ftf _5968_ (
    .a(_1301_),
    .b(_1578_),
    .c(_1575_),
    .y(_1612_)
  );
  al_aoi21 _5969_ (
    .a(_1294_),
    .b(_1612_),
    .c(_1611_),
    .y(_1613_)
  );
  al_and3fft _5970_ (
    .a(_1606_),
    .b(_1610_),
    .c(_1613_),
    .y(_1614_)
  );
  al_aoi21ftf _5971_ (
    .a(_0380_),
    .b(_1595_),
    .c(_1614_),
    .y(_1615_)
  );
  al_ao21 _5972_ (
    .a(_1561_),
    .b(_1615_),
    .c(_1560_),
    .y(_1616_)
  );
  al_mux2h _5973_ (
    .a(\DFF_776.Q ),
    .b(_1616_),
    .s(\DFF_1504.Q ),
    .y(\DFF_776.D )
  );
  al_mux2h _5974_ (
    .a(\DFF_777.Q ),
    .b(_1616_),
    .s(\DFF_1505.Q ),
    .y(\DFF_777.D )
  );
  al_mux2h _5975_ (
    .a(\DFF_778.Q ),
    .b(_1616_),
    .s(\DFF_1506.Q ),
    .y(\DFF_778.D )
  );
  al_nor2ft _5976_ (
    .a(_0054_),
    .b(_0008_),
    .y(_1617_)
  );
  al_aoi21ftf _5977_ (
    .a(_0390_),
    .b(_1614_),
    .c(_1595_),
    .y(_1618_)
  );
  al_ao21 _5978_ (
    .a(_1561_),
    .b(_1618_),
    .c(_1617_),
    .y(_1619_)
  );
  al_mux2h _5979_ (
    .a(\DFF_773.Q ),
    .b(_1619_),
    .s(\DFF_1504.Q ),
    .y(\DFF_773.D )
  );
  al_mux2h _5980_ (
    .a(\DFF_774.Q ),
    .b(_1619_),
    .s(\DFF_1505.Q ),
    .y(\DFF_774.D )
  );
  al_mux2h _5981_ (
    .a(\DFF_775.Q ),
    .b(_1619_),
    .s(\DFF_1506.Q ),
    .y(\DFF_775.D )
  );
  al_oa21ftf _5982_ (
    .a(_0050_),
    .b(_1472_),
    .c(_0035_),
    .y(_1620_)
  );
  al_aoi21ftf _5983_ (
    .a(_0050_),
    .b(_1472_),
    .c(_1620_),
    .y(\DFF_818.D )
  );
  al_and3 _5984_ (
    .a(\DFF_941.Q ),
    .b(\DFF_942.Q ),
    .c(_1323_),
    .y(_1621_)
  );
  al_aoi21 _5985_ (
    .a(\DFF_941.Q ),
    .b(_1323_),
    .c(\DFF_942.Q ),
    .y(_1622_)
  );
  al_nor3ftt _5986_ (
    .a(_0778_),
    .b(_1621_),
    .c(_1622_),
    .y(\DFF_942.D )
  );
  al_nor2 _5987_ (
    .a(_0086_),
    .b(_0008_),
    .y(_1623_)
  );
  al_nand2 _5988_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_1044.Q ),
    .y(_1624_)
  );
  al_aoi21ttf _5989_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_1046.Q ),
    .c(_1624_),
    .y(_1625_)
  );
  al_ao21ftf _5990_ (
    .a(_0025_),
    .b(\DFF_1042.Q ),
    .c(_1625_),
    .y(_1626_)
  );
  al_nand2 _5991_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_1032.Q ),
    .y(_1627_)
  );
  al_aoi21ttf _5992_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_1034.Q ),
    .c(_1627_),
    .y(_1628_)
  );
  al_aoi21ftf _5993_ (
    .a(_0025_),
    .b(\DFF_1030.Q ),
    .c(_1628_),
    .y(_1629_)
  );
  al_nand2 _5994_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_1038.Q ),
    .y(_1630_)
  );
  al_nand2 _5995_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_1036.Q ),
    .y(_1631_)
  );
  al_and2 _5996_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_1040.Q ),
    .y(_1632_)
  );
  al_and3ftt _5997_ (
    .a(_1632_),
    .b(_1630_),
    .c(_1631_),
    .y(_1633_)
  );
  al_oai21ftf _5998_ (
    .a(_1363_),
    .b(_1629_),
    .c(_1633_),
    .y(_1634_)
  );
  al_oai21ftf _5999_ (
    .a(_1629_),
    .b(_1382_),
    .c(_1634_),
    .y(_1635_)
  );
  al_mux2l _6000_ (
    .a(_1357_),
    .b(_1370_),
    .s(_1629_),
    .y(_1636_)
  );
  al_ao21 _6001_ (
    .a(_1636_),
    .b(_1635_),
    .c(_1626_),
    .y(_1637_)
  );
  al_nand2 _6002_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_1050.Q ),
    .y(_1638_)
  );
  al_aoi21ttf _6003_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_1052.Q ),
    .c(_1638_),
    .y(_1639_)
  );
  al_ao21ftf _6004_ (
    .a(_0025_),
    .b(\DFF_1048.Q ),
    .c(_1639_),
    .y(_1640_)
  );
  al_and3fft _6005_ (
    .a(_1367_),
    .b(_1640_),
    .c(_1360_),
    .y(_1641_)
  );
  al_and2 _6006_ (
    .a(_1633_),
    .b(_1626_),
    .y(_1642_)
  );
  al_or3ftt _6007_ (
    .a(_1642_),
    .b(_1629_),
    .c(_1369_),
    .y(_1643_)
  );
  al_nand3ftt _6008_ (
    .a(_1640_),
    .b(_1357_),
    .c(_1360_),
    .y(_1644_)
  );
  al_or3ftt _6009_ (
    .a(_1633_),
    .b(_1360_),
    .c(_1367_),
    .y(_1645_)
  );
  al_ao21 _6010_ (
    .a(_1645_),
    .b(_1644_),
    .c(_1629_),
    .y(_1646_)
  );
  al_inv _6011_ (
    .a(_1633_),
    .y(_1647_)
  );
  al_and2 _6012_ (
    .a(_1363_),
    .b(_1629_),
    .y(_1648_)
  );
  al_nand3fft _6013_ (
    .a(_1360_),
    .b(_1647_),
    .c(_1648_),
    .y(_1649_)
  );
  al_nor2 _6014_ (
    .a(_1360_),
    .b(_1367_),
    .y(_1650_)
  );
  al_nand2ft _6015_ (
    .a(_1360_),
    .b(_1640_),
    .y(_1651_)
  );
  al_and3fft _6016_ (
    .a(_1357_),
    .b(_1651_),
    .c(_1629_),
    .y(_1652_)
  );
  al_aoi21 _6017_ (
    .a(_1650_),
    .b(_1642_),
    .c(_1652_),
    .y(_1653_)
  );
  al_and3 _6018_ (
    .a(_1646_),
    .b(_1649_),
    .c(_1653_),
    .y(_1654_)
  );
  al_and3ftt _6019_ (
    .a(_1641_),
    .b(_1643_),
    .c(_1654_),
    .y(_1655_)
  );
  al_nand3 _6020_ (
    .a(_1626_),
    .b(_1647_),
    .c(_1648_),
    .y(_1656_)
  );
  al_and3fft _6021_ (
    .a(_1633_),
    .b(_1629_),
    .c(_1626_),
    .y(_1657_)
  );
  al_ao21ftf _6022_ (
    .a(_1367_),
    .b(_1657_),
    .c(_1656_),
    .y(_1658_)
  );
  al_and2ft _6023_ (
    .a(_1633_),
    .b(_1640_),
    .y(_1659_)
  );
  al_or3ftt _6024_ (
    .a(_1659_),
    .b(_1629_),
    .c(_1370_),
    .y(_1660_)
  );
  al_aoi21ttf _6025_ (
    .a(_1360_),
    .b(_1658_),
    .c(_1660_),
    .y(_1661_)
  );
  al_and3 _6026_ (
    .a(_1637_),
    .b(_1661_),
    .c(_1655_),
    .y(_1662_)
  );
  al_and3ftt _6027_ (
    .a(_1363_),
    .b(_1360_),
    .c(_1642_),
    .y(_1663_)
  );
  al_oa21ttf _6028_ (
    .a(_1369_),
    .b(_1656_),
    .c(_1663_),
    .y(_1664_)
  );
  al_aoi21ftf _6029_ (
    .a(_1357_),
    .b(_1657_),
    .c(_1664_),
    .y(_1665_)
  );
  al_ao21ftf _6030_ (
    .a(_1629_),
    .b(_1659_),
    .c(_1360_),
    .y(_1666_)
  );
  al_nand3 _6031_ (
    .a(_1382_),
    .b(_1651_),
    .c(_1666_),
    .y(_1667_)
  );
  al_or3 _6032_ (
    .a(_1360_),
    .b(_1363_),
    .c(_1626_),
    .y(_1668_)
  );
  al_aoi21ttf _6033_ (
    .a(_1659_),
    .b(_1650_),
    .c(_1668_),
    .y(_1669_)
  );
  al_aoi21ftf _6034_ (
    .a(_1370_),
    .b(_1633_),
    .c(_1669_),
    .y(_1670_)
  );
  al_or3fft _6035_ (
    .a(_1633_),
    .b(_1360_),
    .c(_1367_),
    .y(_1671_)
  );
  al_and3ftt _6036_ (
    .a(_1626_),
    .b(_1357_),
    .c(_1360_),
    .y(_1672_)
  );
  al_aoi21ttf _6037_ (
    .a(_1363_),
    .b(_1672_),
    .c(_1671_),
    .y(_1673_)
  );
  al_mux2h _6038_ (
    .a(_1673_),
    .b(_1670_),
    .s(_1629_),
    .y(_1674_)
  );
  al_and3 _6039_ (
    .a(_1667_),
    .b(_1665_),
    .c(_1674_),
    .y(_1675_)
  );
  al_aoi21ttf _6040_ (
    .a(_0404_),
    .b(_0414_),
    .c(_0008_),
    .y(_1676_)
  );
  al_aoi21ftf _6041_ (
    .a(_0404_),
    .b(_1675_),
    .c(_1676_),
    .y(_1677_)
  );
  al_ao21 _6042_ (
    .a(_1662_),
    .b(_1677_),
    .c(_1623_),
    .y(_1678_)
  );
  al_mux2h _6043_ (
    .a(\DFF_1126.Q ),
    .b(_1678_),
    .s(\DFF_1504.Q ),
    .y(\DFF_1126.D )
  );
  al_mux2h _6044_ (
    .a(\DFF_1127.Q ),
    .b(_1678_),
    .s(\DFF_1505.Q ),
    .y(\DFF_1127.D )
  );
  al_mux2h _6045_ (
    .a(\DFF_1128.Q ),
    .b(_1678_),
    .s(\DFF_1506.Q ),
    .y(\DFF_1128.D )
  );
  al_and2 _6046_ (
    .a(_1676_),
    .b(_1675_),
    .y(_1679_)
  );
  al_ao21ftf _6047_ (
    .a(_0414_),
    .b(_1662_),
    .c(_1679_),
    .y(_1680_)
  );
  al_ao21ftf _6048_ (
    .a(_0082_),
    .b(_0009_),
    .c(_1680_),
    .y(_1681_)
  );
  al_mux2h _6049_ (
    .a(\DFF_1123.Q ),
    .b(_1681_),
    .s(\DFF_1504.Q ),
    .y(\DFF_1123.D )
  );
  al_mux2h _6050_ (
    .a(\DFF_1124.Q ),
    .b(_1681_),
    .s(\DFF_1505.Q ),
    .y(\DFF_1124.D )
  );
  al_mux2h _6051_ (
    .a(\DFF_1125.Q ),
    .b(_1681_),
    .s(\DFF_1506.Q ),
    .y(\DFF_1125.D )
  );
  al_aoi21 _6052_ (
    .a(_0077_),
    .b(_1482_),
    .c(_0062_),
    .y(_1682_)
  );
  al_aoi21ftf _6053_ (
    .a(_1482_),
    .b(\DFF_1168.Q ),
    .c(_1682_),
    .y(\DFF_1168.D )
  );
  al_and3 _6054_ (
    .a(\DFF_1291.Q ),
    .b(\DFF_1292.Q ),
    .c(_1385_),
    .y(_1683_)
  );
  al_aoi21 _6055_ (
    .a(\DFF_1291.Q ),
    .b(_1385_),
    .c(\DFF_1292.Q ),
    .y(_1684_)
  );
  al_nor3ftt _6056_ (
    .a(_0778_),
    .b(_1683_),
    .c(_1684_),
    .y(\DFF_1292.D )
  );
  al_nor2 _6057_ (
    .a(_0111_),
    .b(_0008_),
    .y(_1685_)
  );
  al_nand2 _6058_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_1382.Q ),
    .y(_1686_)
  );
  al_aoi21ttf _6059_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_1384.Q ),
    .c(_1686_),
    .y(_1687_)
  );
  al_aoi21ftf _6060_ (
    .a(_0025_),
    .b(\DFF_1380.Q ),
    .c(_1687_),
    .y(_1688_)
  );
  al_nand2 _6061_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_1400.Q ),
    .y(_1689_)
  );
  al_aoi21ttf _6062_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_1402.Q ),
    .c(_1689_),
    .y(_1690_)
  );
  al_aoi21ftf _6063_ (
    .a(_0025_),
    .b(\DFF_1398.Q ),
    .c(_1690_),
    .y(_1691_)
  );
  al_nand3ftt _6064_ (
    .a(_1431_),
    .b(_1420_),
    .c(_1691_),
    .y(_1692_)
  );
  al_nand2 _6065_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_1394.Q ),
    .y(_1693_)
  );
  al_nand2 _6066_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_1392.Q ),
    .y(_1694_)
  );
  al_and2 _6067_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_1396.Q ),
    .y(_1695_)
  );
  al_and3ftt _6068_ (
    .a(_1695_),
    .b(_1693_),
    .c(_1694_),
    .y(_1696_)
  );
  al_nand2 _6069_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_1388.Q ),
    .y(_1697_)
  );
  al_aoi21ttf _6070_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_1390.Q ),
    .c(_1697_),
    .y(_1698_)
  );
  al_aoi21ftf _6071_ (
    .a(_0025_),
    .b(\DFF_1386.Q ),
    .c(_1698_),
    .y(_1699_)
  );
  al_nand2ft _6072_ (
    .a(_1696_),
    .b(_1699_),
    .y(_1700_)
  );
  al_or3 _6073_ (
    .a(_1420_),
    .b(_1431_),
    .c(_1700_),
    .y(_1701_)
  );
  al_ao21 _6074_ (
    .a(_1692_),
    .b(_1701_),
    .c(_1688_),
    .y(_1702_)
  );
  al_or2 _6075_ (
    .a(_1696_),
    .b(_1699_),
    .y(_1703_)
  );
  al_nor3fft _6076_ (
    .a(_1423_),
    .b(_1688_),
    .c(_1703_),
    .y(_1704_)
  );
  al_nand3 _6077_ (
    .a(_1427_),
    .b(_1420_),
    .c(_1691_),
    .y(_1705_)
  );
  al_aoi21ttf _6078_ (
    .a(_1420_),
    .b(_1704_),
    .c(_1705_),
    .y(_1706_)
  );
  al_or2 _6079_ (
    .a(_1420_),
    .b(_1691_),
    .y(_1707_)
  );
  al_or3fft _6080_ (
    .a(_1431_),
    .b(_1688_),
    .c(_1707_),
    .y(_1708_)
  );
  al_and3 _6081_ (
    .a(_1708_),
    .b(_1702_),
    .c(_1706_),
    .y(_1709_)
  );
  al_or3 _6082_ (
    .a(_1427_),
    .b(_1423_),
    .c(_1688_),
    .y(_1710_)
  );
  al_inv _6083_ (
    .a(_1688_),
    .y(_1711_)
  );
  al_oa21ftf _6084_ (
    .a(_1423_),
    .b(_1688_),
    .c(_1699_),
    .y(_1712_)
  );
  al_ao21ttf _6085_ (
    .a(_1688_),
    .b(_1445_),
    .c(_1712_),
    .y(_1713_)
  );
  al_aoi21ftf _6086_ (
    .a(_1711_),
    .b(_1431_),
    .c(_1713_),
    .y(_1714_)
  );
  al_ao21ttf _6087_ (
    .a(_1710_),
    .b(_1714_),
    .c(_1696_),
    .y(_1715_)
  );
  al_or3 _6088_ (
    .a(_1699_),
    .b(_1688_),
    .c(_1691_),
    .y(_1716_)
  );
  al_or3 _6089_ (
    .a(_1696_),
    .b(_1699_),
    .c(_1688_),
    .y(_1717_)
  );
  al_or3fft _6090_ (
    .a(_1420_),
    .b(_1427_),
    .c(_1717_),
    .y(_1718_)
  );
  al_oa21 _6091_ (
    .a(_1433_),
    .b(_1716_),
    .c(_1718_),
    .y(_1719_)
  );
  al_nand2ft _6092_ (
    .a(_1688_),
    .b(_1699_),
    .y(_1720_)
  );
  al_ao21 _6093_ (
    .a(_1700_),
    .b(_1720_),
    .c(_1428_),
    .y(_1721_)
  );
  al_nand3 _6094_ (
    .a(_1699_),
    .b(_1688_),
    .c(_1424_),
    .y(_1722_)
  );
  al_nand3 _6095_ (
    .a(_1722_),
    .b(_1721_),
    .c(_1719_),
    .y(_1723_)
  );
  al_and3ftt _6096_ (
    .a(_1723_),
    .b(_1709_),
    .c(_1715_),
    .y(_1724_)
  );
  al_or2ft _6097_ (
    .a(_1431_),
    .b(_1717_),
    .y(_1725_)
  );
  al_aoi21ftf _6098_ (
    .a(_1434_),
    .b(_1704_),
    .c(_1725_),
    .y(_1726_)
  );
  al_aoi21 _6099_ (
    .a(_1420_),
    .b(_1716_),
    .c(_1445_),
    .y(_1727_)
  );
  al_and3fft _6100_ (
    .a(_1423_),
    .b(_1700_),
    .c(_1420_),
    .y(_1728_)
  );
  al_aoi21 _6101_ (
    .a(_1707_),
    .b(_1727_),
    .c(_1728_),
    .y(_1729_)
  );
  al_nor3fft _6102_ (
    .a(_1696_),
    .b(_1420_),
    .c(_1431_),
    .y(_1730_)
  );
  al_nand3ftt _6103_ (
    .a(_1688_),
    .b(_1423_),
    .c(_1730_),
    .y(_1731_)
  );
  al_or3 _6104_ (
    .a(_1699_),
    .b(_1691_),
    .c(_1428_),
    .y(_1732_)
  );
  al_or3ftt _6105_ (
    .a(_1696_),
    .b(_1420_),
    .c(_1423_),
    .y(_1733_)
  );
  al_ao21 _6106_ (
    .a(_1733_),
    .b(_1732_),
    .c(_1711_),
    .y(_1734_)
  );
  al_or3fft _6107_ (
    .a(_1699_),
    .b(_1688_),
    .c(_1433_),
    .y(_1735_)
  );
  al_and2 _6108_ (
    .a(_1427_),
    .b(_1420_),
    .y(_1736_)
  );
  al_aoi21ftf _6109_ (
    .a(_1720_),
    .b(_1736_),
    .c(_1735_),
    .y(_1737_)
  );
  al_and3 _6110_ (
    .a(_1731_),
    .b(_1737_),
    .c(_1734_),
    .y(_1738_)
  );
  al_and3 _6111_ (
    .a(_1726_),
    .b(_1729_),
    .c(_1738_),
    .y(_1739_)
  );
  al_aoi21ttf _6112_ (
    .a(_0427_),
    .b(_0437_),
    .c(_0008_),
    .y(_1740_)
  );
  al_aoi21ftf _6113_ (
    .a(_0427_),
    .b(_1739_),
    .c(_1740_),
    .y(_1741_)
  );
  al_ao21 _6114_ (
    .a(_1724_),
    .b(_1741_),
    .c(_1685_),
    .y(_1742_)
  );
  al_mux2h _6115_ (
    .a(\DFF_1476.Q ),
    .b(_1742_),
    .s(\DFF_1504.Q ),
    .y(\DFF_1476.D )
  );
  al_mux2h _6116_ (
    .a(\DFF_1477.Q ),
    .b(_1742_),
    .s(\DFF_1505.Q ),
    .y(\DFF_1477.D )
  );
  al_mux2h _6117_ (
    .a(\DFF_1478.Q ),
    .b(_1742_),
    .s(\DFF_1506.Q ),
    .y(\DFF_1478.D )
  );
  al_nor2 _6118_ (
    .a(_0107_),
    .b(_0008_),
    .y(_1743_)
  );
  al_aoi21ftf _6119_ (
    .a(_0437_),
    .b(_1724_),
    .c(_1739_),
    .y(_1744_)
  );
  al_ao21 _6120_ (
    .a(_1740_),
    .b(_1744_),
    .c(_1743_),
    .y(_1745_)
  );
  al_mux2h _6121_ (
    .a(\DFF_1473.Q ),
    .b(_1745_),
    .s(\DFF_1504.Q ),
    .y(\DFF_1473.D )
  );
  al_mux2h _6122_ (
    .a(\DFF_1474.Q ),
    .b(_1745_),
    .s(\DFF_1505.Q ),
    .y(\DFF_1474.D )
  );
  al_mux2h _6123_ (
    .a(\DFF_1475.Q ),
    .b(_1745_),
    .s(\DFF_1506.Q ),
    .y(\DFF_1475.D )
  );
  al_aoi21 _6124_ (
    .a(_0103_),
    .b(_1493_),
    .c(_0088_),
    .y(_1746_)
  );
  al_aoi21ftf _6125_ (
    .a(_1493_),
    .b(\DFF_1518.Q ),
    .c(_1746_),
    .y(\DFF_1518.D )
  );
  al_mux2h _6126_ (
    .a(\DFF_110.Q ),
    .b(\DFF_750.D ),
    .s(\DFF_1504.Q ),
    .y(\DFF_110.D )
  );
  al_mux2h _6127_ (
    .a(\DFF_111.Q ),
    .b(\DFF_750.D ),
    .s(\DFF_1505.Q ),
    .y(\DFF_111.D )
  );
  al_mux2h _6128_ (
    .a(\DFF_112.Q ),
    .b(\DFF_750.D ),
    .s(\DFF_1506.Q ),
    .y(\DFF_112.D )
  );
  al_and3fft _6129_ (
    .a(\DFF_156.Q ),
    .b(_1451_),
    .c(\DFF_151.Q ),
    .y(_1747_)
  );
  al_or3 _6130_ (
    .a(\DFF_158.Q ),
    .b(\DFF_159.Q ),
    .c(\DFF_157.Q ),
    .y(_1748_)
  );
  al_nand3ftt _6131_ (
    .a(_1748_),
    .b(\DFF_107.Q ),
    .c(_1747_),
    .y(_1749_)
  );
  al_or3 _6132_ (
    .a(\DFF_151.Q ),
    .b(\DFF_156.Q ),
    .c(_1451_),
    .y(_1750_)
  );
  al_nor2 _6133_ (
    .a(\DFF_158.Q ),
    .b(\DFF_159.Q ),
    .y(_1751_)
  );
  al_and3fft _6134_ (
    .a(\DFF_157.Q ),
    .b(_1750_),
    .c(_1751_),
    .y(_1752_)
  );
  al_oai21 _6135_ (
    .a(\DFF_1624.Q ),
    .b(\DFF_1634.Q ),
    .c(_1752_),
    .y(_1753_)
  );
  al_oa21 _6136_ (
    .a(\DFF_141.Q ),
    .b(_1453_),
    .c(_1753_),
    .y(_1754_)
  );
  al_and2 _6137_ (
    .a(_1450_),
    .b(_1747_),
    .y(_1755_)
  );
  al_and3fft _6138_ (
    .a(\DFF_158.Q ),
    .b(\DFF_159.Q ),
    .c(\DFF_157.Q ),
    .y(_1756_)
  );
  al_nand3 _6139_ (
    .a(\DFF_108.Q ),
    .b(_1756_),
    .c(_1747_),
    .y(_1757_)
  );
  al_aoi21ttf _6140_ (
    .a(\DFF_109.Q ),
    .b(_1755_),
    .c(_1757_),
    .y(_1758_)
  );
  al_and3 _6141_ (
    .a(_1749_),
    .b(_1758_),
    .c(_1754_),
    .y(_1759_)
  );
  al_nand2ft _6142_ (
    .a(\DFF_157.Q ),
    .b(\DFF_159.Q ),
    .y(_1760_)
  );
  al_and2ft _6143_ (
    .a(_1760_),
    .b(_1452_),
    .y(_1761_)
  );
  al_and3fft _6144_ (
    .a(\DFF_158.Q ),
    .b(\DFF_157.Q ),
    .c(\DFF_159.Q ),
    .y(_1762_)
  );
  al_and3 _6145_ (
    .a(\DFF_111.Q ),
    .b(_1762_),
    .c(_1747_),
    .y(_1763_)
  );
  al_and3ftt _6146_ (
    .a(\DFF_158.Q ),
    .b(\DFF_159.Q ),
    .c(\DFF_157.Q ),
    .y(_1764_)
  );
  al_nand3 _6147_ (
    .a(\DFF_112.Q ),
    .b(_1764_),
    .c(_1747_),
    .y(_1765_)
  );
  al_nand3fft _6148_ (
    .a(_1761_),
    .b(_1763_),
    .c(_1765_),
    .y(_1766_)
  );
  al_and3ftt _6149_ (
    .a(_1760_),
    .b(\DFF_158.Q ),
    .c(_1747_),
    .y(_1767_)
  );
  al_ao21ttf _6150_ (
    .a(\DFF_113.Q ),
    .b(_1767_),
    .c(_1449_),
    .y(_1768_)
  );
  al_nor3fft _6151_ (
    .a(\DFF_151.Q ),
    .b(\DFF_156.Q ),
    .c(_1451_),
    .y(_1769_)
  );
  al_nand3 _6152_ (
    .a(\DFF_116.Q ),
    .b(_1756_),
    .c(_1769_),
    .y(_1770_)
  );
  al_aoi21ftf _6153_ (
    .a(_1750_),
    .b(_1762_),
    .c(_1770_),
    .y(_1771_)
  );
  al_or3ftt _6154_ (
    .a(_1771_),
    .b(_1768_),
    .c(_1766_),
    .y(_1772_)
  );
  al_and3ftt _6155_ (
    .a(\DFF_159.Q ),
    .b(\DFF_158.Q ),
    .c(\DFF_157.Q ),
    .y(_1773_)
  );
  al_nand3 _6156_ (
    .a(\DFF_118.Q ),
    .b(_1773_),
    .c(_1769_),
    .y(_1774_)
  );
  al_nand3ftt _6157_ (
    .a(_1748_),
    .b(\DFF_115.Q ),
    .c(_1769_),
    .y(_1775_)
  );
  al_nand3 _6158_ (
    .a(\DFF_117.Q ),
    .b(_1450_),
    .c(_1769_),
    .y(_1776_)
  );
  al_and3 _6159_ (
    .a(\DFF_158.Q ),
    .b(\DFF_159.Q ),
    .c(\DFF_157.Q ),
    .y(_1777_)
  );
  al_nand3 _6160_ (
    .a(\DFF_114.Q ),
    .b(_1777_),
    .c(_1747_),
    .y(_1778_)
  );
  al_and3 _6161_ (
    .a(\DFF_110.Q ),
    .b(_1773_),
    .c(_1747_),
    .y(_1779_)
  );
  al_and3ftt _6162_ (
    .a(_1779_),
    .b(_1776_),
    .c(_1778_),
    .y(_1780_)
  );
  al_and3 _6163_ (
    .a(_1774_),
    .b(_1775_),
    .c(_1780_),
    .y(_1781_)
  );
  al_and3ftt _6164_ (
    .a(_1772_),
    .b(_1781_),
    .c(_1759_),
    .y(\DFF_141.D )
  );
  al_inv _6165_ (
    .a(\DFF_141.D ),
    .y(\DFF_159.D )
  );
  al_inv _6166_ (
    .a(\DFF_243.Q ),
    .y(_1782_)
  );
  al_inv _6167_ (
    .a(\DFF_242.Q ),
    .y(_1783_)
  );
  al_nand3fft _6168_ (
    .a(_1782_),
    .b(_1783_),
    .c(_1454_),
    .y(_1784_)
  );
  al_ao21 _6169_ (
    .a(\DFF_242.Q ),
    .b(_1454_),
    .c(\DFF_243.Q ),
    .y(_1785_)
  );
  al_and3 _6170_ (
    .a(_0778_),
    .b(_1784_),
    .c(_1785_),
    .y(\DFF_243.D )
  );
  al_nand2 _6171_ (
    .a(\DFF_266.Q ),
    .b(\DFF_1428.Q ),
    .y(_1786_)
  );
  al_aoi21ttf _6172_ (
    .a(\DFF_267.Q ),
    .b(\DFF_1429.Q ),
    .c(_1786_),
    .y(_1787_)
  );
  al_ao21ftf _6173_ (
    .a(_1197_),
    .b(\DFF_265.Q ),
    .c(_1787_),
    .y(_1788_)
  );
  al_nand2ft _6174_ (
    .a(\DFF_271.Q ),
    .b(\DFF_1427.Q ),
    .y(_1789_)
  );
  al_aoi21ftf _6175_ (
    .a(\DFF_273.Q ),
    .b(\DFF_1429.Q ),
    .c(_1789_),
    .y(_1790_)
  );
  al_aoi21ftf _6176_ (
    .a(\DFF_272.Q ),
    .b(\DFF_1428.Q ),
    .c(_1790_),
    .y(_1791_)
  );
  al_nor3fft _6177_ (
    .a(_0161_),
    .b(_0165_),
    .c(_0462_),
    .y(_1792_)
  );
  al_nor2 _6178_ (
    .a(_1102_),
    .b(_0847_),
    .y(_1793_)
  );
  al_ao21ftf _6179_ (
    .a(_1793_),
    .b(_1792_),
    .c(_0170_),
    .y(_1794_)
  );
  al_aoi21ftf _6180_ (
    .a(_0170_),
    .b(_1792_),
    .c(_1794_),
    .y(_1795_)
  );
  al_ao21 _6181_ (
    .a(_1791_),
    .b(_1795_),
    .c(_1102_),
    .y(_1796_)
  );
  al_and3ftt _6182_ (
    .a(_1788_),
    .b(\DFF_1302.Q ),
    .c(_1795_),
    .y(_1797_)
  );
  al_ao21 _6183_ (
    .a(_1788_),
    .b(_1796_),
    .c(_1797_),
    .y(_1798_)
  );
  al_mux2h _6184_ (
    .a(\DFF_265.Q ),
    .b(_1798_),
    .s(\DFF_1427.Q ),
    .y(\DFF_265.D )
  );
  al_mux2h _6185_ (
    .a(\DFF_266.Q ),
    .b(_1798_),
    .s(\DFF_1428.Q ),
    .y(\DFF_266.D )
  );
  al_mux2h _6186_ (
    .a(\DFF_267.Q ),
    .b(_1798_),
    .s(\DFF_1429.Q ),
    .y(\DFF_267.D )
  );
  al_ao21 _6187_ (
    .a(\DFF_1427.Q ),
    .b(_1797_),
    .c(\DFF_271.Q ),
    .y(_1799_)
  );
  al_and2 _6188_ (
    .a(\DFF_1302.Q ),
    .b(_1788_),
    .y(_1800_)
  );
  al_and3 _6189_ (
    .a(_1791_),
    .b(_1800_),
    .c(_1795_),
    .y(_1801_)
  );
  al_aoi21ftf _6190_ (
    .a(_1197_),
    .b(_1801_),
    .c(_1799_),
    .y(\DFF_271.D )
  );
  al_ao21 _6191_ (
    .a(\DFF_1428.Q ),
    .b(_1797_),
    .c(\DFF_272.Q ),
    .y(_1802_)
  );
  al_aoi21ftf _6192_ (
    .a(_0246_),
    .b(_1801_),
    .c(_1802_),
    .y(\DFF_272.D )
  );
  al_ao21 _6193_ (
    .a(\DFF_1429.Q ),
    .b(_1797_),
    .c(\DFF_273.Q ),
    .y(_1803_)
  );
  al_aoi21ftf _6194_ (
    .a(_0344_),
    .b(_1801_),
    .c(_1803_),
    .y(\DFF_273.D )
  );
  al_inv _6195_ (
    .a(\DFF_593.Q ),
    .y(_1804_)
  );
  al_oa21ftf _6196_ (
    .a(_1804_),
    .b(_1558_),
    .c(_0449_),
    .y(_1805_)
  );
  al_aoi21ftf _6197_ (
    .a(_1804_),
    .b(_1558_),
    .c(_1805_),
    .y(\DFF_593.D )
  );
  al_nand2 _6198_ (
    .a(\DFF_616.Q ),
    .b(\DFF_1428.Q ),
    .y(_1806_)
  );
  al_aoi21ttf _6199_ (
    .a(\DFF_617.Q ),
    .b(\DFF_1429.Q ),
    .c(_1806_),
    .y(_1807_)
  );
  al_ao21ftf _6200_ (
    .a(_1197_),
    .b(\DFF_615.Q ),
    .c(_1807_),
    .y(_1808_)
  );
  al_or3fft _6201_ (
    .a(_0913_),
    .b(_0917_),
    .c(_0540_),
    .y(_1809_)
  );
  al_aoi21 _6202_ (
    .a(\DFF_1302.Q ),
    .b(_0926_),
    .c(\DFF_666.D ),
    .y(_1810_)
  );
  al_mux2l _6203_ (
    .a(\DFF_666.D ),
    .b(_1810_),
    .s(_1809_),
    .y(_1811_)
  );
  al_nand2ft _6204_ (
    .a(\DFF_621.Q ),
    .b(\DFF_1427.Q ),
    .y(_1812_)
  );
  al_aoi21ftf _6205_ (
    .a(\DFF_623.Q ),
    .b(\DFF_1429.Q ),
    .c(_1812_),
    .y(_1813_)
  );
  al_aoi21ftf _6206_ (
    .a(\DFF_622.Q ),
    .b(\DFF_1428.Q ),
    .c(_1813_),
    .y(_1814_)
  );
  al_ao21 _6207_ (
    .a(_1814_),
    .b(_1811_),
    .c(_1102_),
    .y(_1815_)
  );
  al_and3ftt _6208_ (
    .a(_1808_),
    .b(\DFF_1302.Q ),
    .c(_1811_),
    .y(_1816_)
  );
  al_ao21 _6209_ (
    .a(_1808_),
    .b(_1815_),
    .c(_1816_),
    .y(_1817_)
  );
  al_mux2h _6210_ (
    .a(\DFF_615.Q ),
    .b(_1817_),
    .s(\DFF_1427.Q ),
    .y(\DFF_615.D )
  );
  al_mux2h _6211_ (
    .a(\DFF_616.Q ),
    .b(_1817_),
    .s(\DFF_1428.Q ),
    .y(\DFF_616.D )
  );
  al_mux2h _6212_ (
    .a(\DFF_617.Q ),
    .b(_1817_),
    .s(\DFF_1429.Q ),
    .y(\DFF_617.D )
  );
  al_ao21 _6213_ (
    .a(\DFF_1427.Q ),
    .b(_1816_),
    .c(\DFF_621.Q ),
    .y(_1818_)
  );
  al_and2 _6214_ (
    .a(\DFF_1302.Q ),
    .b(_1808_),
    .y(_1819_)
  );
  al_and3 _6215_ (
    .a(_1814_),
    .b(_1819_),
    .c(_1811_),
    .y(_1820_)
  );
  al_aoi21ftf _6216_ (
    .a(_1197_),
    .b(_1820_),
    .c(_1818_),
    .y(\DFF_621.D )
  );
  al_ao21 _6217_ (
    .a(\DFF_1428.Q ),
    .b(_1816_),
    .c(\DFF_622.Q ),
    .y(_1821_)
  );
  al_aoi21ftf _6218_ (
    .a(_0246_),
    .b(_1820_),
    .c(_1821_),
    .y(\DFF_622.D )
  );
  al_ao21 _6219_ (
    .a(\DFF_1429.Q ),
    .b(_1816_),
    .c(\DFF_623.Q ),
    .y(_1822_)
  );
  al_aoi21ftf _6220_ (
    .a(_0344_),
    .b(_1820_),
    .c(_1822_),
    .y(\DFF_623.D )
  );
  al_or3fft _6221_ (
    .a(\DFF_943.Q ),
    .b(\DFF_942.Q ),
    .c(_1474_),
    .y(_1823_)
  );
  al_oai21ftf _6222_ (
    .a(\DFF_942.Q ),
    .b(_1474_),
    .c(\DFF_943.Q ),
    .y(_1824_)
  );
  al_and3 _6223_ (
    .a(_0778_),
    .b(_1823_),
    .c(_1824_),
    .y(\DFF_943.D )
  );
  al_inv _6224_ (
    .a(\DFF_1028.Q ),
    .y(_1825_)
  );
  al_mux2h _6225_ (
    .a(\DFF_1017.Q ),
    .b(\DFF_667.D ),
    .s(\DFF_1428.Q ),
    .y(_1826_)
  );
  al_mux2h _6226_ (
    .a(_1825_),
    .b(_1826_),
    .s(\DFF_1016.Q ),
    .y(\DFF_1017.D )
  );
  al_nand2 _6227_ (
    .a(\DFF_966.Q ),
    .b(\DFF_1428.Q ),
    .y(_1827_)
  );
  al_aoi21ttf _6228_ (
    .a(\DFF_967.Q ),
    .b(\DFF_1429.Q ),
    .c(_1827_),
    .y(_1828_)
  );
  al_ao21ftf _6229_ (
    .a(_1197_),
    .b(\DFF_965.Q ),
    .c(_1828_),
    .y(_1829_)
  );
  al_nand2ft _6230_ (
    .a(\DFF_971.Q ),
    .b(\DFF_1427.Q ),
    .y(_1830_)
  );
  al_aoi21ftf _6231_ (
    .a(\DFF_973.Q ),
    .b(\DFF_1429.Q ),
    .c(_1830_),
    .y(_1831_)
  );
  al_aoi21ftf _6232_ (
    .a(\DFF_972.Q ),
    .b(\DFF_1428.Q ),
    .c(_1831_),
    .y(_1832_)
  );
  al_or2 _6233_ (
    .a(_0215_),
    .b(_0217_),
    .y(_1833_)
  );
  al_and3 _6234_ (
    .a(_0953_),
    .b(_1833_),
    .c(_0618_),
    .y(_1834_)
  );
  al_or2 _6235_ (
    .a(_0222_),
    .b(_1834_),
    .y(_1835_)
  );
  al_and2 _6236_ (
    .a(_0222_),
    .b(_1834_),
    .y(_1836_)
  );
  al_or2 _6237_ (
    .a(_1102_),
    .b(_1005_),
    .y(_1837_)
  );
  al_ao21ttf _6238_ (
    .a(_1837_),
    .b(_1836_),
    .c(_1835_),
    .y(_1838_)
  );
  al_ao21 _6239_ (
    .a(_1832_),
    .b(_1838_),
    .c(_1102_),
    .y(_1839_)
  );
  al_nor2 _6240_ (
    .a(_1102_),
    .b(_1829_),
    .y(_1840_)
  );
  al_and2 _6241_ (
    .a(_1840_),
    .b(_1838_),
    .y(_1841_)
  );
  al_ao21 _6242_ (
    .a(_1829_),
    .b(_1839_),
    .c(_1841_),
    .y(_1842_)
  );
  al_mux2h _6243_ (
    .a(\DFF_965.Q ),
    .b(_1842_),
    .s(\DFF_1427.Q ),
    .y(\DFF_965.D )
  );
  al_mux2h _6244_ (
    .a(\DFF_966.Q ),
    .b(_1842_),
    .s(\DFF_1428.Q ),
    .y(\DFF_966.D )
  );
  al_mux2h _6245_ (
    .a(\DFF_967.Q ),
    .b(_1842_),
    .s(\DFF_1429.Q ),
    .y(\DFF_967.D )
  );
  al_ao21 _6246_ (
    .a(\DFF_1427.Q ),
    .b(_1841_),
    .c(\DFF_971.Q ),
    .y(_1843_)
  );
  al_and2 _6247_ (
    .a(\DFF_1302.Q ),
    .b(_1829_),
    .y(_1844_)
  );
  al_and3 _6248_ (
    .a(_1832_),
    .b(_1844_),
    .c(_1838_),
    .y(_1845_)
  );
  al_aoi21ftf _6249_ (
    .a(_1197_),
    .b(_1845_),
    .c(_1843_),
    .y(\DFF_971.D )
  );
  al_ao21 _6250_ (
    .a(\DFF_1428.Q ),
    .b(_1841_),
    .c(\DFF_972.Q ),
    .y(_1846_)
  );
  al_aoi21ftf _6251_ (
    .a(_0246_),
    .b(_1845_),
    .c(_1846_),
    .y(\DFF_972.D )
  );
  al_ao21 _6252_ (
    .a(\DFF_1429.Q ),
    .b(_1841_),
    .c(\DFF_973.Q ),
    .y(_1847_)
  );
  al_aoi21ftf _6253_ (
    .a(_0344_),
    .b(_1845_),
    .c(_1847_),
    .y(\DFF_973.D )
  );
  al_and2ft _6254_ (
    .a(\DFF_1133.Q ),
    .b(\DFF_1132.Q ),
    .y(_1848_)
  );
  al_oai21ftf _6255_ (
    .a(\DFF_1142.Q ),
    .b(\DFF_1505.Q ),
    .c(\DFF_1132.Q ),
    .y(_1849_)
  );
  al_ao21 _6256_ (
    .a(\DFF_1505.Q ),
    .b(\DFF_792.D ),
    .c(_1849_),
    .y(_1850_)
  );
  al_and2ft _6257_ (
    .a(_1848_),
    .b(_1850_),
    .y(\DFF_1142.D )
  );
  al_and2ft _6258_ (
    .a(\DFF_1099.Q ),
    .b(\DFF_1102.Q ),
    .y(_1851_)
  );
  al_oai21ftf _6259_ (
    .a(\DFF_1100.Q ),
    .b(\DFF_1504.Q ),
    .c(\DFF_1102.Q ),
    .y(_1852_)
  );
  al_ao21 _6260_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_750.D ),
    .c(_1852_),
    .y(_1853_)
  );
  al_nand2ft _6261_ (
    .a(_1851_),
    .b(_1853_),
    .y(_1854_)
  );
  al_inv _6262_ (
    .a(_1854_),
    .y(\DFF_1100.D )
  );
  al_inv _6263_ (
    .a(\DFF_1293.Q ),
    .y(_1855_)
  );
  al_oa21ftf _6264_ (
    .a(_1855_),
    .b(_1683_),
    .c(_0449_),
    .y(_1856_)
  );
  al_aoi21ftf _6265_ (
    .a(_1855_),
    .b(_1683_),
    .c(_1856_),
    .y(\DFF_1293.D )
  );
  al_nand2 _6266_ (
    .a(\DFF_1316.Q ),
    .b(\DFF_1428.Q ),
    .y(_1857_)
  );
  al_aoi21ttf _6267_ (
    .a(\DFF_1317.Q ),
    .b(\DFF_1429.Q ),
    .c(_1857_),
    .y(_1858_)
  );
  al_ao21ftf _6268_ (
    .a(_1197_),
    .b(\DFF_1315.Q ),
    .c(_1858_),
    .y(_1859_)
  );
  al_nand2ft _6269_ (
    .a(\DFF_1321.Q ),
    .b(\DFF_1427.Q ),
    .y(_1860_)
  );
  al_aoi21ftf _6270_ (
    .a(\DFF_1323.Q ),
    .b(\DFF_1429.Q ),
    .c(_1860_),
    .y(_1861_)
  );
  al_aoi21ftf _6271_ (
    .a(\DFF_1322.Q ),
    .b(\DFF_1428.Q ),
    .c(_1861_),
    .y(_1862_)
  );
  al_and3 _6272_ (
    .a(_0236_),
    .b(_0240_),
    .c(_0699_),
    .y(_1863_)
  );
  al_or2 _6273_ (
    .a(_0245_),
    .b(_1863_),
    .y(_1864_)
  );
  al_or2 _6274_ (
    .a(_1102_),
    .b(_1084_),
    .y(_1865_)
  );
  al_and2 _6275_ (
    .a(_0245_),
    .b(_1863_),
    .y(_1866_)
  );
  al_ao21ttf _6276_ (
    .a(_1865_),
    .b(_1866_),
    .c(_1864_),
    .y(_1867_)
  );
  al_ao21 _6277_ (
    .a(_1862_),
    .b(_1867_),
    .c(_1102_),
    .y(_1868_)
  );
  al_nor2 _6278_ (
    .a(_1102_),
    .b(_1859_),
    .y(_1869_)
  );
  al_and2 _6279_ (
    .a(_1869_),
    .b(_1867_),
    .y(_1870_)
  );
  al_ao21 _6280_ (
    .a(_1859_),
    .b(_1868_),
    .c(_1870_),
    .y(_1871_)
  );
  al_mux2h _6281_ (
    .a(\DFF_1315.Q ),
    .b(_1871_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1315.D )
  );
  al_mux2h _6282_ (
    .a(\DFF_1316.Q ),
    .b(_1871_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1316.D )
  );
  al_mux2h _6283_ (
    .a(\DFF_1317.Q ),
    .b(_1871_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1317.D )
  );
  al_ao21 _6284_ (
    .a(\DFF_1427.Q ),
    .b(_1870_),
    .c(\DFF_1321.Q ),
    .y(_1872_)
  );
  al_and2 _6285_ (
    .a(\DFF_1302.Q ),
    .b(_1859_),
    .y(_1873_)
  );
  al_and3 _6286_ (
    .a(_1862_),
    .b(_1873_),
    .c(_1867_),
    .y(_1874_)
  );
  al_aoi21ftf _6287_ (
    .a(_1197_),
    .b(_1874_),
    .c(_1872_),
    .y(\DFF_1321.D )
  );
  al_ao21 _6288_ (
    .a(\DFF_1428.Q ),
    .b(_1870_),
    .c(\DFF_1322.Q ),
    .y(_1875_)
  );
  al_aoi21ftf _6289_ (
    .a(_0246_),
    .b(_1874_),
    .c(_1875_),
    .y(\DFF_1322.D )
  );
  al_ao21 _6290_ (
    .a(\DFF_1429.Q ),
    .b(_1870_),
    .c(\DFF_1323.Q ),
    .y(_1876_)
  );
  al_aoi21ftf _6291_ (
    .a(_0344_),
    .b(_1874_),
    .c(_1876_),
    .y(\DFF_1323.D )
  );
  al_inv _6292_ (
    .a(\DFF_244.Q ),
    .y(_1877_)
  );
  al_nand3fft _6293_ (
    .a(_1782_),
    .b(_1877_),
    .c(_1496_),
    .y(_1878_)
  );
  al_nand2 _6294_ (
    .a(_1877_),
    .b(_1784_),
    .y(_1879_)
  );
  al_and3 _6295_ (
    .a(_0778_),
    .b(_1879_),
    .c(_1878_),
    .y(\DFF_244.D )
  );
  al_nand2 _6296_ (
    .a(\DFF_222.Q ),
    .b(\DFF_1428.Q ),
    .y(_1880_)
  );
  al_aoi21ttf _6297_ (
    .a(\DFF_223.Q ),
    .b(\DFF_1429.Q ),
    .c(_1880_),
    .y(_1881_)
  );
  al_aoi21ftf _6298_ (
    .a(_1197_),
    .b(\DFF_221.Q ),
    .c(_1881_),
    .y(_1882_)
  );
  al_nor2 _6299_ (
    .a(\DFF_70.Q ),
    .b(_1882_),
    .y(_1883_)
  );
  al_and2 _6300_ (
    .a(\DFF_70.Q ),
    .b(_1882_),
    .y(_1884_)
  );
  al_nand2 _6301_ (
    .a(\DFF_227.Q ),
    .b(\DFF_1427.Q ),
    .y(_1885_)
  );
  al_nand2 _6302_ (
    .a(\DFF_228.Q ),
    .b(\DFF_1428.Q ),
    .y(_1886_)
  );
  al_aoi21ttf _6303_ (
    .a(\DFF_229.Q ),
    .b(\DFF_1429.Q ),
    .c(_1886_),
    .y(_1887_)
  );
  al_ao21 _6304_ (
    .a(_1885_),
    .b(_1887_),
    .c(\DFF_298.D ),
    .y(_1888_)
  );
  al_and3 _6305_ (
    .a(\DFF_298.D ),
    .b(_1885_),
    .c(_1887_),
    .y(_1889_)
  );
  al_nand2ft _6306_ (
    .a(_1889_),
    .b(_1888_),
    .y(_1890_)
  );
  al_nand3fft _6307_ (
    .a(_1884_),
    .b(_1883_),
    .c(_1890_),
    .y(_1891_)
  );
  al_nand2 _6308_ (
    .a(\DFF_206.Q ),
    .b(\DFF_1427.Q ),
    .y(_1892_)
  );
  al_nand2 _6309_ (
    .a(\DFF_207.Q ),
    .b(\DFF_1428.Q ),
    .y(_1893_)
  );
  al_aoi21ttf _6310_ (
    .a(\DFF_208.Q ),
    .b(\DFF_1429.Q ),
    .c(_1893_),
    .y(_1894_)
  );
  al_ao21 _6311_ (
    .a(_1892_),
    .b(_1894_),
    .c(\DFF_312.D ),
    .y(_1895_)
  );
  al_and3 _6312_ (
    .a(\DFF_312.D ),
    .b(_1892_),
    .c(_1894_),
    .y(_1896_)
  );
  al_nand2ft _6313_ (
    .a(_1896_),
    .b(_1895_),
    .y(_1897_)
  );
  al_nand2 _6314_ (
    .a(\DFF_225.Q ),
    .b(\DFF_1428.Q ),
    .y(_1898_)
  );
  al_aoi21ttf _6315_ (
    .a(\DFF_226.Q ),
    .b(\DFF_1429.Q ),
    .c(_1898_),
    .y(_1899_)
  );
  al_ao21ftf _6316_ (
    .a(_1197_),
    .b(\DFF_224.Q ),
    .c(_1899_),
    .y(_1900_)
  );
  al_and2 _6317_ (
    .a(\DFF_68.Q ),
    .b(_1900_),
    .y(_1901_)
  );
  al_or2 _6318_ (
    .a(\DFF_68.Q ),
    .b(_1900_),
    .y(_1902_)
  );
  al_nand2ft _6319_ (
    .a(_1901_),
    .b(_1902_),
    .y(_1903_)
  );
  al_nand2 _6320_ (
    .a(\DFF_212.Q ),
    .b(\DFF_1427.Q ),
    .y(_1904_)
  );
  al_nand2 _6321_ (
    .a(\DFF_213.Q ),
    .b(\DFF_1428.Q ),
    .y(_1905_)
  );
  al_aoi21ttf _6322_ (
    .a(\DFF_214.Q ),
    .b(\DFF_1429.Q ),
    .c(_1905_),
    .y(_1906_)
  );
  al_ao21 _6323_ (
    .a(_1904_),
    .b(_1906_),
    .c(\DFF_308.D ),
    .y(_1907_)
  );
  al_and3 _6324_ (
    .a(\DFF_308.D ),
    .b(_1904_),
    .c(_1906_),
    .y(_1908_)
  );
  al_nand2ft _6325_ (
    .a(_1908_),
    .b(_1907_),
    .y(_1909_)
  );
  al_nand2 _6326_ (
    .a(\DFF_231.Q ),
    .b(\DFF_1428.Q ),
    .y(_1910_)
  );
  al_aoi21ttf _6327_ (
    .a(\DFF_232.Q ),
    .b(\DFF_1429.Q ),
    .c(_1910_),
    .y(_1911_)
  );
  al_ao21ftf _6328_ (
    .a(_1197_),
    .b(\DFF_230.Q ),
    .c(_1911_),
    .y(_1912_)
  );
  al_nand2ft _6329_ (
    .a(_0161_),
    .b(_1912_),
    .y(_1913_)
  );
  al_nand2ft _6330_ (
    .a(_1912_),
    .b(_0161_),
    .y(_1914_)
  );
  al_and3 _6331_ (
    .a(_1913_),
    .b(_1914_),
    .c(_1909_),
    .y(_1915_)
  );
  al_and3 _6332_ (
    .a(_1897_),
    .b(_1903_),
    .c(_1915_),
    .y(_1916_)
  );
  al_nand2 _6333_ (
    .a(\DFF_215.Q ),
    .b(\DFF_1427.Q ),
    .y(_1917_)
  );
  al_nand2 _6334_ (
    .a(\DFF_216.Q ),
    .b(\DFF_1428.Q ),
    .y(_1918_)
  );
  al_aoi21ttf _6335_ (
    .a(\DFF_217.Q ),
    .b(\DFF_1429.Q ),
    .c(_1918_),
    .y(_1919_)
  );
  al_ao21 _6336_ (
    .a(_1917_),
    .b(_1919_),
    .c(\DFF_306.D ),
    .y(_1920_)
  );
  al_and3 _6337_ (
    .a(\DFF_306.D ),
    .b(_1917_),
    .c(_1919_),
    .y(_1921_)
  );
  al_nand2ft _6338_ (
    .a(_1921_),
    .b(_1920_),
    .y(_1922_)
  );
  al_nand2 _6339_ (
    .a(\DFF_233.Q ),
    .b(\DFF_1427.Q ),
    .y(_1923_)
  );
  al_nand2 _6340_ (
    .a(\DFF_234.Q ),
    .b(\DFF_1428.Q ),
    .y(_1924_)
  );
  al_aoi21ttf _6341_ (
    .a(\DFF_235.Q ),
    .b(\DFF_1429.Q ),
    .c(_1924_),
    .y(_1925_)
  );
  al_ao21 _6342_ (
    .a(_1923_),
    .b(_1925_),
    .c(_0165_),
    .y(_1926_)
  );
  al_nand3 _6343_ (
    .a(_1923_),
    .b(_1925_),
    .c(_0165_),
    .y(_1927_)
  );
  al_and2 _6344_ (
    .a(_1927_),
    .b(_1926_),
    .y(_1928_)
  );
  al_nand2 _6345_ (
    .a(\DFF_219.Q ),
    .b(\DFF_1428.Q ),
    .y(_1929_)
  );
  al_aoi21ttf _6346_ (
    .a(\DFF_220.Q ),
    .b(\DFF_1429.Q ),
    .c(_1929_),
    .y(_1930_)
  );
  al_ao21ftf _6347_ (
    .a(_1197_),
    .b(\DFF_218.Q ),
    .c(_1930_),
    .y(_1931_)
  );
  al_and2 _6348_ (
    .a(\DFF_304.D ),
    .b(_1931_),
    .y(_1932_)
  );
  al_or2 _6349_ (
    .a(\DFF_304.D ),
    .b(_1931_),
    .y(_1933_)
  );
  al_nand2 _6350_ (
    .a(\DFF_209.Q ),
    .b(\DFF_1427.Q ),
    .y(_1934_)
  );
  al_nand2 _6351_ (
    .a(\DFF_210.Q ),
    .b(\DFF_1428.Q ),
    .y(_1935_)
  );
  al_aoi21ttf _6352_ (
    .a(\DFF_211.Q ),
    .b(\DFF_1429.Q ),
    .c(_1935_),
    .y(_1936_)
  );
  al_ao21 _6353_ (
    .a(_1934_),
    .b(_1936_),
    .c(\DFF_310.D ),
    .y(_1937_)
  );
  al_and3 _6354_ (
    .a(\DFF_310.D ),
    .b(_1934_),
    .c(_1936_),
    .y(_1938_)
  );
  al_and2ft _6355_ (
    .a(_1938_),
    .b(_1937_),
    .y(_1939_)
  );
  al_or3ftt _6356_ (
    .a(_1933_),
    .b(_1932_),
    .c(_1939_),
    .y(_1940_)
  );
  al_nor3fft _6357_ (
    .a(_1922_),
    .b(_1928_),
    .c(_1940_),
    .y(_1941_)
  );
  al_nand3ftt _6358_ (
    .a(_1891_),
    .b(_1941_),
    .c(_1916_),
    .y(_1942_)
  );
  al_ao21 _6359_ (
    .a(_0847_),
    .b(_1942_),
    .c(_0276_),
    .y(_1943_)
  );
  al_and2 _6360_ (
    .a(_0156_),
    .b(_1943_),
    .y(_1944_)
  );
  al_inv _6361_ (
    .a(_0273_),
    .y(_1945_)
  );
  al_or2 _6362_ (
    .a(_1884_),
    .b(_1883_),
    .y(_1946_)
  );
  al_ao21ftf _6363_ (
    .a(_1939_),
    .b(_1890_),
    .c(_1946_),
    .y(_1947_)
  );
  al_ao21ftf _6364_ (
    .a(_1938_),
    .b(_1937_),
    .c(_1922_),
    .y(_1948_)
  );
  al_ao21ttf _6365_ (
    .a(_1926_),
    .b(_1927_),
    .c(_1948_),
    .y(_1949_)
  );
  al_aoi21ttf _6366_ (
    .a(_1922_),
    .b(_1928_),
    .c(_1891_),
    .y(_1950_)
  );
  al_ao21ttf _6367_ (
    .a(_1949_),
    .b(_1947_),
    .c(_1950_),
    .y(_1951_)
  );
  al_nand3fft _6368_ (
    .a(_1884_),
    .b(_1883_),
    .c(_1922_),
    .y(_1952_)
  );
  al_nand3 _6369_ (
    .a(_1927_),
    .b(_1926_),
    .c(_1890_),
    .y(_1953_)
  );
  al_and3 _6370_ (
    .a(_1939_),
    .b(_1953_),
    .c(_1952_),
    .y(_1954_)
  );
  al_and2ft _6371_ (
    .a(_1954_),
    .b(_1951_),
    .y(_1955_)
  );
  al_nand2ft _6372_ (
    .a(_1932_),
    .b(_1933_),
    .y(_1956_)
  );
  al_ao21ttf _6373_ (
    .a(_1897_),
    .b(_1903_),
    .c(_1956_),
    .y(_1957_)
  );
  al_ao21ftf _6374_ (
    .a(_1908_),
    .b(_1907_),
    .c(_1897_),
    .y(_1958_)
  );
  al_aoi21ttf _6375_ (
    .a(_1913_),
    .b(_1914_),
    .c(_1958_),
    .y(_1959_)
  );
  al_aoi21ftt _6376_ (
    .a(_1956_),
    .b(_1903_),
    .c(_1915_),
    .y(_1960_)
  );
  al_ao21ftf _6377_ (
    .a(_1959_),
    .b(_1957_),
    .c(_1960_),
    .y(_1961_)
  );
  al_nand3 _6378_ (
    .a(_1913_),
    .b(_1914_),
    .c(_1903_),
    .y(_1962_)
  );
  al_nand3ftt _6379_ (
    .a(_1932_),
    .b(_1933_),
    .c(_1909_),
    .y(_1963_)
  );
  al_nand3ftt _6380_ (
    .a(_1897_),
    .b(_1963_),
    .c(_1962_),
    .y(_1964_)
  );
  al_ao21 _6381_ (
    .a(_1964_),
    .b(_1961_),
    .c(_0848_),
    .y(_1965_)
  );
  al_oa21 _6382_ (
    .a(_0848_),
    .b(_1955_),
    .c(_1965_),
    .y(_1966_)
  );
  al_mux2h _6383_ (
    .a(_1945_),
    .b(_1966_),
    .s(_0270_),
    .y(_1967_)
  );
  al_nand3 _6384_ (
    .a(_0267_),
    .b(_0851_),
    .c(_1967_),
    .y(_1968_)
  );
  al_mux2h _6385_ (
    .a(\DFF_292.Q ),
    .b(_1968_),
    .s(_1944_),
    .y(\DFF_292.D )
  );
  al_and2 _6386_ (
    .a(_0157_),
    .b(_1943_),
    .y(_1969_)
  );
  al_mux2h _6387_ (
    .a(\DFF_293.Q ),
    .b(_1968_),
    .s(_1969_),
    .y(\DFF_293.D )
  );
  al_and2 _6388_ (
    .a(_0158_),
    .b(_1943_),
    .y(_1970_)
  );
  al_mux2h _6389_ (
    .a(\DFF_294.Q ),
    .b(_1968_),
    .s(_1970_),
    .y(\DFF_294.D )
  );
  al_or3fft _6390_ (
    .a(\DFF_1302.Q ),
    .b(_1788_),
    .c(_1791_),
    .y(_1971_)
  );
  al_ao21ftf _6391_ (
    .a(_1793_),
    .b(_1971_),
    .c(_1792_),
    .y(_1972_)
  );
  al_ao21ftf _6392_ (
    .a(_0170_),
    .b(_1971_),
    .c(_1972_),
    .y(_1973_)
  );
  al_mux2h _6393_ (
    .a(\DFF_268.Q ),
    .b(_1973_),
    .s(\DFF_1427.Q ),
    .y(\DFF_268.D )
  );
  al_mux2h _6394_ (
    .a(\DFF_269.Q ),
    .b(_1973_),
    .s(\DFF_1428.Q ),
    .y(\DFF_269.D )
  );
  al_mux2h _6395_ (
    .a(\DFF_270.Q ),
    .b(_1973_),
    .s(\DFF_1429.Q ),
    .y(\DFF_270.D )
  );
  al_nand3 _6396_ (
    .a(\DFF_593.Q ),
    .b(\DFF_594.Q ),
    .c(_1558_),
    .y(_1974_)
  );
  al_ao21 _6397_ (
    .a(\DFF_593.Q ),
    .b(_1558_),
    .c(\DFF_594.Q ),
    .y(_1975_)
  );
  al_and3 _6398_ (
    .a(_0778_),
    .b(_1974_),
    .c(_1975_),
    .y(\DFF_594.D )
  );
  al_nand2 _6399_ (
    .a(\DFF_556.Q ),
    .b(\DFF_1427.Q ),
    .y(_1976_)
  );
  al_nand2 _6400_ (
    .a(\DFF_557.Q ),
    .b(\DFF_1428.Q ),
    .y(_1977_)
  );
  al_aoi21ttf _6401_ (
    .a(\DFF_558.Q ),
    .b(\DFF_1429.Q ),
    .c(_1977_),
    .y(_1978_)
  );
  al_aoi21 _6402_ (
    .a(_1976_),
    .b(_1978_),
    .c(\DFF_62.Q ),
    .y(_1979_)
  );
  al_and3 _6403_ (
    .a(\DFF_62.Q ),
    .b(_1976_),
    .c(_1978_),
    .y(_1980_)
  );
  al_nor2 _6404_ (
    .a(_1980_),
    .b(_1979_),
    .y(_1981_)
  );
  al_nand2 _6405_ (
    .a(\DFF_562.Q ),
    .b(\DFF_1427.Q ),
    .y(_1982_)
  );
  al_nand2 _6406_ (
    .a(\DFF_563.Q ),
    .b(\DFF_1428.Q ),
    .y(_1983_)
  );
  al_aoi21ttf _6407_ (
    .a(\DFF_564.Q ),
    .b(\DFF_1429.Q ),
    .c(_1983_),
    .y(_1984_)
  );
  al_aoi21 _6408_ (
    .a(_1982_),
    .b(_1984_),
    .c(\DFF_58.Q ),
    .y(_1985_)
  );
  al_nand3 _6409_ (
    .a(\DFF_58.Q ),
    .b(_1982_),
    .c(_1984_),
    .y(_1986_)
  );
  al_nand3ftt _6410_ (
    .a(_1985_),
    .b(_1986_),
    .c(_1981_),
    .y(_1987_)
  );
  al_nand2 _6411_ (
    .a(\DFF_571.Q ),
    .b(\DFF_1427.Q ),
    .y(_1988_)
  );
  al_nand2 _6412_ (
    .a(\DFF_572.Q ),
    .b(\DFF_1428.Q ),
    .y(_1989_)
  );
  al_aoi21ttf _6413_ (
    .a(\DFF_573.Q ),
    .b(\DFF_1429.Q ),
    .c(_1989_),
    .y(_1990_)
  );
  al_ao21 _6414_ (
    .a(_1988_),
    .b(_1990_),
    .c(\DFF_652.D ),
    .y(_1991_)
  );
  al_and3 _6415_ (
    .a(\DFF_652.D ),
    .b(_1988_),
    .c(_1990_),
    .y(_1992_)
  );
  al_nand2ft _6416_ (
    .a(_1992_),
    .b(_1991_),
    .y(_1993_)
  );
  al_nand2 _6417_ (
    .a(\DFF_577.Q ),
    .b(\DFF_1427.Q ),
    .y(_1994_)
  );
  al_nand2 _6418_ (
    .a(\DFF_578.Q ),
    .b(\DFF_1428.Q ),
    .y(_1995_)
  );
  al_aoi21ttf _6419_ (
    .a(\DFF_579.Q ),
    .b(\DFF_1429.Q ),
    .c(_1995_),
    .y(_1996_)
  );
  al_ao21 _6420_ (
    .a(_1994_),
    .b(_1996_),
    .c(\DFF_48.Q ),
    .y(_1997_)
  );
  al_nand3 _6421_ (
    .a(\DFF_48.Q ),
    .b(_1994_),
    .c(_1996_),
    .y(_1998_)
  );
  al_nand3 _6422_ (
    .a(_1997_),
    .b(_1998_),
    .c(_1993_),
    .y(_1999_)
  );
  al_nand2 _6423_ (
    .a(\DFF_565.Q ),
    .b(\DFF_1427.Q ),
    .y(_2000_)
  );
  al_nand2 _6424_ (
    .a(\DFF_566.Q ),
    .b(\DFF_1428.Q ),
    .y(_2001_)
  );
  al_aoi21ttf _6425_ (
    .a(\DFF_567.Q ),
    .b(\DFF_1429.Q ),
    .c(_2001_),
    .y(_2002_)
  );
  al_ao21 _6426_ (
    .a(_2000_),
    .b(_2002_),
    .c(\DFF_656.D ),
    .y(_2003_)
  );
  al_and3 _6427_ (
    .a(\DFF_656.D ),
    .b(_2000_),
    .c(_2002_),
    .y(_2004_)
  );
  al_nand2ft _6428_ (
    .a(_2004_),
    .b(_2003_),
    .y(_2005_)
  );
  al_nand2 _6429_ (
    .a(\DFF_559.Q ),
    .b(\DFF_1427.Q ),
    .y(_2006_)
  );
  al_nand2 _6430_ (
    .a(\DFF_560.Q ),
    .b(\DFF_1428.Q ),
    .y(_2007_)
  );
  al_aoi21ttf _6431_ (
    .a(\DFF_561.Q ),
    .b(\DFF_1429.Q ),
    .c(_2007_),
    .y(_2008_)
  );
  al_ao21 _6432_ (
    .a(_2006_),
    .b(_2008_),
    .c(\DFF_660.D ),
    .y(_2009_)
  );
  al_and3 _6433_ (
    .a(\DFF_660.D ),
    .b(_2006_),
    .c(_2008_),
    .y(_2010_)
  );
  al_aoi21ftf _6434_ (
    .a(_2010_),
    .b(_2009_),
    .c(_2005_),
    .y(_2011_)
  );
  al_and3fft _6435_ (
    .a(_1999_),
    .b(_1987_),
    .c(_2011_),
    .y(_2012_)
  );
  al_nand2 _6436_ (
    .a(\DFF_583.Q ),
    .b(\DFF_1427.Q ),
    .y(_2013_)
  );
  al_nand2 _6437_ (
    .a(\DFF_584.Q ),
    .b(\DFF_1428.Q ),
    .y(_2014_)
  );
  al_aoi21ttf _6438_ (
    .a(\DFF_585.Q ),
    .b(\DFF_1429.Q ),
    .c(_2014_),
    .y(_2015_)
  );
  al_ao21ttf _6439_ (
    .a(_2013_),
    .b(_2015_),
    .c(_0195_),
    .y(_2016_)
  );
  al_and3 _6440_ (
    .a(_2013_),
    .b(_2015_),
    .c(_0917_),
    .y(_2017_)
  );
  al_nand2ft _6441_ (
    .a(_2017_),
    .b(_2016_),
    .y(_2018_)
  );
  al_nand2 _6442_ (
    .a(\DFF_580.Q ),
    .b(\DFF_1427.Q ),
    .y(_2019_)
  );
  al_nand2 _6443_ (
    .a(\DFF_581.Q ),
    .b(\DFF_1428.Q ),
    .y(_2020_)
  );
  al_aoi21ttf _6444_ (
    .a(\DFF_582.Q ),
    .b(\DFF_1429.Q ),
    .c(_2020_),
    .y(_2021_)
  );
  al_ao21ttf _6445_ (
    .a(_2019_),
    .b(_2021_),
    .c(_0191_),
    .y(_2022_)
  );
  al_nand3 _6446_ (
    .a(_2019_),
    .b(_2021_),
    .c(_0913_),
    .y(_2023_)
  );
  al_nand2 _6447_ (
    .a(_2023_),
    .b(_2022_),
    .y(_2024_)
  );
  al_nand2 _6448_ (
    .a(\DFF_568.Q ),
    .b(\DFF_1427.Q ),
    .y(_2025_)
  );
  al_nand2 _6449_ (
    .a(\DFF_569.Q ),
    .b(\DFF_1428.Q ),
    .y(_2026_)
  );
  al_aoi21ttf _6450_ (
    .a(\DFF_570.Q ),
    .b(\DFF_1429.Q ),
    .c(_2026_),
    .y(_2027_)
  );
  al_ao21 _6451_ (
    .a(_2025_),
    .b(_2027_),
    .c(\DFF_654.D ),
    .y(_2028_)
  );
  al_and3 _6452_ (
    .a(\DFF_654.D ),
    .b(_2025_),
    .c(_2027_),
    .y(_2029_)
  );
  al_nand2ft _6453_ (
    .a(_2029_),
    .b(_2028_),
    .y(_2030_)
  );
  al_nand2 _6454_ (
    .a(\DFF_574.Q ),
    .b(\DFF_1427.Q ),
    .y(_2031_)
  );
  al_nand2 _6455_ (
    .a(\DFF_575.Q ),
    .b(\DFF_1428.Q ),
    .y(_2032_)
  );
  al_aoi21ttf _6456_ (
    .a(\DFF_576.Q ),
    .b(\DFF_1429.Q ),
    .c(_2032_),
    .y(_2033_)
  );
  al_ao21 _6457_ (
    .a(_2031_),
    .b(_2033_),
    .c(\DFF_650.D ),
    .y(_2034_)
  );
  al_and3 _6458_ (
    .a(\DFF_650.D ),
    .b(_2031_),
    .c(_2033_),
    .y(_2035_)
  );
  al_aoi21ftf _6459_ (
    .a(_2035_),
    .b(_2034_),
    .c(_2030_),
    .y(_2036_)
  );
  al_and3fft _6460_ (
    .a(_2018_),
    .b(_2024_),
    .c(_2036_),
    .y(_2037_)
  );
  al_ao21 _6461_ (
    .a(_2037_),
    .b(_2012_),
    .c(_0926_),
    .y(_2038_)
  );
  al_aoi21ftf _6462_ (
    .a(_0292_),
    .b(_2038_),
    .c(_0156_),
    .y(_2039_)
  );
  al_nand3ftt _6463_ (
    .a(_2017_),
    .b(_2016_),
    .c(_2005_),
    .y(_2040_)
  );
  al_nand2ft _6464_ (
    .a(_2010_),
    .b(_2009_),
    .y(_2041_)
  );
  al_and2 _6465_ (
    .a(_1998_),
    .b(_1997_),
    .y(_2042_)
  );
  al_aoi21 _6466_ (
    .a(_2041_),
    .b(_2042_),
    .c(_1993_),
    .y(_2043_)
  );
  al_aoi21ttf _6467_ (
    .a(_2005_),
    .b(_2041_),
    .c(_2018_),
    .y(_2044_)
  );
  al_ao21 _6468_ (
    .a(_1999_),
    .b(_2044_),
    .c(_2043_),
    .y(_2045_)
  );
  al_aoi21 _6469_ (
    .a(_1993_),
    .b(_2005_),
    .c(_2041_),
    .y(_2046_)
  );
  al_aoi21ftf _6470_ (
    .a(_2018_),
    .b(_2042_),
    .c(_2046_),
    .y(_2047_)
  );
  al_aoi21 _6471_ (
    .a(_2040_),
    .b(_2045_),
    .c(_2047_),
    .y(_2048_)
  );
  al_or3 _6472_ (
    .a(_1102_),
    .b(_0926_),
    .c(_2048_),
    .y(_2049_)
  );
  al_or2 _6473_ (
    .a(_1102_),
    .b(_0926_),
    .y(_2050_)
  );
  al_nand2ft _6474_ (
    .a(_2035_),
    .b(_2034_),
    .y(_2051_)
  );
  al_nor2ft _6475_ (
    .a(_1986_),
    .b(_1985_),
    .y(_2052_)
  );
  al_aoi21 _6476_ (
    .a(_2030_),
    .b(_2052_),
    .c(_1981_),
    .y(_2053_)
  );
  al_ao21ftf _6477_ (
    .a(_2024_),
    .b(_2051_),
    .c(_2053_),
    .y(_2054_)
  );
  al_and2ft _6478_ (
    .a(_2029_),
    .b(_2028_),
    .y(_2055_)
  );
  al_nand3 _6479_ (
    .a(_2022_),
    .b(_2023_),
    .c(_2052_),
    .y(_2056_)
  );
  al_nand3fft _6480_ (
    .a(_1979_),
    .b(_1980_),
    .c(_2051_),
    .y(_2057_)
  );
  al_nand3 _6481_ (
    .a(_2055_),
    .b(_2057_),
    .c(_2056_),
    .y(_2058_)
  );
  al_aoi21ttf _6482_ (
    .a(_1981_),
    .b(_2052_),
    .c(_2024_),
    .y(_2059_)
  );
  al_aoi21ftf _6483_ (
    .a(_2036_),
    .b(_2059_),
    .c(_2058_),
    .y(_2060_)
  );
  al_ao21 _6484_ (
    .a(_2054_),
    .b(_2060_),
    .c(_2050_),
    .y(_2061_)
  );
  al_and3 _6485_ (
    .a(_0284_),
    .b(_2061_),
    .c(_2049_),
    .y(_2062_)
  );
  al_and2ft _6486_ (
    .a(_0923_),
    .b(_0921_),
    .y(_2063_)
  );
  al_and3 _6487_ (
    .a(_0893_),
    .b(_0892_),
    .c(_2063_),
    .y(_2064_)
  );
  al_oa21ttf _6488_ (
    .a(_0874_),
    .b(_0873_),
    .c(_2050_),
    .y(_2065_)
  );
  al_nand3 _6489_ (
    .a(_0888_),
    .b(_2064_),
    .c(_2065_),
    .y(_2066_)
  );
  al_nand2ft _6490_ (
    .a(_0917_),
    .b(_0902_),
    .y(_2067_)
  );
  al_and2 _6491_ (
    .a(_0914_),
    .b(_0912_),
    .y(_2068_)
  );
  al_nand3 _6492_ (
    .a(_2067_),
    .b(_2068_),
    .c(_0869_),
    .y(_2069_)
  );
  al_or2ft _6493_ (
    .a(_0899_),
    .b(_0898_),
    .y(_2070_)
  );
  al_ao21ftt _6494_ (
    .a(_0902_),
    .b(_0917_),
    .c(_0881_),
    .y(_2071_)
  );
  al_nor2 _6495_ (
    .a(_0915_),
    .b(_0906_),
    .y(_2072_)
  );
  al_nor3fft _6496_ (
    .a(_2072_),
    .b(_2070_),
    .c(_2071_),
    .y(_2073_)
  );
  al_and3fft _6497_ (
    .a(_2069_),
    .b(_2066_),
    .c(_2073_),
    .y(_2074_)
  );
  al_nand2ft _6498_ (
    .a(_0281_),
    .b(_2074_),
    .y(_2075_)
  );
  al_oai21ftf _6499_ (
    .a(_0291_),
    .b(_2062_),
    .c(_2075_),
    .y(_2076_)
  );
  al_mux2h _6500_ (
    .a(\DFF_642.Q ),
    .b(_2076_),
    .s(_2039_),
    .y(\DFF_642.D )
  );
  al_aoi21ftf _6501_ (
    .a(_0292_),
    .b(_2038_),
    .c(_0157_),
    .y(_2077_)
  );
  al_mux2h _6502_ (
    .a(\DFF_643.Q ),
    .b(_2076_),
    .s(_2077_),
    .y(\DFF_643.D )
  );
  al_aoi21ftf _6503_ (
    .a(_0292_),
    .b(_2038_),
    .c(_0158_),
    .y(_2078_)
  );
  al_mux2h _6504_ (
    .a(\DFF_644.Q ),
    .b(_2076_),
    .s(_2078_),
    .y(\DFF_644.D )
  );
  al_or3fft _6505_ (
    .a(\DFF_1302.Q ),
    .b(_1808_),
    .c(_1814_),
    .y(_2079_)
  );
  al_ao21ttf _6506_ (
    .a(\DFF_666.D ),
    .b(_2079_),
    .c(_1809_),
    .y(_2080_)
  );
  al_aoi21ttf _6507_ (
    .a(_1810_),
    .b(_2079_),
    .c(_2080_),
    .y(_2081_)
  );
  al_mux2h _6508_ (
    .a(\DFF_618.Q ),
    .b(_2081_),
    .s(\DFF_1427.Q ),
    .y(\DFF_618.D )
  );
  al_mux2h _6509_ (
    .a(\DFF_619.Q ),
    .b(_2081_),
    .s(\DFF_1428.Q ),
    .y(\DFF_619.D )
  );
  al_mux2h _6510_ (
    .a(\DFF_620.Q ),
    .b(_2081_),
    .s(\DFF_1429.Q ),
    .y(\DFF_620.D )
  );
  al_nand3 _6511_ (
    .a(\DFF_943.Q ),
    .b(\DFF_944.Q ),
    .c(_1621_),
    .y(_2082_)
  );
  al_ao21 _6512_ (
    .a(\DFF_943.Q ),
    .b(_1621_),
    .c(\DFF_944.Q ),
    .y(_2083_)
  );
  al_and3 _6513_ (
    .a(_0778_),
    .b(_2082_),
    .c(_2083_),
    .y(\DFF_944.D )
  );
  al_inv _6514_ (
    .a(_1005_),
    .y(_2084_)
  );
  al_nand2 _6515_ (
    .a(\DFF_918.Q ),
    .b(\DFF_1427.Q ),
    .y(_2085_)
  );
  al_nand2 _6516_ (
    .a(\DFF_919.Q ),
    .b(\DFF_1428.Q ),
    .y(_2086_)
  );
  al_aoi21ttf _6517_ (
    .a(\DFF_920.Q ),
    .b(\DFF_1429.Q ),
    .c(_2086_),
    .y(_2087_)
  );
  al_ao21 _6518_ (
    .a(_2085_),
    .b(_2087_),
    .c(\DFF_41.Q ),
    .y(_2088_)
  );
  al_and3 _6519_ (
    .a(\DFF_41.Q ),
    .b(_2085_),
    .c(_2087_),
    .y(_2089_)
  );
  al_nand2 _6520_ (
    .a(\DFF_924.Q ),
    .b(\DFF_1427.Q ),
    .y(_2090_)
  );
  al_nand2 _6521_ (
    .a(\DFF_925.Q ),
    .b(\DFF_1428.Q ),
    .y(_2091_)
  );
  al_aoi21ttf _6522_ (
    .a(\DFF_926.Q ),
    .b(\DFF_1429.Q ),
    .c(_2091_),
    .y(_2092_)
  );
  al_ao21 _6523_ (
    .a(_2090_),
    .b(_2092_),
    .c(\DFF_1000.D ),
    .y(_2093_)
  );
  al_and3 _6524_ (
    .a(\DFF_1000.D ),
    .b(_2090_),
    .c(_2092_),
    .y(_2094_)
  );
  al_nand2ft _6525_ (
    .a(_2094_),
    .b(_2093_),
    .y(_2095_)
  );
  al_and3ftt _6526_ (
    .a(_2089_),
    .b(_2088_),
    .c(_2095_),
    .y(_2096_)
  );
  al_nand2 _6527_ (
    .a(\DFF_909.Q ),
    .b(\DFF_1427.Q ),
    .y(_2097_)
  );
  al_nand2 _6528_ (
    .a(\DFF_910.Q ),
    .b(\DFF_1428.Q ),
    .y(_2098_)
  );
  al_aoi21ttf _6529_ (
    .a(\DFF_911.Q ),
    .b(\DFF_1429.Q ),
    .c(_2098_),
    .y(_2099_)
  );
  al_ao21 _6530_ (
    .a(_2097_),
    .b(_2099_),
    .c(\DFF_1010.D ),
    .y(_2100_)
  );
  al_and3 _6531_ (
    .a(\DFF_1010.D ),
    .b(_2097_),
    .c(_2099_),
    .y(_2101_)
  );
  al_nand2ft _6532_ (
    .a(_2101_),
    .b(_2100_),
    .y(_2102_)
  );
  al_nand2 _6533_ (
    .a(\DFF_906.Q ),
    .b(\DFF_1427.Q ),
    .y(_2103_)
  );
  al_nand2 _6534_ (
    .a(\DFF_907.Q ),
    .b(\DFF_1428.Q ),
    .y(_2104_)
  );
  al_aoi21ttf _6535_ (
    .a(\DFF_908.Q ),
    .b(\DFF_1429.Q ),
    .c(_2104_),
    .y(_2105_)
  );
  al_aoi21 _6536_ (
    .a(_2103_),
    .b(_2105_),
    .c(\DFF_45.Q ),
    .y(_2106_)
  );
  al_and3 _6537_ (
    .a(\DFF_45.Q ),
    .b(_2103_),
    .c(_2105_),
    .y(_2107_)
  );
  al_nor2 _6538_ (
    .a(_2107_),
    .b(_2106_),
    .y(_2108_)
  );
  al_and3 _6539_ (
    .a(_2102_),
    .b(_2108_),
    .c(_2096_),
    .y(_2109_)
  );
  al_nand2 _6540_ (
    .a(\DFF_930.Q ),
    .b(\DFF_1427.Q ),
    .y(_2110_)
  );
  al_nand2 _6541_ (
    .a(\DFF_931.Q ),
    .b(\DFF_1428.Q ),
    .y(_2111_)
  );
  al_aoi21ttf _6542_ (
    .a(\DFF_932.Q ),
    .b(\DFF_1429.Q ),
    .c(_2111_),
    .y(_2112_)
  );
  al_ao21ttf _6543_ (
    .a(_2110_),
    .b(_2112_),
    .c(_0214_),
    .y(_2113_)
  );
  al_and3 _6544_ (
    .a(_2110_),
    .b(_2112_),
    .c(_0953_),
    .y(_2114_)
  );
  al_nand2 _6545_ (
    .a(\DFF_912.Q ),
    .b(\DFF_1427.Q ),
    .y(_2115_)
  );
  al_nand2 _6546_ (
    .a(\DFF_913.Q ),
    .b(\DFF_1428.Q ),
    .y(_2116_)
  );
  al_aoi21ttf _6547_ (
    .a(\DFF_914.Q ),
    .b(\DFF_1429.Q ),
    .c(_2116_),
    .y(_2117_)
  );
  al_ao21 _6548_ (
    .a(_2115_),
    .b(_2117_),
    .c(\DFF_1008.D ),
    .y(_2118_)
  );
  al_and3 _6549_ (
    .a(\DFF_1008.D ),
    .b(_2115_),
    .c(_2117_),
    .y(_2119_)
  );
  al_nand2ft _6550_ (
    .a(_2119_),
    .b(_2118_),
    .y(_2120_)
  );
  al_nand3ftt _6551_ (
    .a(_2114_),
    .b(_2113_),
    .c(_2120_),
    .y(_2121_)
  );
  al_nand2 _6552_ (
    .a(\DFF_921.Q ),
    .b(\DFF_1427.Q ),
    .y(_2122_)
  );
  al_nand2 _6553_ (
    .a(\DFF_922.Q ),
    .b(\DFF_1428.Q ),
    .y(_2123_)
  );
  al_aoi21ttf _6554_ (
    .a(\DFF_923.Q ),
    .b(\DFF_1429.Q ),
    .c(_2123_),
    .y(_2124_)
  );
  al_aoi21 _6555_ (
    .a(_2122_),
    .b(_2124_),
    .c(\DFF_40.Q ),
    .y(_2125_)
  );
  al_and3 _6556_ (
    .a(\DFF_40.Q ),
    .b(_2122_),
    .c(_2124_),
    .y(_2126_)
  );
  al_nand2 _6557_ (
    .a(\DFF_915.Q ),
    .b(\DFF_1427.Q ),
    .y(_2127_)
  );
  al_nand2 _6558_ (
    .a(\DFF_916.Q ),
    .b(\DFF_1428.Q ),
    .y(_2128_)
  );
  al_aoi21ttf _6559_ (
    .a(\DFF_917.Q ),
    .b(\DFF_1429.Q ),
    .c(_2128_),
    .y(_2129_)
  );
  al_ao21 _6560_ (
    .a(_2127_),
    .b(_2129_),
    .c(\DFF_1006.D ),
    .y(_2130_)
  );
  al_and3 _6561_ (
    .a(\DFF_1006.D ),
    .b(_2127_),
    .c(_2129_),
    .y(_2131_)
  );
  al_nand2ft _6562_ (
    .a(_2131_),
    .b(_2130_),
    .y(_2132_)
  );
  al_nand3fft _6563_ (
    .a(_2125_),
    .b(_2126_),
    .c(_2132_),
    .y(_2133_)
  );
  al_nand2 _6564_ (
    .a(\DFF_927.Q ),
    .b(\DFF_1427.Q ),
    .y(_2134_)
  );
  al_nand2 _6565_ (
    .a(\DFF_928.Q ),
    .b(\DFF_1428.Q ),
    .y(_2135_)
  );
  al_aoi21ttf _6566_ (
    .a(\DFF_929.Q ),
    .b(\DFF_1429.Q ),
    .c(_2135_),
    .y(_2136_)
  );
  al_ao21 _6567_ (
    .a(_2134_),
    .b(_2136_),
    .c(\DFF_998.D ),
    .y(_2137_)
  );
  al_and3 _6568_ (
    .a(\DFF_998.D ),
    .b(_2134_),
    .c(_2136_),
    .y(_2138_)
  );
  al_nand2ft _6569_ (
    .a(_2138_),
    .b(_2137_),
    .y(_2139_)
  );
  al_nand2 _6570_ (
    .a(\DFF_933.Q ),
    .b(\DFF_1427.Q ),
    .y(_2140_)
  );
  al_nand2 _6571_ (
    .a(\DFF_934.Q ),
    .b(\DFF_1428.Q ),
    .y(_2141_)
  );
  al_aoi21ttf _6572_ (
    .a(\DFF_935.Q ),
    .b(\DFF_1429.Q ),
    .c(_2141_),
    .y(_2142_)
  );
  al_nand2 _6573_ (
    .a(_2140_),
    .b(_2142_),
    .y(_2143_)
  );
  al_nand3fft _6574_ (
    .a(_0215_),
    .b(_0217_),
    .c(_2143_),
    .y(_2144_)
  );
  al_nand3 _6575_ (
    .a(_2140_),
    .b(_2142_),
    .c(_1833_),
    .y(_2145_)
  );
  al_and3 _6576_ (
    .a(_2144_),
    .b(_2145_),
    .c(_2139_),
    .y(_2146_)
  );
  al_and3fft _6577_ (
    .a(_2133_),
    .b(_2121_),
    .c(_2146_),
    .y(_2147_)
  );
  al_ao21 _6578_ (
    .a(_2109_),
    .b(_2147_),
    .c(_2084_),
    .y(_2148_)
  );
  al_aoi21ftf _6579_ (
    .a(_0308_),
    .b(_2148_),
    .c(_0156_),
    .y(_2149_)
  );
  al_nand2ft _6580_ (
    .a(_0304_),
    .b(_0306_),
    .y(_2150_)
  );
  al_and2ft _6581_ (
    .a(_2101_),
    .b(_2100_),
    .y(_2151_)
  );
  al_nor3fft _6582_ (
    .a(_2151_),
    .b(_2133_),
    .c(_2146_),
    .y(_2152_)
  );
  al_nand2 _6583_ (
    .a(_2145_),
    .b(_2144_),
    .y(_2153_)
  );
  al_nand3fft _6584_ (
    .a(_2125_),
    .b(_2126_),
    .c(_2139_),
    .y(_2154_)
  );
  al_aoi21ftf _6585_ (
    .a(_2131_),
    .b(_2130_),
    .c(_2102_),
    .y(_2155_)
  );
  al_or3fft _6586_ (
    .a(_2153_),
    .b(_2154_),
    .c(_2155_),
    .y(_2156_)
  );
  al_or2 _6587_ (
    .a(_2126_),
    .b(_2125_),
    .y(_2157_)
  );
  al_nand3 _6588_ (
    .a(_2144_),
    .b(_2145_),
    .c(_2132_),
    .y(_2158_)
  );
  al_ao21ftf _6589_ (
    .a(_2138_),
    .b(_2137_),
    .c(_2102_),
    .y(_2159_)
  );
  al_nand3 _6590_ (
    .a(_2157_),
    .b(_2158_),
    .c(_2159_),
    .y(_2160_)
  );
  al_and3ftt _6591_ (
    .a(_2152_),
    .b(_2156_),
    .c(_2160_),
    .y(_2161_)
  );
  al_or3fft _6592_ (
    .a(\DFF_1302.Q ),
    .b(_1005_),
    .c(_2161_),
    .y(_2162_)
  );
  al_and2ft _6593_ (
    .a(_2089_),
    .b(_2088_),
    .y(_2163_)
  );
  al_ao21ftf _6594_ (
    .a(_2094_),
    .b(_2093_),
    .c(_2108_),
    .y(_2164_)
  );
  al_nand3ftt _6595_ (
    .a(_2163_),
    .b(_2121_),
    .c(_2164_),
    .y(_2165_)
  );
  al_ao21 _6596_ (
    .a(_2120_),
    .b(_2163_),
    .c(_2108_),
    .y(_2166_)
  );
  al_nand2ft _6597_ (
    .a(_2114_),
    .b(_2113_),
    .y(_2167_)
  );
  al_ao21ttf _6598_ (
    .a(_2095_),
    .b(_2163_),
    .c(_2167_),
    .y(_2168_)
  );
  al_nand3fft _6599_ (
    .a(_2106_),
    .b(_2107_),
    .c(_2120_),
    .y(_2169_)
  );
  al_aoi21ftf _6600_ (
    .a(_2167_),
    .b(_2095_),
    .c(_2169_),
    .y(_2170_)
  );
  al_ao21ttf _6601_ (
    .a(_2166_),
    .b(_2168_),
    .c(_2170_),
    .y(_2171_)
  );
  al_ao21 _6602_ (
    .a(_2165_),
    .b(_2171_),
    .c(_1006_),
    .y(_2172_)
  );
  al_and3 _6603_ (
    .a(_0301_),
    .b(_2172_),
    .c(_2162_),
    .y(_2173_)
  );
  al_inv _6604_ (
    .a(_0298_),
    .y(_2174_)
  );
  al_nand2 _6605_ (
    .a(_2174_),
    .b(_1010_),
    .y(_2175_)
  );
  al_oai21ftf _6606_ (
    .a(_2150_),
    .b(_2173_),
    .c(_2175_),
    .y(_2176_)
  );
  al_mux2h _6607_ (
    .a(\DFF_992.Q ),
    .b(_2176_),
    .s(_2149_),
    .y(\DFF_992.D )
  );
  al_aoi21ftf _6608_ (
    .a(_0308_),
    .b(_2148_),
    .c(_0157_),
    .y(_2177_)
  );
  al_mux2h _6609_ (
    .a(\DFF_993.Q ),
    .b(_2176_),
    .s(_2177_),
    .y(\DFF_993.D )
  );
  al_aoi21ftf _6610_ (
    .a(_0308_),
    .b(_2148_),
    .c(_0158_),
    .y(_2178_)
  );
  al_mux2h _6611_ (
    .a(\DFF_994.Q ),
    .b(_2176_),
    .s(_2178_),
    .y(\DFF_994.D )
  );
  al_inv _6612_ (
    .a(_0222_),
    .y(\DFF_1016.D )
  );
  al_and3fft _6613_ (
    .a(_1102_),
    .b(_1005_),
    .c(_0222_),
    .y(_2179_)
  );
  al_oai21ftt _6614_ (
    .a(_1832_),
    .b(_2179_),
    .c(_1844_),
    .y(_2180_)
  );
  al_oai21ftf _6615_ (
    .a(_1835_),
    .b(_1836_),
    .c(_2180_),
    .y(_2181_)
  );
  al_nand3 _6616_ (
    .a(_2179_),
    .b(_1840_),
    .c(_1834_),
    .y(_2182_)
  );
  al_and3 _6617_ (
    .a(\DFF_1016.D ),
    .b(_2182_),
    .c(_2181_),
    .y(_2183_)
  );
  al_ao21 _6618_ (
    .a(_2182_),
    .b(_2181_),
    .c(\DFF_1016.D ),
    .y(_2184_)
  );
  al_nand2ft _6619_ (
    .a(_2183_),
    .b(_2184_),
    .y(_2185_)
  );
  al_mux2h _6620_ (
    .a(\DFF_968.Q ),
    .b(_2185_),
    .s(\DFF_1427.Q ),
    .y(\DFF_968.D )
  );
  al_mux2h _6621_ (
    .a(\DFF_969.Q ),
    .b(_2185_),
    .s(\DFF_1428.Q ),
    .y(\DFF_969.D )
  );
  al_mux2h _6622_ (
    .a(\DFF_970.Q ),
    .b(_2185_),
    .s(\DFF_1429.Q ),
    .y(\DFF_970.D )
  );
  al_nand3 _6623_ (
    .a(\DFF_1293.Q ),
    .b(\DFF_1294.Q ),
    .c(_1683_),
    .y(_2186_)
  );
  al_ao21 _6624_ (
    .a(\DFF_1293.Q ),
    .b(_1683_),
    .c(\DFF_1294.Q ),
    .y(_2187_)
  );
  al_and3 _6625_ (
    .a(_0778_),
    .b(_2186_),
    .c(_2187_),
    .y(\DFF_1294.D )
  );
  al_nand2 _6626_ (
    .a(\DFF_1281.Q ),
    .b(\DFF_1428.Q ),
    .y(_2188_)
  );
  al_aoi21ttf _6627_ (
    .a(\DFF_1282.Q ),
    .b(\DFF_1429.Q ),
    .c(_2188_),
    .y(_2189_)
  );
  al_ao21ftf _6628_ (
    .a(_1197_),
    .b(\DFF_1280.Q ),
    .c(_2189_),
    .y(_2190_)
  );
  al_and2ft _6629_ (
    .a(_0236_),
    .b(_2190_),
    .y(_2191_)
  );
  al_nor2ft _6630_ (
    .a(_0236_),
    .b(_2190_),
    .y(_2192_)
  );
  al_nand2 _6631_ (
    .a(\DFF_1274.Q ),
    .b(\DFF_1427.Q ),
    .y(_2193_)
  );
  al_nand2 _6632_ (
    .a(\DFF_1275.Q ),
    .b(\DFF_1428.Q ),
    .y(_2194_)
  );
  al_aoi21ttf _6633_ (
    .a(\DFF_1276.Q ),
    .b(\DFF_1429.Q ),
    .c(_2194_),
    .y(_2195_)
  );
  al_ao21 _6634_ (
    .a(_2193_),
    .b(_2195_),
    .c(\DFF_1350.D ),
    .y(_2196_)
  );
  al_and3 _6635_ (
    .a(\DFF_1350.D ),
    .b(_2193_),
    .c(_2195_),
    .y(_2197_)
  );
  al_nand2ft _6636_ (
    .a(_2197_),
    .b(_2196_),
    .y(_2198_)
  );
  al_and3fft _6637_ (
    .a(_2191_),
    .b(_2192_),
    .c(_2198_),
    .y(_2199_)
  );
  al_nand2 _6638_ (
    .a(\DFF_1260.Q ),
    .b(\DFF_1428.Q ),
    .y(_2200_)
  );
  al_aoi21ttf _6639_ (
    .a(\DFF_1261.Q ),
    .b(\DFF_1429.Q ),
    .c(_2200_),
    .y(_2201_)
  );
  al_ao21ftf _6640_ (
    .a(_1197_),
    .b(\DFF_1259.Q ),
    .c(_2201_),
    .y(_2202_)
  );
  al_and2 _6641_ (
    .a(\DFF_1360.D ),
    .b(_2202_),
    .y(_2203_)
  );
  al_aoi21ftf _6642_ (
    .a(_1197_),
    .b(\DFF_1259.Q ),
    .c(_2201_),
    .y(_2204_)
  );
  al_and2 _6643_ (
    .a(\DFF_89.Q ),
    .b(_2204_),
    .y(_2205_)
  );
  al_nor2 _6644_ (
    .a(_2203_),
    .b(_2205_),
    .y(_2206_)
  );
  al_nand2 _6645_ (
    .a(\DFF_1257.Q ),
    .b(\DFF_1428.Q ),
    .y(_2207_)
  );
  al_aoi21ttf _6646_ (
    .a(\DFF_1258.Q ),
    .b(\DFF_1429.Q ),
    .c(_2207_),
    .y(_2208_)
  );
  al_ao21ftf _6647_ (
    .a(_1197_),
    .b(\DFF_1256.Q ),
    .c(_2208_),
    .y(_2209_)
  );
  al_and2 _6648_ (
    .a(\DFF_90.Q ),
    .b(_2209_),
    .y(_2210_)
  );
  al_aoi21ftf _6649_ (
    .a(_1197_),
    .b(\DFF_1256.Q ),
    .c(_2208_),
    .y(_2211_)
  );
  al_nand2 _6650_ (
    .a(\DFF_1362.D ),
    .b(_2211_),
    .y(_2212_)
  );
  al_nand2ft _6651_ (
    .a(_2210_),
    .b(_2212_),
    .y(_2213_)
  );
  al_and3 _6652_ (
    .a(_2213_),
    .b(_2206_),
    .c(_2199_),
    .y(_2214_)
  );
  al_nand2 _6653_ (
    .a(\DFF_1269.Q ),
    .b(\DFF_1428.Q ),
    .y(_2215_)
  );
  al_aoi21ttf _6654_ (
    .a(\DFF_1270.Q ),
    .b(\DFF_1429.Q ),
    .c(_2215_),
    .y(_2216_)
  );
  al_ao21ftf _6655_ (
    .a(_1197_),
    .b(\DFF_1268.Q ),
    .c(_2216_),
    .y(_2217_)
  );
  al_and2 _6656_ (
    .a(\DFF_86.Q ),
    .b(_2217_),
    .y(_2218_)
  );
  al_or2 _6657_ (
    .a(\DFF_86.Q ),
    .b(_2217_),
    .y(_2219_)
  );
  al_nand2 _6658_ (
    .a(\DFF_1262.Q ),
    .b(\DFF_1427.Q ),
    .y(_2220_)
  );
  al_nand2 _6659_ (
    .a(\DFF_1263.Q ),
    .b(\DFF_1428.Q ),
    .y(_2221_)
  );
  al_aoi21ttf _6660_ (
    .a(\DFF_1264.Q ),
    .b(\DFF_1429.Q ),
    .c(_2221_),
    .y(_2222_)
  );
  al_ao21 _6661_ (
    .a(_2220_),
    .b(_2222_),
    .c(\DFF_1358.D ),
    .y(_2223_)
  );
  al_and3 _6662_ (
    .a(\DFF_1358.D ),
    .b(_2220_),
    .c(_2222_),
    .y(_2224_)
  );
  al_nand2ft _6663_ (
    .a(_2224_),
    .b(_2223_),
    .y(_2225_)
  );
  al_oa21ftt _6664_ (
    .a(_2219_),
    .b(_2218_),
    .c(_2225_),
    .y(_2226_)
  );
  al_nand2 _6665_ (
    .a(\DFF_1265.Q ),
    .b(\DFF_1427.Q ),
    .y(_2227_)
  );
  al_nand2 _6666_ (
    .a(\DFF_1266.Q ),
    .b(\DFF_1428.Q ),
    .y(_2228_)
  );
  al_aoi21ttf _6667_ (
    .a(\DFF_1267.Q ),
    .b(\DFF_1429.Q ),
    .c(_2228_),
    .y(_2229_)
  );
  al_ao21 _6668_ (
    .a(_2227_),
    .b(_2229_),
    .c(\DFF_1356.D ),
    .y(_2230_)
  );
  al_and3 _6669_ (
    .a(\DFF_1356.D ),
    .b(_2227_),
    .c(_2229_),
    .y(_2231_)
  );
  al_nand2ft _6670_ (
    .a(_2231_),
    .b(_2230_),
    .y(_2232_)
  );
  al_nand2 _6671_ (
    .a(\DFF_1272.Q ),
    .b(\DFF_1428.Q ),
    .y(_2233_)
  );
  al_aoi21ttf _6672_ (
    .a(\DFF_1273.Q ),
    .b(\DFF_1429.Q ),
    .c(_2233_),
    .y(_2234_)
  );
  al_aoi21ftf _6673_ (
    .a(_1197_),
    .b(\DFF_1271.Q ),
    .c(_2234_),
    .y(_2235_)
  );
  al_nor2 _6674_ (
    .a(\DFF_85.Q ),
    .b(_2235_),
    .y(_2236_)
  );
  al_and2 _6675_ (
    .a(\DFF_85.Q ),
    .b(_2235_),
    .y(_2237_)
  );
  al_nor2 _6676_ (
    .a(_2237_),
    .b(_2236_),
    .y(_2238_)
  );
  al_nand2 _6677_ (
    .a(\DFF_1277.Q ),
    .b(\DFF_1427.Q ),
    .y(_2239_)
  );
  al_nand2 _6678_ (
    .a(\DFF_1278.Q ),
    .b(\DFF_1428.Q ),
    .y(_2240_)
  );
  al_aoi21ttf _6679_ (
    .a(\DFF_1279.Q ),
    .b(\DFF_1429.Q ),
    .c(_2240_),
    .y(_2241_)
  );
  al_ao21 _6680_ (
    .a(_2239_),
    .b(_2241_),
    .c(\DFF_1348.D ),
    .y(_2242_)
  );
  al_and3 _6681_ (
    .a(\DFF_1348.D ),
    .b(_2239_),
    .c(_2241_),
    .y(_2243_)
  );
  al_nand2ft _6682_ (
    .a(_2243_),
    .b(_2242_),
    .y(_2244_)
  );
  al_nand2 _6683_ (
    .a(\DFF_1283.Q ),
    .b(\DFF_1427.Q ),
    .y(_2245_)
  );
  al_nand2 _6684_ (
    .a(\DFF_1284.Q ),
    .b(\DFF_1428.Q ),
    .y(_2246_)
  );
  al_aoi21ttf _6685_ (
    .a(\DFF_1285.Q ),
    .b(\DFF_1429.Q ),
    .c(_2246_),
    .y(_2247_)
  );
  al_ao21 _6686_ (
    .a(_2245_),
    .b(_2247_),
    .c(_0240_),
    .y(_2248_)
  );
  al_and3 _6687_ (
    .a(_2245_),
    .b(_2247_),
    .c(_0240_),
    .y(_2249_)
  );
  al_and3ftt _6688_ (
    .a(_2249_),
    .b(_2248_),
    .c(_2244_),
    .y(_2250_)
  );
  al_and3 _6689_ (
    .a(_2232_),
    .b(_2250_),
    .c(_2238_),
    .y(_2251_)
  );
  al_nand3 _6690_ (
    .a(_2226_),
    .b(_2251_),
    .c(_2214_),
    .y(_2252_)
  );
  al_ao21 _6691_ (
    .a(_1084_),
    .b(_2252_),
    .c(_0323_),
    .y(_2253_)
  );
  al_and2 _6692_ (
    .a(_0156_),
    .b(_2253_),
    .y(_2254_)
  );
  al_or2 _6693_ (
    .a(_0320_),
    .b(_0317_),
    .y(_2255_)
  );
  al_nand2 _6694_ (
    .a(\DFF_1302.Q ),
    .b(_1084_),
    .y(_2256_)
  );
  al_and3ftt _6695_ (
    .a(_2249_),
    .b(_2248_),
    .c(_2232_),
    .y(_2257_)
  );
  al_ao21 _6696_ (
    .a(_2244_),
    .b(_2206_),
    .c(_2238_),
    .y(_2258_)
  );
  al_and2ft _6697_ (
    .a(_2249_),
    .b(_2248_),
    .y(_2259_)
  );
  al_nand3fft _6698_ (
    .a(_2237_),
    .b(_2236_),
    .c(_2244_),
    .y(_2260_)
  );
  al_nand3fft _6699_ (
    .a(_2203_),
    .b(_2205_),
    .c(_2232_),
    .y(_2261_)
  );
  al_nand3ftt _6700_ (
    .a(_2259_),
    .b(_2260_),
    .c(_2261_),
    .y(_2262_)
  );
  al_ao21 _6701_ (
    .a(_2258_),
    .b(_2262_),
    .c(_2257_),
    .y(_2263_)
  );
  al_and3fft _6702_ (
    .a(_2236_),
    .b(_2237_),
    .c(_2232_),
    .y(_2264_)
  );
  al_or3 _6703_ (
    .a(_2250_),
    .b(_2206_),
    .c(_2264_),
    .y(_2265_)
  );
  al_ao21 _6704_ (
    .a(_2265_),
    .b(_2263_),
    .c(_2256_),
    .y(_2266_)
  );
  al_nand2ft _6705_ (
    .a(_2218_),
    .b(_2219_),
    .y(_2267_)
  );
  al_ao21 _6706_ (
    .a(_2198_),
    .b(_2213_),
    .c(_2267_),
    .y(_2268_)
  );
  al_oai21ftt _6707_ (
    .a(_2212_),
    .b(_2210_),
    .c(_2225_),
    .y(_2269_)
  );
  al_oai21 _6708_ (
    .a(_2191_),
    .b(_2192_),
    .c(_2269_),
    .y(_2270_)
  );
  al_nand3fft _6709_ (
    .a(_2191_),
    .b(_2192_),
    .c(_2225_),
    .y(_2271_)
  );
  al_aoi21ttf _6710_ (
    .a(_2198_),
    .b(_2267_),
    .c(_2271_),
    .y(_2272_)
  );
  al_ao21ttf _6711_ (
    .a(_2270_),
    .b(_2268_),
    .c(_2272_),
    .y(_2273_)
  );
  al_or3 _6712_ (
    .a(_2213_),
    .b(_2226_),
    .c(_2199_),
    .y(_2274_)
  );
  al_ao21 _6713_ (
    .a(_2274_),
    .b(_2273_),
    .c(_2256_),
    .y(_2275_)
  );
  al_and3 _6714_ (
    .a(_0317_),
    .b(_2275_),
    .c(_2266_),
    .y(_2276_)
  );
  al_nand2 _6715_ (
    .a(_0314_),
    .b(_1088_),
    .y(_2277_)
  );
  al_oai21ftf _6716_ (
    .a(_2255_),
    .b(_2276_),
    .c(_2277_),
    .y(_2278_)
  );
  al_mux2h _6717_ (
    .a(\DFF_1342.Q ),
    .b(_2278_),
    .s(_2254_),
    .y(\DFF_1342.D )
  );
  al_and2 _6718_ (
    .a(_0157_),
    .b(_2253_),
    .y(_2279_)
  );
  al_mux2h _6719_ (
    .a(\DFF_1343.Q ),
    .b(_2278_),
    .s(_2279_),
    .y(\DFF_1343.D )
  );
  al_and2 _6720_ (
    .a(_0158_),
    .b(_2253_),
    .y(_2280_)
  );
  al_mux2h _6721_ (
    .a(\DFF_1344.Q ),
    .b(_2278_),
    .s(_2280_),
    .y(\DFF_1344.D )
  );
  al_inv _6722_ (
    .a(_0245_),
    .y(\DFF_1366.D )
  );
  al_and3fft _6723_ (
    .a(_1102_),
    .b(_1084_),
    .c(_0245_),
    .y(_2281_)
  );
  al_oai21ftt _6724_ (
    .a(_1862_),
    .b(_2281_),
    .c(_1873_),
    .y(_2282_)
  );
  al_oai21ftf _6725_ (
    .a(_1864_),
    .b(_1866_),
    .c(_2282_),
    .y(_2283_)
  );
  al_nand3 _6726_ (
    .a(_2281_),
    .b(_1869_),
    .c(_1863_),
    .y(_2284_)
  );
  al_and3 _6727_ (
    .a(\DFF_1366.D ),
    .b(_2284_),
    .c(_2283_),
    .y(_2285_)
  );
  al_ao21 _6728_ (
    .a(_2284_),
    .b(_2283_),
    .c(\DFF_1366.D ),
    .y(_2286_)
  );
  al_nand2ft _6729_ (
    .a(_2285_),
    .b(_2286_),
    .y(_2287_)
  );
  al_mux2h _6730_ (
    .a(\DFF_1318.Q ),
    .b(_2287_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1318.D )
  );
  al_mux2h _6731_ (
    .a(\DFF_1319.Q ),
    .b(_2287_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1319.D )
  );
  al_mux2h _6732_ (
    .a(\DFF_1320.Q ),
    .b(_2287_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1320.D )
  );
  al_nand3ftt _6733_ (
    .a(\DFF_160.Q ),
    .b(_1450_),
    .c(_1452_),
    .y(_2288_)
  );
  al_nand3fft _6734_ (
    .a(\DFF_1624.Q ),
    .b(\DFF_1634.Q ),
    .c(_1762_),
    .y(_2289_)
  );
  al_nand2ft _6735_ (
    .a(\DFF_160.Q ),
    .b(_1764_),
    .y(_2290_)
  );
  al_ao21ttf _6736_ (
    .a(_2290_),
    .b(_2289_),
    .c(_1769_),
    .y(_2291_)
  );
  al_nand2 _6737_ (
    .a(_1751_),
    .b(_1452_),
    .y(_2292_)
  );
  al_nor3fft _6738_ (
    .a(_1449_),
    .b(_2292_),
    .c(_1752_),
    .y(_2293_)
  );
  al_and3 _6739_ (
    .a(_2291_),
    .b(_2288_),
    .c(_2293_),
    .y(\DFF_160.D )
  );
  al_inv _6740_ (
    .a(\DFF_160.D ),
    .y(\DFF_157.D )
  );
  al_aoi21ftf _6741_ (
    .a(\DFF_245.Q ),
    .b(_1878_),
    .c(_0778_),
    .y(_2294_)
  );
  al_aoi21ftf _6742_ (
    .a(_1878_),
    .b(\DFF_245.Q ),
    .c(_2294_),
    .y(\DFF_245.D )
  );
  al_nand3ftt _6743_ (
    .a(_0267_),
    .b(_0273_),
    .c(_0270_),
    .y(_2295_)
  );
  al_ao21ftt _6744_ (
    .a(_1954_),
    .b(_1951_),
    .c(_0848_),
    .y(_2296_)
  );
  al_oai21 _6745_ (
    .a(_0273_),
    .b(_0270_),
    .c(_0267_),
    .y(_2297_)
  );
  al_ao21 _6746_ (
    .a(_2296_),
    .b(_1965_),
    .c(_2297_),
    .y(_2298_)
  );
  al_and2 _6747_ (
    .a(_0783_),
    .b(_0851_),
    .y(_2299_)
  );
  al_aoi21 _6748_ (
    .a(_2295_),
    .b(_2298_),
    .c(_2299_),
    .y(_2300_)
  );
  al_mux2h _6749_ (
    .a(\DFF_283.Q ),
    .b(_2300_),
    .s(\DFF_1427.Q ),
    .y(\DFF_283.D )
  );
  al_mux2h _6750_ (
    .a(\DFF_284.Q ),
    .b(_2300_),
    .s(\DFF_1428.Q ),
    .y(\DFF_284.D )
  );
  al_mux2h _6751_ (
    .a(\DFF_285.Q ),
    .b(_2300_),
    .s(\DFF_1429.Q ),
    .y(\DFF_285.D )
  );
  al_aoi21ftf _6752_ (
    .a(\DFF_595.Q ),
    .b(_1974_),
    .c(_0778_),
    .y(_2301_)
  );
  al_aoi21ftf _6753_ (
    .a(_1974_),
    .b(\DFF_595.Q ),
    .c(_2301_),
    .y(\DFF_595.D )
  );
  al_nand3 _6754_ (
    .a(_0287_),
    .b(_0281_),
    .c(_0284_),
    .y(_2302_)
  );
  al_oai21ttf _6755_ (
    .a(_0287_),
    .b(_0284_),
    .c(_0281_),
    .y(_2303_)
  );
  al_ao21 _6756_ (
    .a(_2061_),
    .b(_2049_),
    .c(_2303_),
    .y(_2304_)
  );
  al_and2 _6757_ (
    .a(_0863_),
    .b(_2074_),
    .y(_2305_)
  );
  al_aoi21 _6758_ (
    .a(_2302_),
    .b(_2304_),
    .c(_2305_),
    .y(_2306_)
  );
  al_mux2h _6759_ (
    .a(\DFF_633.Q ),
    .b(_2306_),
    .s(\DFF_1427.Q ),
    .y(\DFF_633.D )
  );
  al_mux2h _6760_ (
    .a(\DFF_634.Q ),
    .b(_2306_),
    .s(\DFF_1428.Q ),
    .y(\DFF_634.D )
  );
  al_mux2h _6761_ (
    .a(\DFF_635.Q ),
    .b(_2306_),
    .s(\DFF_1429.Q ),
    .y(\DFF_635.D )
  );
  al_aoi21ftf _6762_ (
    .a(\DFF_945.Q ),
    .b(_2082_),
    .c(_0778_),
    .y(_2307_)
  );
  al_aoi21ftf _6763_ (
    .a(_2082_),
    .b(\DFF_945.Q ),
    .c(_2307_),
    .y(\DFF_945.D )
  );
  al_nand3 _6764_ (
    .a(_0298_),
    .b(_0304_),
    .c(_0301_),
    .y(_2308_)
  );
  al_oai21ftf _6765_ (
    .a(_0306_),
    .b(_0304_),
    .c(_0298_),
    .y(_2309_)
  );
  al_ao21 _6766_ (
    .a(_2172_),
    .b(_2162_),
    .c(_2309_),
    .y(_2310_)
  );
  al_and2 _6767_ (
    .a(_0978_),
    .b(_0977_),
    .y(_2311_)
  );
  al_or2ft _6768_ (
    .a(_1002_),
    .b(_1001_),
    .y(_2312_)
  );
  al_and3fft _6769_ (
    .a(_1006_),
    .b(_0952_),
    .c(_0951_),
    .y(_2313_)
  );
  al_and3ftt _6770_ (
    .a(_2312_),
    .b(_2311_),
    .c(_2313_),
    .y(_2314_)
  );
  al_and3 _6771_ (
    .a(_0973_),
    .b(_0997_),
    .c(_0991_),
    .y(_2315_)
  );
  al_and3fft _6772_ (
    .a(_0945_),
    .b(_0946_),
    .c(_0984_),
    .y(_2316_)
  );
  al_and3 _6773_ (
    .a(_0966_),
    .b(_2316_),
    .c(_2315_),
    .y(_2317_)
  );
  al_and3 _6774_ (
    .a(_0941_),
    .b(_2314_),
    .c(_2317_),
    .y(_2318_)
  );
  al_aoi21 _6775_ (
    .a(_2308_),
    .b(_2310_),
    .c(_2318_),
    .y(_2319_)
  );
  al_mux2h _6776_ (
    .a(\DFF_983.Q ),
    .b(_2319_),
    .s(\DFF_1427.Q ),
    .y(\DFF_983.D )
  );
  al_mux2h _6777_ (
    .a(\DFF_984.Q ),
    .b(_2319_),
    .s(\DFF_1428.Q ),
    .y(\DFF_984.D )
  );
  al_mux2h _6778_ (
    .a(\DFF_985.Q ),
    .b(_2319_),
    .s(\DFF_1429.Q ),
    .y(\DFF_985.D )
  );
  al_aoi21ftf _6779_ (
    .a(\DFF_1295.Q ),
    .b(_2186_),
    .c(_0778_),
    .y(_2320_)
  );
  al_aoi21ftf _6780_ (
    .a(_2186_),
    .b(\DFF_1295.Q ),
    .c(_2320_),
    .y(\DFF_1295.D )
  );
  al_nand3ftt _6781_ (
    .a(_0314_),
    .b(_0320_),
    .c(_0317_),
    .y(_2321_)
  );
  al_oai21 _6782_ (
    .a(_0320_),
    .b(_0317_),
    .c(_0314_),
    .y(_2322_)
  );
  al_ao21 _6783_ (
    .a(_2275_),
    .b(_2266_),
    .c(_2322_),
    .y(_2323_)
  );
  al_and2 _6784_ (
    .a(_1018_),
    .b(_1088_),
    .y(_2324_)
  );
  al_aoi21 _6785_ (
    .a(_2321_),
    .b(_2323_),
    .c(_2324_),
    .y(_2325_)
  );
  al_mux2h _6786_ (
    .a(\DFF_1333.Q ),
    .b(_2325_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1333.D )
  );
  al_mux2h _6787_ (
    .a(\DFF_1334.Q ),
    .b(_2325_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1334.D )
  );
  al_mux2h _6788_ (
    .a(\DFF_1335.Q ),
    .b(_2325_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1335.D )
  );
  al_nand3fft _6789_ (
    .a(_0025_),
    .b(_1851_),
    .c(_1853_),
    .y(_2326_)
  );
  al_ao21ftf _6790_ (
    .a(\DFF_1504.Q ),
    .b(\DFF_113.Q ),
    .c(_2326_),
    .y(\DFF_113.D )
  );
  al_mux2h _6791_ (
    .a(\DFF_114.Q ),
    .b(\DFF_1100.D ),
    .s(\DFF_1505.Q ),
    .y(\DFF_114.D )
  );
  al_mux2h _6792_ (
    .a(\DFF_115.Q ),
    .b(\DFF_1100.D ),
    .s(\DFF_1506.Q ),
    .y(\DFF_115.D )
  );
  al_oa21ftt _6793_ (
    .a(\DFF_1367.Q ),
    .b(\DFF_1428.Q ),
    .c(\DFF_1366.Q ),
    .y(_2327_)
  );
  al_ao21ttf _6794_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_1017.D ),
    .c(_2327_),
    .y(_2328_)
  );
  al_aoi21ftf _6795_ (
    .a(\DFF_1366.Q ),
    .b(\DFF_1378.Q ),
    .c(_2328_),
    .y(\DFF_1367.D )
  );
  al_and2ft _6796_ (
    .a(\DFF_1483.Q ),
    .b(\DFF_1482.Q ),
    .y(_2329_)
  );
  al_nand3fft _6797_ (
    .a(_0353_),
    .b(_1848_),
    .c(_1850_),
    .y(_2330_)
  );
  al_oa21ftf _6798_ (
    .a(\DFF_1492.Q ),
    .b(\DFF_1505.Q ),
    .c(\DFF_1482.Q ),
    .y(_2331_)
  );
  al_aoi21 _6799_ (
    .a(_2331_),
    .b(_2330_),
    .c(_2329_),
    .y(\DFF_1492.D )
  );
  al_oa21ftf _6800_ (
    .a(\DFF_1450.Q ),
    .b(\DFF_1504.Q ),
    .c(\DFF_1452.Q ),
    .y(_2332_)
  );
  al_nand2 _6801_ (
    .a(_2332_),
    .b(_2326_),
    .y(_2333_)
  );
  al_ao21ftf _6802_ (
    .a(\DFF_1449.Q ),
    .b(\DFF_1452.Q ),
    .c(_2333_),
    .y(_2334_)
  );
  al_inv _6803_ (
    .a(_2334_),
    .y(\DFF_1450.D )
  );
  al_and3ftt _6804_ (
    .a(_0789_),
    .b(_0833_),
    .c(_0795_),
    .y(_2335_)
  );
  al_and3 _6805_ (
    .a(_0839_),
    .b(_0820_),
    .c(_2335_),
    .y(_2336_)
  );
  al_or2 _6806_ (
    .a(_0844_),
    .b(_0843_),
    .y(_2337_)
  );
  al_nor3fft _6807_ (
    .a(_0801_),
    .b(_0814_),
    .c(_2337_),
    .y(_2338_)
  );
  al_and3 _6808_ (
    .a(\DFF_1302.Q ),
    .b(_0847_),
    .c(_0806_),
    .y(_2339_)
  );
  al_and3ftt _6809_ (
    .a(_0805_),
    .b(_2339_),
    .c(_0826_),
    .y(_2340_)
  );
  al_and2 _6810_ (
    .a(_2338_),
    .b(_2340_),
    .y(_2341_)
  );
  al_nand3 _6811_ (
    .a(_0783_),
    .b(_2336_),
    .c(_2341_),
    .y(_2342_)
  );
  al_or3fft _6812_ (
    .a(\DFF_1302.Q ),
    .b(_0267_),
    .c(_0847_),
    .y(_2343_)
  );
  al_and3 _6813_ (
    .a(_2338_),
    .b(_2340_),
    .c(_2336_),
    .y(_2344_)
  );
  al_nand2ft _6814_ (
    .a(\DFF_294.Q ),
    .b(\DFF_1429.Q ),
    .y(_2345_)
  );
  al_aoi21ftf _6815_ (
    .a(\DFF_293.Q ),
    .b(\DFF_1428.Q ),
    .c(_2345_),
    .y(_2346_)
  );
  al_ao21ftf _6816_ (
    .a(\DFF_292.Q ),
    .b(\DFF_1427.Q ),
    .c(_2346_),
    .y(_2347_)
  );
  al_nand3 _6817_ (
    .a(_0276_),
    .b(_2347_),
    .c(_2344_),
    .y(_2348_)
  );
  al_and3 _6818_ (
    .a(_2343_),
    .b(_2342_),
    .c(_2348_),
    .y(_2349_)
  );
  al_and2ft _6819_ (
    .a(_0273_),
    .b(_0270_),
    .y(_2350_)
  );
  al_and3 _6820_ (
    .a(_0267_),
    .b(_2347_),
    .c(_0851_),
    .y(_2351_)
  );
  al_nand3 _6821_ (
    .a(_2350_),
    .b(_2351_),
    .c(_1966_),
    .y(_2352_)
  );
  al_ao21 _6822_ (
    .a(_2349_),
    .b(_2352_),
    .c(\DFF_312.D ),
    .y(_2353_)
  );
  al_and2 _6823_ (
    .a(_1892_),
    .b(_1894_),
    .y(_2354_)
  );
  al_and2 _6824_ (
    .a(_1885_),
    .b(_1887_),
    .y(_2355_)
  );
  al_and3fft _6825_ (
    .a(_1900_),
    .b(_1931_),
    .c(_2355_),
    .y(_2356_)
  );
  al_and3 _6826_ (
    .a(_2354_),
    .b(_1882_),
    .c(_2356_),
    .y(_2357_)
  );
  al_nand2 _6827_ (
    .a(_1923_),
    .b(_1925_),
    .y(_2358_)
  );
  al_nand2 _6828_ (
    .a(_1904_),
    .b(_1906_),
    .y(_2359_)
  );
  al_nand2 _6829_ (
    .a(_1917_),
    .b(_1919_),
    .y(_2360_)
  );
  al_and2 _6830_ (
    .a(_1934_),
    .b(_1936_),
    .y(_2361_)
  );
  al_and3fft _6831_ (
    .a(_2359_),
    .b(_2360_),
    .c(_2361_),
    .y(_2362_)
  );
  al_nand3fft _6832_ (
    .a(_1912_),
    .b(_2358_),
    .c(_2362_),
    .y(_2363_)
  );
  al_nor3fft _6833_ (
    .a(_0275_),
    .b(_2357_),
    .c(_2363_),
    .y(_2364_)
  );
  al_and3 _6834_ (
    .a(_0273_),
    .b(_2360_),
    .c(_1198_),
    .y(_2365_)
  );
  al_aoi21ttf _6835_ (
    .a(_1934_),
    .b(_1936_),
    .c(_2358_),
    .y(_2366_)
  );
  al_and3 _6836_ (
    .a(_2359_),
    .b(_1912_),
    .c(_2366_),
    .y(_2367_)
  );
  al_and2 _6837_ (
    .a(_2367_),
    .b(_2357_),
    .y(_2368_)
  );
  al_aoi21 _6838_ (
    .a(_2365_),
    .b(_2368_),
    .c(_2364_),
    .y(_2369_)
  );
  al_and3 _6839_ (
    .a(_2349_),
    .b(_2369_),
    .c(_2352_),
    .y(_2370_)
  );
  al_ao21ftt _6840_ (
    .a(_0267_),
    .b(_0270_),
    .c(_2354_),
    .y(_2371_)
  );
  al_and3ftt _6841_ (
    .a(_0267_),
    .b(_0270_),
    .c(_2354_),
    .y(_2372_)
  );
  al_nand2ft _6842_ (
    .a(_2372_),
    .b(_2371_),
    .y(_2373_)
  );
  al_ao21ttf _6843_ (
    .a(_2373_),
    .b(_2370_),
    .c(_2353_),
    .y(_2374_)
  );
  al_mux2h _6844_ (
    .a(\DFF_206.Q ),
    .b(_2374_),
    .s(\DFF_1427.Q ),
    .y(\DFF_206.D )
  );
  al_mux2h _6845_ (
    .a(\DFF_207.Q ),
    .b(_2374_),
    .s(\DFF_1428.Q ),
    .y(\DFF_207.D )
  );
  al_mux2h _6846_ (
    .a(\DFF_208.Q ),
    .b(_2374_),
    .s(\DFF_1429.Q ),
    .y(\DFF_208.D )
  );
  al_ao21 _6847_ (
    .a(_2349_),
    .b(_2352_),
    .c(\DFF_304.D ),
    .y(_2375_)
  );
  al_nand2ft _6848_ (
    .a(_2360_),
    .b(_2295_),
    .y(_2376_)
  );
  al_nand2ft _6849_ (
    .a(_2365_),
    .b(_2376_),
    .y(_2377_)
  );
  al_and3ftt _6850_ (
    .a(_0267_),
    .b(_0273_),
    .c(_0270_),
    .y(_2378_)
  );
  al_mux2h _6851_ (
    .a(_2378_),
    .b(_0275_),
    .s(_2354_),
    .y(_2379_)
  );
  al_nand2 _6852_ (
    .a(_2361_),
    .b(_2295_),
    .y(_2380_)
  );
  al_and3ftt _6853_ (
    .a(_2361_),
    .b(_0273_),
    .c(_1198_),
    .y(_2381_)
  );
  al_aoi21ftf _6854_ (
    .a(_2381_),
    .b(_2380_),
    .c(_2379_),
    .y(_2382_)
  );
  al_nand2ft _6855_ (
    .a(_2359_),
    .b(_2295_),
    .y(_2383_)
  );
  al_and3 _6856_ (
    .a(_0273_),
    .b(_2359_),
    .c(_1198_),
    .y(_2384_)
  );
  al_aoi21ftf _6857_ (
    .a(_2384_),
    .b(_2383_),
    .c(_2382_),
    .y(_2385_)
  );
  al_ao21ttf _6858_ (
    .a(_2377_),
    .b(_2385_),
    .c(_1931_),
    .y(_2386_)
  );
  al_and3ftt _6859_ (
    .a(_1931_),
    .b(_2377_),
    .c(_2385_),
    .y(_2387_)
  );
  al_nand2ft _6860_ (
    .a(_2387_),
    .b(_2386_),
    .y(_2388_)
  );
  al_ao21ttf _6861_ (
    .a(_2388_),
    .b(_2370_),
    .c(_2375_),
    .y(_2389_)
  );
  al_mux2h _6862_ (
    .a(\DFF_218.Q ),
    .b(_2389_),
    .s(\DFF_1427.Q ),
    .y(\DFF_218.D )
  );
  al_mux2h _6863_ (
    .a(\DFF_219.Q ),
    .b(_2389_),
    .s(\DFF_1428.Q ),
    .y(\DFF_219.D )
  );
  al_mux2h _6864_ (
    .a(\DFF_220.Q ),
    .b(_2389_),
    .s(\DFF_1429.Q ),
    .y(\DFF_220.D )
  );
  al_ao21 _6865_ (
    .a(_2349_),
    .b(_2352_),
    .c(\DFF_300.D ),
    .y(_2390_)
  );
  al_nand2ft _6866_ (
    .a(_2384_),
    .b(_2383_),
    .y(_2391_)
  );
  al_and3 _6867_ (
    .a(_2377_),
    .b(_2391_),
    .c(_2382_),
    .y(_2392_)
  );
  al_and2ft _6868_ (
    .a(_1931_),
    .b(_2295_),
    .y(_2393_)
  );
  al_and3 _6869_ (
    .a(_0273_),
    .b(_1931_),
    .c(_1198_),
    .y(_2394_)
  );
  al_mux2h _6870_ (
    .a(_2394_),
    .b(_2393_),
    .s(_1882_),
    .y(_2395_)
  );
  al_ao21ttf _6871_ (
    .a(_2395_),
    .b(_2392_),
    .c(_1900_),
    .y(_2396_)
  );
  al_and3ftt _6872_ (
    .a(_1900_),
    .b(_2395_),
    .c(_2392_),
    .y(_2397_)
  );
  al_nand2ft _6873_ (
    .a(_2397_),
    .b(_2396_),
    .y(_2398_)
  );
  al_ao21ttf _6874_ (
    .a(_2398_),
    .b(_2370_),
    .c(_2390_),
    .y(_2399_)
  );
  al_mux2h _6875_ (
    .a(\DFF_224.Q ),
    .b(_2399_),
    .s(\DFF_1427.Q ),
    .y(\DFF_224.D )
  );
  al_mux2h _6876_ (
    .a(\DFF_225.Q ),
    .b(_2399_),
    .s(\DFF_1428.Q ),
    .y(\DFF_225.D )
  );
  al_mux2h _6877_ (
    .a(\DFF_226.Q ),
    .b(_2399_),
    .s(\DFF_1429.Q ),
    .y(\DFF_226.D )
  );
  al_ao21 _6878_ (
    .a(_2349_),
    .b(_2352_),
    .c(\DFF_302.D ),
    .y(_2400_)
  );
  al_or2 _6879_ (
    .a(_2394_),
    .b(_2393_),
    .y(_2401_)
  );
  al_ao21 _6880_ (
    .a(_2401_),
    .b(_2392_),
    .c(_1882_),
    .y(_2402_)
  );
  al_and3 _6881_ (
    .a(_1882_),
    .b(_2401_),
    .c(_2392_),
    .y(_2403_)
  );
  al_nand2ft _6882_ (
    .a(_2403_),
    .b(_2402_),
    .y(_2404_)
  );
  al_ao21ttf _6883_ (
    .a(_2404_),
    .b(_2370_),
    .c(_2400_),
    .y(_2405_)
  );
  al_mux2h _6884_ (
    .a(\DFF_221.Q ),
    .b(_2405_),
    .s(\DFF_1427.Q ),
    .y(\DFF_221.D )
  );
  al_mux2h _6885_ (
    .a(\DFF_222.Q ),
    .b(_2405_),
    .s(\DFF_1428.Q ),
    .y(\DFF_222.D )
  );
  al_mux2h _6886_ (
    .a(\DFF_223.Q ),
    .b(_2405_),
    .s(\DFF_1429.Q ),
    .y(\DFF_223.D )
  );
  al_ao21 _6887_ (
    .a(_2349_),
    .b(_2352_),
    .c(\DFF_298.D ),
    .y(_2406_)
  );
  al_and3 _6888_ (
    .a(_2377_),
    .b(_2395_),
    .c(_2385_),
    .y(_2407_)
  );
  al_nand2ft _6889_ (
    .a(_1900_),
    .b(_2295_),
    .y(_2408_)
  );
  al_and3 _6890_ (
    .a(_0273_),
    .b(_1900_),
    .c(_1198_),
    .y(_2409_)
  );
  al_nand2ft _6891_ (
    .a(_2409_),
    .b(_2408_),
    .y(_2410_)
  );
  al_and3 _6892_ (
    .a(_2355_),
    .b(_2410_),
    .c(_2407_),
    .y(_2411_)
  );
  al_ao21 _6893_ (
    .a(_2410_),
    .b(_2407_),
    .c(_2355_),
    .y(_2412_)
  );
  al_nand2ft _6894_ (
    .a(_2411_),
    .b(_2412_),
    .y(_2413_)
  );
  al_ao21ttf _6895_ (
    .a(_2413_),
    .b(_2370_),
    .c(_2406_),
    .y(_2414_)
  );
  al_mux2h _6896_ (
    .a(\DFF_227.Q ),
    .b(_2414_),
    .s(\DFF_1427.Q ),
    .y(\DFF_227.D )
  );
  al_mux2h _6897_ (
    .a(\DFF_228.Q ),
    .b(_2414_),
    .s(\DFF_1428.Q ),
    .y(\DFF_228.D )
  );
  al_mux2h _6898_ (
    .a(\DFF_229.Q ),
    .b(_2414_),
    .s(\DFF_1429.Q ),
    .y(\DFF_229.D )
  );
  al_or3fft _6899_ (
    .a(\DFF_1302.Q ),
    .b(_0926_),
    .c(_0281_),
    .y(_2415_)
  );
  al_nand2ft _6900_ (
    .a(\DFF_643.Q ),
    .b(\DFF_1428.Q ),
    .y(_2416_)
  );
  al_aoi21ftf _6901_ (
    .a(\DFF_644.Q ),
    .b(\DFF_1429.Q ),
    .c(_2416_),
    .y(_2417_)
  );
  al_ao21ftf _6902_ (
    .a(\DFF_642.Q ),
    .b(\DFF_1427.Q ),
    .c(_2417_),
    .y(_2418_)
  );
  al_nand3 _6903_ (
    .a(_0292_),
    .b(_2418_),
    .c(_2074_),
    .y(_2419_)
  );
  al_nor3fft _6904_ (
    .a(_2415_),
    .b(_2419_),
    .c(_2305_),
    .y(_2420_)
  );
  al_nand2ft _6905_ (
    .a(_0287_),
    .b(_0284_),
    .y(_2421_)
  );
  al_oa21 _6906_ (
    .a(_0874_),
    .b(_0873_),
    .c(_0888_),
    .y(_2422_)
  );
  al_and3fft _6907_ (
    .a(_2050_),
    .b(_2071_),
    .c(_2067_),
    .y(_2423_)
  );
  al_and3 _6908_ (
    .a(_2064_),
    .b(_2422_),
    .c(_2423_),
    .y(_2424_)
  );
  al_oai21 _6909_ (
    .a(_0868_),
    .b(_0867_),
    .c(_2072_),
    .y(_2425_)
  );
  al_nor3fft _6910_ (
    .a(_2068_),
    .b(_2070_),
    .c(_2425_),
    .y(_2426_)
  );
  al_and3 _6911_ (
    .a(_2418_),
    .b(_2426_),
    .c(_2424_),
    .y(_2427_)
  );
  al_nand3fft _6912_ (
    .a(_0281_),
    .b(_2421_),
    .c(_2427_),
    .y(_2428_)
  );
  al_or3fft _6913_ (
    .a(_2061_),
    .b(_2049_),
    .c(_2428_),
    .y(_2429_)
  );
  al_ao21 _6914_ (
    .a(_2420_),
    .b(_2429_),
    .c(\DFF_662.D ),
    .y(_2430_)
  );
  al_and2 _6915_ (
    .a(_0281_),
    .b(_0284_),
    .y(_2431_)
  );
  al_and2 _6916_ (
    .a(_1988_),
    .b(_1990_),
    .y(_2432_)
  );
  al_nand2 _6917_ (
    .a(_2025_),
    .b(_2027_),
    .y(_2433_)
  );
  al_and2 _6918_ (
    .a(_1976_),
    .b(_1978_),
    .y(_2434_)
  );
  al_nand2 _6919_ (
    .a(_1994_),
    .b(_1996_),
    .y(_2435_)
  );
  al_nand2 _6920_ (
    .a(_2031_),
    .b(_2033_),
    .y(_2436_)
  );
  al_and3fft _6921_ (
    .a(_2435_),
    .b(_2436_),
    .c(_2434_),
    .y(_2437_)
  );
  al_nand3ftt _6922_ (
    .a(_2433_),
    .b(_2432_),
    .c(_2437_),
    .y(_2438_)
  );
  al_nand2 _6923_ (
    .a(_2000_),
    .b(_2002_),
    .y(_2439_)
  );
  al_and2 _6924_ (
    .a(_2006_),
    .b(_2008_),
    .y(_2440_)
  );
  al_nand2 _6925_ (
    .a(_1982_),
    .b(_1984_),
    .y(_2441_)
  );
  al_and3fft _6926_ (
    .a(_2439_),
    .b(_2441_),
    .c(_2440_),
    .y(_2442_)
  );
  al_nand2 _6927_ (
    .a(_2013_),
    .b(_2015_),
    .y(_2443_)
  );
  al_nor3fft _6928_ (
    .a(_2019_),
    .b(_2021_),
    .c(_2443_),
    .y(_2444_)
  );
  al_or3fft _6929_ (
    .a(_2442_),
    .b(_2444_),
    .c(_2438_),
    .y(_2445_)
  );
  al_or2ft _6930_ (
    .a(_2439_),
    .b(_2302_),
    .y(_2446_)
  );
  al_nand2 _6931_ (
    .a(_2019_),
    .b(_2021_),
    .y(_2447_)
  );
  al_aoi21ttf _6932_ (
    .a(_2006_),
    .b(_2008_),
    .c(_2441_),
    .y(_2448_)
  );
  al_and3 _6933_ (
    .a(_2443_),
    .b(_2447_),
    .c(_2448_),
    .y(_2449_)
  );
  al_or3ftt _6934_ (
    .a(_2449_),
    .b(_2438_),
    .c(_2446_),
    .y(_2450_)
  );
  al_oai21ftt _6935_ (
    .a(_2302_),
    .b(_2445_),
    .c(_2450_),
    .y(_2451_)
  );
  al_nand2 _6936_ (
    .a(_2431_),
    .b(_2451_),
    .y(_2452_)
  );
  al_and3 _6937_ (
    .a(_2452_),
    .b(_2420_),
    .c(_2429_),
    .y(_2453_)
  );
  al_aoi21 _6938_ (
    .a(_0281_),
    .b(_0284_),
    .c(_2434_),
    .y(_2454_)
  );
  al_nand3 _6939_ (
    .a(_0281_),
    .b(_0284_),
    .c(_2434_),
    .y(_2455_)
  );
  al_nand2ft _6940_ (
    .a(_2454_),
    .b(_2455_),
    .y(_2456_)
  );
  al_ao21ttf _6941_ (
    .a(_2456_),
    .b(_2453_),
    .c(_2430_),
    .y(_2457_)
  );
  al_mux2h _6942_ (
    .a(\DFF_556.Q ),
    .b(_2457_),
    .s(\DFF_1427.Q ),
    .y(\DFF_556.D )
  );
  al_mux2h _6943_ (
    .a(\DFF_557.Q ),
    .b(_2457_),
    .s(\DFF_1428.Q ),
    .y(\DFF_557.D )
  );
  al_mux2h _6944_ (
    .a(\DFF_558.Q ),
    .b(_2457_),
    .s(\DFF_1429.Q ),
    .y(\DFF_558.D )
  );
  al_ao21 _6945_ (
    .a(_2420_),
    .b(_2429_),
    .c(\DFF_654.D ),
    .y(_2458_)
  );
  al_and2ft _6946_ (
    .a(_2439_),
    .b(_2302_),
    .y(_2459_)
  );
  al_nand2ft _6947_ (
    .a(_2459_),
    .b(_2446_),
    .y(_2460_)
  );
  al_mux2l _6948_ (
    .a(_0289_),
    .b(_2302_),
    .s(_2434_),
    .y(_2461_)
  );
  al_nand2 _6949_ (
    .a(_2440_),
    .b(_2302_),
    .y(_2462_)
  );
  al_or2 _6950_ (
    .a(_2440_),
    .b(_2302_),
    .y(_2463_)
  );
  al_aoi21 _6951_ (
    .a(_2462_),
    .b(_2463_),
    .c(_2461_),
    .y(_2464_)
  );
  al_nand2ft _6952_ (
    .a(_2441_),
    .b(_2302_),
    .y(_2465_)
  );
  al_nor2ft _6953_ (
    .a(_2441_),
    .b(_2302_),
    .y(_2466_)
  );
  al_aoi21ftf _6954_ (
    .a(_2466_),
    .b(_2465_),
    .c(_2464_),
    .y(_2467_)
  );
  al_and3ftt _6955_ (
    .a(_2433_),
    .b(_2460_),
    .c(_2467_),
    .y(_2468_)
  );
  al_ao21ttf _6956_ (
    .a(_2460_),
    .b(_2467_),
    .c(_2433_),
    .y(_2469_)
  );
  al_nand2ft _6957_ (
    .a(_2468_),
    .b(_2469_),
    .y(_2470_)
  );
  al_ao21ttf _6958_ (
    .a(_2470_),
    .b(_2453_),
    .c(_2458_),
    .y(_2471_)
  );
  al_mux2h _6959_ (
    .a(\DFF_568.Q ),
    .b(_2471_),
    .s(\DFF_1427.Q ),
    .y(\DFF_568.D )
  );
  al_mux2h _6960_ (
    .a(\DFF_569.Q ),
    .b(_2471_),
    .s(\DFF_1428.Q ),
    .y(\DFF_569.D )
  );
  al_mux2h _6961_ (
    .a(\DFF_570.Q ),
    .b(_2471_),
    .s(\DFF_1429.Q ),
    .y(\DFF_570.D )
  );
  al_ao21 _6962_ (
    .a(_2420_),
    .b(_2429_),
    .c(\DFF_650.D ),
    .y(_2472_)
  );
  al_or2ft _6963_ (
    .a(_2465_),
    .b(_2466_),
    .y(_2473_)
  );
  al_and3 _6964_ (
    .a(_2460_),
    .b(_2464_),
    .c(_2473_),
    .y(_2474_)
  );
  al_and2ft _6965_ (
    .a(_2433_),
    .b(_2302_),
    .y(_2475_)
  );
  al_nor2ft _6966_ (
    .a(_2433_),
    .b(_2302_),
    .y(_2476_)
  );
  al_mux2l _6967_ (
    .a(_2475_),
    .b(_2476_),
    .s(_2432_),
    .y(_2477_)
  );
  al_and3ftt _6968_ (
    .a(_2436_),
    .b(_2477_),
    .c(_2474_),
    .y(_2478_)
  );
  al_ao21ttf _6969_ (
    .a(_2477_),
    .b(_2474_),
    .c(_2436_),
    .y(_2479_)
  );
  al_nand2ft _6970_ (
    .a(_2478_),
    .b(_2479_),
    .y(_2480_)
  );
  al_ao21ttf _6971_ (
    .a(_2480_),
    .b(_2453_),
    .c(_2472_),
    .y(_2481_)
  );
  al_mux2h _6972_ (
    .a(\DFF_574.Q ),
    .b(_2481_),
    .s(\DFF_1427.Q ),
    .y(\DFF_574.D )
  );
  al_mux2h _6973_ (
    .a(\DFF_575.Q ),
    .b(_2481_),
    .s(\DFF_1428.Q ),
    .y(\DFF_575.D )
  );
  al_mux2h _6974_ (
    .a(\DFF_576.Q ),
    .b(_2481_),
    .s(\DFF_1429.Q ),
    .y(\DFF_576.D )
  );
  al_ao21 _6975_ (
    .a(_2420_),
    .b(_2429_),
    .c(\DFF_652.D ),
    .y(_2482_)
  );
  al_or2 _6976_ (
    .a(_2475_),
    .b(_2476_),
    .y(_2483_)
  );
  al_and3 _6977_ (
    .a(_2432_),
    .b(_2483_),
    .c(_2474_),
    .y(_2484_)
  );
  al_ao21 _6978_ (
    .a(_2483_),
    .b(_2474_),
    .c(_2432_),
    .y(_2485_)
  );
  al_nand2ft _6979_ (
    .a(_2484_),
    .b(_2485_),
    .y(_2486_)
  );
  al_ao21ttf _6980_ (
    .a(_2486_),
    .b(_2453_),
    .c(_2482_),
    .y(_2487_)
  );
  al_mux2h _6981_ (
    .a(\DFF_571.Q ),
    .b(_2487_),
    .s(\DFF_1427.Q ),
    .y(\DFF_571.D )
  );
  al_mux2h _6982_ (
    .a(\DFF_572.Q ),
    .b(_2487_),
    .s(\DFF_1428.Q ),
    .y(\DFF_572.D )
  );
  al_mux2h _6983_ (
    .a(\DFF_573.Q ),
    .b(_2487_),
    .s(\DFF_1429.Q ),
    .y(\DFF_573.D )
  );
  al_ao21 _6984_ (
    .a(_2420_),
    .b(_2429_),
    .c(\DFF_648.D ),
    .y(_2488_)
  );
  al_and3 _6985_ (
    .a(_2460_),
    .b(_2477_),
    .c(_2467_),
    .y(_2489_)
  );
  al_and2ft _6986_ (
    .a(_2436_),
    .b(_2302_),
    .y(_2490_)
  );
  al_nor2ft _6987_ (
    .a(_2436_),
    .b(_2302_),
    .y(_2491_)
  );
  al_or2 _6988_ (
    .a(_2490_),
    .b(_2491_),
    .y(_2492_)
  );
  al_and3ftt _6989_ (
    .a(_2435_),
    .b(_2492_),
    .c(_2489_),
    .y(_2493_)
  );
  al_ao21ttf _6990_ (
    .a(_2492_),
    .b(_2489_),
    .c(_2435_),
    .y(_2494_)
  );
  al_nand2ft _6991_ (
    .a(_2493_),
    .b(_2494_),
    .y(_2495_)
  );
  al_ao21ttf _6992_ (
    .a(_2495_),
    .b(_2453_),
    .c(_2488_),
    .y(_2496_)
  );
  al_mux2h _6993_ (
    .a(\DFF_577.Q ),
    .b(_2496_),
    .s(\DFF_1427.Q ),
    .y(\DFF_577.D )
  );
  al_mux2h _6994_ (
    .a(\DFF_578.Q ),
    .b(_2496_),
    .s(\DFF_1428.Q ),
    .y(\DFF_578.D )
  );
  al_mux2h _6995_ (
    .a(\DFF_579.Q ),
    .b(_2496_),
    .s(\DFF_1429.Q ),
    .y(\DFF_579.D )
  );
  al_or3 _6996_ (
    .a(_1102_),
    .b(_0298_),
    .c(_1005_),
    .y(_2497_)
  );
  al_and2ft _6997_ (
    .a(_0304_),
    .b(_0301_),
    .y(_2498_)
  );
  al_nand2ft _6998_ (
    .a(\DFF_993.Q ),
    .b(\DFF_1428.Q ),
    .y(_2499_)
  );
  al_aoi21ftf _6999_ (
    .a(\DFF_994.Q ),
    .b(\DFF_1429.Q ),
    .c(_2499_),
    .y(_2500_)
  );
  al_ao21ftf _7000_ (
    .a(\DFF_992.Q ),
    .b(\DFF_1427.Q ),
    .c(_2500_),
    .y(_2501_)
  );
  al_and3 _7001_ (
    .a(_2501_),
    .b(_2314_),
    .c(_2317_),
    .y(_2502_)
  );
  al_and3 _7002_ (
    .a(_2174_),
    .b(_2498_),
    .c(_2502_),
    .y(_2503_)
  );
  al_nand3 _7003_ (
    .a(_2172_),
    .b(_2162_),
    .c(_2503_),
    .y(_2504_)
  );
  al_aoi21 _7004_ (
    .a(_0308_),
    .b(_2502_),
    .c(_2318_),
    .y(_2505_)
  );
  al_and3 _7005_ (
    .a(_2497_),
    .b(_2505_),
    .c(_2504_),
    .y(_2506_)
  );
  al_and2 _7006_ (
    .a(_2122_),
    .b(_2124_),
    .y(_2507_)
  );
  al_and2 _7007_ (
    .a(_2134_),
    .b(_2136_),
    .y(_2508_)
  );
  al_and2 _7008_ (
    .a(_2085_),
    .b(_2087_),
    .y(_2509_)
  );
  al_nand2 _7009_ (
    .a(_2090_),
    .b(_2092_),
    .y(_2510_)
  );
  al_nand2 _7010_ (
    .a(_2103_),
    .b(_2105_),
    .y(_2511_)
  );
  al_and3fft _7011_ (
    .a(_2510_),
    .b(_2511_),
    .c(_2509_),
    .y(_2512_)
  );
  al_and3 _7012_ (
    .a(_2507_),
    .b(_2508_),
    .c(_2512_),
    .y(_2513_)
  );
  al_nand2 _7013_ (
    .a(_2097_),
    .b(_2099_),
    .y(_2514_)
  );
  al_nand2 _7014_ (
    .a(_2110_),
    .b(_2112_),
    .y(_2515_)
  );
  al_nor3fft _7015_ (
    .a(_0298_),
    .b(_0304_),
    .c(_0306_),
    .y(_2516_)
  );
  al_and3 _7016_ (
    .a(_2514_),
    .b(_2515_),
    .c(_2516_),
    .y(_2517_)
  );
  al_and2 _7017_ (
    .a(_2115_),
    .b(_2117_),
    .y(_2518_)
  );
  al_and2 _7018_ (
    .a(_2127_),
    .b(_2129_),
    .y(_2519_)
  );
  al_and3fft _7019_ (
    .a(_2518_),
    .b(_2519_),
    .c(_2143_),
    .y(_2520_)
  );
  al_nand3 _7020_ (
    .a(_2520_),
    .b(_2517_),
    .c(_2513_),
    .y(_2521_)
  );
  al_nor3fft _7021_ (
    .a(_2097_),
    .b(_2099_),
    .c(_0304_),
    .y(_2522_)
  );
  al_nand3fft _7022_ (
    .a(_2515_),
    .b(_2143_),
    .c(_2522_),
    .y(_2523_)
  );
  al_nor2ft _7023_ (
    .a(_0298_),
    .b(_0306_),
    .y(_2524_)
  );
  al_and3 _7024_ (
    .a(_2518_),
    .b(_2519_),
    .c(_2524_),
    .y(_2525_)
  );
  al_and3ftt _7025_ (
    .a(_2523_),
    .b(_2525_),
    .c(_2513_),
    .y(_2526_)
  );
  al_and2ft _7026_ (
    .a(_2526_),
    .b(_2521_),
    .y(_2527_)
  );
  al_ao21ttf _7027_ (
    .a(_0298_),
    .b(_0301_),
    .c(_2511_),
    .y(_2528_)
  );
  al_nor3ftt _7028_ (
    .a(_0298_),
    .b(_0306_),
    .c(_2511_),
    .y(_2529_)
  );
  al_nand2ft _7029_ (
    .a(_2529_),
    .b(_2528_),
    .y(_2530_)
  );
  al_nand3 _7030_ (
    .a(_2527_),
    .b(_2530_),
    .c(_2506_),
    .y(_2531_)
  );
  al_ao21ftf _7031_ (
    .a(_2506_),
    .b(\DFF_45.Q ),
    .c(_2531_),
    .y(_2532_)
  );
  al_mux2h _7032_ (
    .a(\DFF_906.Q ),
    .b(_2532_),
    .s(\DFF_1427.Q ),
    .y(\DFF_906.D )
  );
  al_mux2h _7033_ (
    .a(\DFF_907.Q ),
    .b(_2532_),
    .s(\DFF_1428.Q ),
    .y(\DFF_907.D )
  );
  al_mux2h _7034_ (
    .a(\DFF_908.Q ),
    .b(_2532_),
    .s(\DFF_1429.Q ),
    .y(\DFF_908.D )
  );
  al_and3 _7035_ (
    .a(_0304_),
    .b(_2514_),
    .c(_2524_),
    .y(_2533_)
  );
  al_nand2ft _7036_ (
    .a(_2514_),
    .b(_2308_),
    .y(_2534_)
  );
  al_mux2h _7037_ (
    .a(_2511_),
    .b(_2529_),
    .s(_2308_),
    .y(_2535_)
  );
  al_oa21ftt _7038_ (
    .a(_2534_),
    .b(_2533_),
    .c(_2535_),
    .y(_2536_)
  );
  al_and2 _7039_ (
    .a(_2518_),
    .b(_2308_),
    .y(_2537_)
  );
  al_and3ftt _7040_ (
    .a(_2518_),
    .b(_0304_),
    .c(_2524_),
    .y(_2538_)
  );
  al_mux2h _7041_ (
    .a(_2538_),
    .b(_2537_),
    .s(_2519_),
    .y(_2539_)
  );
  al_ao21 _7042_ (
    .a(_2539_),
    .b(_2536_),
    .c(_2509_),
    .y(_2540_)
  );
  al_and3 _7043_ (
    .a(_2509_),
    .b(_2539_),
    .c(_2536_),
    .y(_2541_)
  );
  al_nand2ft _7044_ (
    .a(_2541_),
    .b(_2540_),
    .y(_2542_)
  );
  al_nand3 _7045_ (
    .a(_2527_),
    .b(_2542_),
    .c(_2506_),
    .y(_2543_)
  );
  al_ao21ftf _7046_ (
    .a(_2506_),
    .b(\DFF_41.Q ),
    .c(_2543_),
    .y(_2544_)
  );
  al_mux2h _7047_ (
    .a(\DFF_918.Q ),
    .b(_2544_),
    .s(\DFF_1427.Q ),
    .y(\DFF_918.D )
  );
  al_mux2h _7048_ (
    .a(\DFF_919.Q ),
    .b(_2544_),
    .s(\DFF_1428.Q ),
    .y(\DFF_919.D )
  );
  al_mux2h _7049_ (
    .a(\DFF_920.Q ),
    .b(_2544_),
    .s(\DFF_1429.Q ),
    .y(\DFF_920.D )
  );
  al_nand2ft _7050_ (
    .a(_2533_),
    .b(_2534_),
    .y(_2545_)
  );
  al_and3 _7051_ (
    .a(_2535_),
    .b(_2545_),
    .c(_2539_),
    .y(_2546_)
  );
  al_nand3 _7052_ (
    .a(_2509_),
    .b(_2507_),
    .c(_2308_),
    .y(_2547_)
  );
  al_and3ftt _7053_ (
    .a(_2509_),
    .b(_0304_),
    .c(_2524_),
    .y(_2548_)
  );
  al_ao21ftf _7054_ (
    .a(_2507_),
    .b(_2548_),
    .c(_2547_),
    .y(_2549_)
  );
  al_and3ftt _7055_ (
    .a(_2510_),
    .b(_2549_),
    .c(_2546_),
    .y(_2550_)
  );
  al_and3 _7056_ (
    .a(_2549_),
    .b(_2536_),
    .c(_2539_),
    .y(_2551_)
  );
  al_or2ft _7057_ (
    .a(_2510_),
    .b(_2551_),
    .y(_2552_)
  );
  al_nand2ft _7058_ (
    .a(_2550_),
    .b(_2552_),
    .y(_2553_)
  );
  al_nand3 _7059_ (
    .a(_2527_),
    .b(_2553_),
    .c(_2506_),
    .y(_2554_)
  );
  al_ao21ftf _7060_ (
    .a(_2506_),
    .b(\DFF_39.Q ),
    .c(_2554_),
    .y(_2555_)
  );
  al_mux2h _7061_ (
    .a(\DFF_924.Q ),
    .b(_2555_),
    .s(\DFF_1427.Q ),
    .y(\DFF_924.D )
  );
  al_mux2h _7062_ (
    .a(\DFF_925.Q ),
    .b(_2555_),
    .s(\DFF_1428.Q ),
    .y(\DFF_925.D )
  );
  al_mux2h _7063_ (
    .a(\DFF_926.Q ),
    .b(_2555_),
    .s(\DFF_1429.Q ),
    .y(\DFF_926.D )
  );
  al_nand2 _7064_ (
    .a(_2509_),
    .b(_2308_),
    .y(_2556_)
  );
  al_ao21ftf _7065_ (
    .a(_2548_),
    .b(_2556_),
    .c(_2546_),
    .y(_2557_)
  );
  al_and2ft _7066_ (
    .a(_2507_),
    .b(_2557_),
    .y(_2558_)
  );
  al_or3fft _7067_ (
    .a(_2122_),
    .b(_2124_),
    .c(_2557_),
    .y(_2559_)
  );
  al_nand2ft _7068_ (
    .a(_2558_),
    .b(_2559_),
    .y(_2560_)
  );
  al_nand3 _7069_ (
    .a(_2527_),
    .b(_2560_),
    .c(_2506_),
    .y(_2561_)
  );
  al_ao21ftf _7070_ (
    .a(_2506_),
    .b(\DFF_40.Q ),
    .c(_2561_),
    .y(_2562_)
  );
  al_mux2h _7071_ (
    .a(\DFF_921.Q ),
    .b(_2562_),
    .s(\DFF_1427.Q ),
    .y(\DFF_921.D )
  );
  al_mux2h _7072_ (
    .a(\DFF_922.Q ),
    .b(_2562_),
    .s(\DFF_1428.Q ),
    .y(\DFF_922.D )
  );
  al_mux2h _7073_ (
    .a(\DFF_923.Q ),
    .b(_2562_),
    .s(\DFF_1429.Q ),
    .y(\DFF_923.D )
  );
  al_nand2ft _7074_ (
    .a(_2510_),
    .b(_2308_),
    .y(_2563_)
  );
  al_and3 _7075_ (
    .a(_0304_),
    .b(_2510_),
    .c(_2524_),
    .y(_2564_)
  );
  al_ao21ftf _7076_ (
    .a(_2564_),
    .b(_2563_),
    .c(_2551_),
    .y(_2565_)
  );
  al_or2ft _7077_ (
    .a(_2508_),
    .b(_2565_),
    .y(_2566_)
  );
  al_and2ft _7078_ (
    .a(_2508_),
    .b(_2565_),
    .y(_2567_)
  );
  al_nand2ft _7079_ (
    .a(_2567_),
    .b(_2566_),
    .y(_2568_)
  );
  al_nand3 _7080_ (
    .a(_2527_),
    .b(_2568_),
    .c(_2506_),
    .y(_2569_)
  );
  al_ao21ftf _7081_ (
    .a(_2506_),
    .b(\DFF_38.Q ),
    .c(_2569_),
    .y(_2570_)
  );
  al_mux2h _7082_ (
    .a(\DFF_927.Q ),
    .b(_2570_),
    .s(\DFF_1427.Q ),
    .y(\DFF_927.D )
  );
  al_mux2h _7083_ (
    .a(\DFF_928.Q ),
    .b(_2570_),
    .s(\DFF_1428.Q ),
    .y(\DFF_928.D )
  );
  al_mux2h _7084_ (
    .a(\DFF_929.Q ),
    .b(_2570_),
    .s(\DFF_1429.Q ),
    .y(\DFF_929.D )
  );
  al_or3fft _7085_ (
    .a(\DFF_1302.Q ),
    .b(_0314_),
    .c(_1084_),
    .y(_2571_)
  );
  al_nand2ft _7086_ (
    .a(\DFF_1343.Q ),
    .b(\DFF_1428.Q ),
    .y(_2572_)
  );
  al_aoi21ftf _7087_ (
    .a(\DFF_1344.Q ),
    .b(\DFF_1429.Q ),
    .c(_2572_),
    .y(_2573_)
  );
  al_ao21ftf _7088_ (
    .a(\DFF_1342.Q ),
    .b(\DFF_1427.Q ),
    .c(_2573_),
    .y(_2574_)
  );
  al_nand3 _7089_ (
    .a(_0323_),
    .b(_2574_),
    .c(_1088_),
    .y(_2575_)
  );
  al_nor3fft _7090_ (
    .a(_2571_),
    .b(_2575_),
    .c(_2324_),
    .y(_2576_)
  );
  al_and2ft _7091_ (
    .a(_0320_),
    .b(_0317_),
    .y(_2577_)
  );
  al_nor2ft _7092_ (
    .a(_1081_),
    .b(_1080_),
    .y(_2578_)
  );
  al_and3fft _7093_ (
    .a(_2256_),
    .b(_1023_),
    .c(_1022_),
    .y(_2579_)
  );
  al_and3 _7094_ (
    .a(_2579_),
    .b(_2578_),
    .c(_1056_),
    .y(_2580_)
  );
  al_aoi21ftf _7095_ (
    .a(_1049_),
    .b(_1048_),
    .c(_1070_),
    .y(_2581_)
  );
  al_and3 _7096_ (
    .a(_1063_),
    .b(_1037_),
    .c(_1043_),
    .y(_2582_)
  );
  al_and3 _7097_ (
    .a(_1076_),
    .b(_2581_),
    .c(_2582_),
    .y(_2583_)
  );
  al_and3 _7098_ (
    .a(_2580_),
    .b(_2574_),
    .c(_2583_),
    .y(_2584_)
  );
  al_and3 _7099_ (
    .a(_0314_),
    .b(_2577_),
    .c(_2584_),
    .y(_2585_)
  );
  al_nand3 _7100_ (
    .a(_2275_),
    .b(_2266_),
    .c(_2585_),
    .y(_2586_)
  );
  al_ao21 _7101_ (
    .a(_2576_),
    .b(_2586_),
    .c(\DFF_1362.D ),
    .y(_2587_)
  );
  al_and2 _7102_ (
    .a(_2193_),
    .b(_2195_),
    .y(_2588_)
  );
  al_and2 _7103_ (
    .a(_2239_),
    .b(_2241_),
    .y(_2589_)
  );
  al_and3ftt _7104_ (
    .a(_2217_),
    .b(_2588_),
    .c(_2589_),
    .y(_2590_)
  );
  al_nand3 _7105_ (
    .a(_2211_),
    .b(_2235_),
    .c(_2590_),
    .y(_2591_)
  );
  al_nand2 _7106_ (
    .a(_2220_),
    .b(_2222_),
    .y(_2592_)
  );
  al_nand2 _7107_ (
    .a(_2227_),
    .b(_2229_),
    .y(_2593_)
  );
  al_nand2 _7108_ (
    .a(_2245_),
    .b(_2247_),
    .y(_2594_)
  );
  al_or3 _7109_ (
    .a(_2592_),
    .b(_2593_),
    .c(_2594_),
    .y(_2595_)
  );
  al_and2ft _7110_ (
    .a(_2190_),
    .b(_2204_),
    .y(_2596_)
  );
  al_and3fft _7111_ (
    .a(_2595_),
    .b(_2591_),
    .c(_2596_),
    .y(_2597_)
  );
  al_nand3 _7112_ (
    .a(_0320_),
    .b(_2593_),
    .c(_1387_),
    .y(_2598_)
  );
  al_aoi21ttf _7113_ (
    .a(_2245_),
    .b(_2247_),
    .c(_2592_),
    .y(_2599_)
  );
  al_nand3 _7114_ (
    .a(_2190_),
    .b(_2202_),
    .c(_2599_),
    .y(_2600_)
  );
  al_or3 _7115_ (
    .a(_2598_),
    .b(_2600_),
    .c(_2591_),
    .y(_2601_)
  );
  al_ao21ttf _7116_ (
    .a(_2321_),
    .b(_2597_),
    .c(_2601_),
    .y(_2602_)
  );
  al_nand2 _7117_ (
    .a(_1387_),
    .b(_2602_),
    .y(_2603_)
  );
  al_and3 _7118_ (
    .a(_2603_),
    .b(_2576_),
    .c(_2586_),
    .y(_2604_)
  );
  al_ao21ftf _7119_ (
    .a(_0314_),
    .b(_0317_),
    .c(_2209_),
    .y(_2605_)
  );
  al_and3fft _7120_ (
    .a(_0314_),
    .b(_2209_),
    .c(_0317_),
    .y(_2606_)
  );
  al_nand2ft _7121_ (
    .a(_2606_),
    .b(_2605_),
    .y(_2607_)
  );
  al_ao21ttf _7122_ (
    .a(_2607_),
    .b(_2604_),
    .c(_2587_),
    .y(_2608_)
  );
  al_mux2h _7123_ (
    .a(\DFF_1256.Q ),
    .b(_2608_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1256.D )
  );
  al_mux2h _7124_ (
    .a(\DFF_1257.Q ),
    .b(_2608_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1257.D )
  );
  al_mux2h _7125_ (
    .a(\DFF_1258.Q ),
    .b(_2608_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1258.D )
  );
  al_ao21 _7126_ (
    .a(_2576_),
    .b(_2586_),
    .c(\DFF_1354.D ),
    .y(_2609_)
  );
  al_and2ft _7127_ (
    .a(_2593_),
    .b(_2321_),
    .y(_2610_)
  );
  al_or2ft _7128_ (
    .a(_2598_),
    .b(_2610_),
    .y(_2611_)
  );
  al_mux2h _7129_ (
    .a(_2209_),
    .b(_2606_),
    .s(_2321_),
    .y(_2612_)
  );
  al_nand2 _7130_ (
    .a(_2204_),
    .b(_2321_),
    .y(_2613_)
  );
  al_nand3 _7131_ (
    .a(_0320_),
    .b(_2202_),
    .c(_1387_),
    .y(_2614_)
  );
  al_aoi21ttf _7132_ (
    .a(_2614_),
    .b(_2613_),
    .c(_2612_),
    .y(_2615_)
  );
  al_nand2ft _7133_ (
    .a(_2592_),
    .b(_2321_),
    .y(_2616_)
  );
  al_and3 _7134_ (
    .a(_0320_),
    .b(_2592_),
    .c(_1387_),
    .y(_2617_)
  );
  al_aoi21ftf _7135_ (
    .a(_2617_),
    .b(_2616_),
    .c(_2615_),
    .y(_2618_)
  );
  al_ao21ttf _7136_ (
    .a(_2611_),
    .b(_2618_),
    .c(_2217_),
    .y(_2619_)
  );
  al_and3ftt _7137_ (
    .a(_2217_),
    .b(_2611_),
    .c(_2618_),
    .y(_2620_)
  );
  al_nand2ft _7138_ (
    .a(_2620_),
    .b(_2619_),
    .y(_2621_)
  );
  al_ao21ttf _7139_ (
    .a(_2621_),
    .b(_2604_),
    .c(_2609_),
    .y(_2622_)
  );
  al_mux2h _7140_ (
    .a(\DFF_1268.Q ),
    .b(_2622_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1268.D )
  );
  al_mux2h _7141_ (
    .a(\DFF_1269.Q ),
    .b(_2622_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1269.D )
  );
  al_mux2h _7142_ (
    .a(\DFF_1270.Q ),
    .b(_2622_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1270.D )
  );
  al_ao21 _7143_ (
    .a(_2576_),
    .b(_2586_),
    .c(\DFF_1350.D ),
    .y(_2623_)
  );
  al_nand2ft _7144_ (
    .a(_2617_),
    .b(_2616_),
    .y(_2624_)
  );
  al_and3 _7145_ (
    .a(_2624_),
    .b(_2611_),
    .c(_2615_),
    .y(_2625_)
  );
  al_and2ft _7146_ (
    .a(_2217_),
    .b(_2321_),
    .y(_2626_)
  );
  al_and3 _7147_ (
    .a(_0320_),
    .b(_2217_),
    .c(_1387_),
    .y(_2627_)
  );
  al_mux2h _7148_ (
    .a(_2627_),
    .b(_2626_),
    .s(_2235_),
    .y(_2628_)
  );
  al_ao21 _7149_ (
    .a(_2628_),
    .b(_2625_),
    .c(_2588_),
    .y(_2629_)
  );
  al_and3 _7150_ (
    .a(_2588_),
    .b(_2628_),
    .c(_2625_),
    .y(_2630_)
  );
  al_nand2ft _7151_ (
    .a(_2630_),
    .b(_2629_),
    .y(_2631_)
  );
  al_ao21ttf _7152_ (
    .a(_2631_),
    .b(_2604_),
    .c(_2623_),
    .y(_2632_)
  );
  al_mux2h _7153_ (
    .a(\DFF_1274.Q ),
    .b(_2632_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1274.D )
  );
  al_mux2h _7154_ (
    .a(\DFF_1275.Q ),
    .b(_2632_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1275.D )
  );
  al_mux2h _7155_ (
    .a(\DFF_1276.Q ),
    .b(_2632_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1276.D )
  );
  al_ao21 _7156_ (
    .a(_2576_),
    .b(_2586_),
    .c(\DFF_1352.D ),
    .y(_2633_)
  );
  al_or2 _7157_ (
    .a(_2627_),
    .b(_2626_),
    .y(_2634_)
  );
  al_ao21 _7158_ (
    .a(_2634_),
    .b(_2625_),
    .c(_2235_),
    .y(_2635_)
  );
  al_and3 _7159_ (
    .a(_2235_),
    .b(_2634_),
    .c(_2625_),
    .y(_2636_)
  );
  al_nand2ft _7160_ (
    .a(_2636_),
    .b(_2635_),
    .y(_2637_)
  );
  al_ao21ttf _7161_ (
    .a(_2637_),
    .b(_2604_),
    .c(_2633_),
    .y(_2638_)
  );
  al_mux2h _7162_ (
    .a(\DFF_1271.Q ),
    .b(_2638_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1271.D )
  );
  al_mux2h _7163_ (
    .a(\DFF_1272.Q ),
    .b(_2638_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1272.D )
  );
  al_mux2h _7164_ (
    .a(\DFF_1273.Q ),
    .b(_2638_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1273.D )
  );
  al_ao21 _7165_ (
    .a(_2576_),
    .b(_2586_),
    .c(\DFF_1348.D ),
    .y(_2639_)
  );
  al_and3 _7166_ (
    .a(_2611_),
    .b(_2628_),
    .c(_2618_),
    .y(_2640_)
  );
  al_nand2 _7167_ (
    .a(_2588_),
    .b(_2321_),
    .y(_2641_)
  );
  al_and3ftt _7168_ (
    .a(_2588_),
    .b(_0320_),
    .c(_1387_),
    .y(_2642_)
  );
  al_nand2ft _7169_ (
    .a(_2642_),
    .b(_2641_),
    .y(_2643_)
  );
  al_and3 _7170_ (
    .a(_2589_),
    .b(_2643_),
    .c(_2640_),
    .y(_2644_)
  );
  al_ao21 _7171_ (
    .a(_2643_),
    .b(_2640_),
    .c(_2589_),
    .y(_2645_)
  );
  al_nand2ft _7172_ (
    .a(_2644_),
    .b(_2645_),
    .y(_2646_)
  );
  al_ao21ttf _7173_ (
    .a(_2646_),
    .b(_2604_),
    .c(_2639_),
    .y(_2647_)
  );
  al_mux2h _7174_ (
    .a(\DFF_1277.Q ),
    .b(_2647_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1277.D )
  );
  al_mux2h _7175_ (
    .a(\DFF_1278.Q ),
    .b(_2647_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1278.D )
  );
  al_mux2h _7176_ (
    .a(\DFF_1279.Q ),
    .b(_2647_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1279.D )
  );
  al_nand3 _7177_ (
    .a(\DFF_1302.Q ),
    .b(_2350_),
    .c(_1966_),
    .y(_2648_)
  );
  al_nand2ft _7178_ (
    .a(_0848_),
    .b(_1942_),
    .y(_2649_)
  );
  al_ao21 _7179_ (
    .a(_0847_),
    .b(_1942_),
    .c(_1102_),
    .y(_2650_)
  );
  al_aoi21 _7180_ (
    .a(_0270_),
    .b(_2650_),
    .c(_1945_),
    .y(_2651_)
  );
  al_ao21ftf _7181_ (
    .a(_0270_),
    .b(_2649_),
    .c(_2651_),
    .y(_2652_)
  );
  al_ao21ttf _7182_ (
    .a(_2648_),
    .b(_2652_),
    .c(_0270_),
    .y(_2653_)
  );
  al_aoi21ttf _7183_ (
    .a(_0783_),
    .b(_0851_),
    .c(_0267_),
    .y(_2654_)
  );
  al_nand3ftt _7184_ (
    .a(_0270_),
    .b(_2648_),
    .c(_2652_),
    .y(_2655_)
  );
  al_and3 _7185_ (
    .a(_2654_),
    .b(_2655_),
    .c(_2653_),
    .y(_2656_)
  );
  al_mux2h _7186_ (
    .a(\DFF_289.Q ),
    .b(_2656_),
    .s(\DFF_1427.Q ),
    .y(\DFF_289.D )
  );
  al_mux2h _7187_ (
    .a(\DFF_290.Q ),
    .b(_2656_),
    .s(\DFF_1428.Q ),
    .y(\DFF_290.D )
  );
  al_mux2h _7188_ (
    .a(\DFF_291.Q ),
    .b(_2656_),
    .s(\DFF_1429.Q ),
    .y(\DFF_291.D )
  );
  al_ao21 _7189_ (
    .a(\DFF_1302.Q ),
    .b(_2062_),
    .c(_0287_),
    .y(_2657_)
  );
  al_aoi21 _7190_ (
    .a(_2037_),
    .b(_2012_),
    .c(_2050_),
    .y(_2658_)
  );
  al_ao21ftf _7191_ (
    .a(_0284_),
    .b(_2658_),
    .c(_0287_),
    .y(_2659_)
  );
  al_ao21 _7192_ (
    .a(_2659_),
    .b(_2657_),
    .c(_0284_),
    .y(_2660_)
  );
  al_or3fft _7193_ (
    .a(_2005_),
    .b(_2041_),
    .c(_1999_),
    .y(_2661_)
  );
  al_nand3fft _7194_ (
    .a(_1987_),
    .b(_2661_),
    .c(_2037_),
    .y(_2662_)
  );
  al_ao21ftf _7195_ (
    .a(_0926_),
    .b(_2662_),
    .c(\DFF_1302.Q ),
    .y(_2663_)
  );
  al_aoi21ttf _7196_ (
    .a(_0287_),
    .b(_2663_),
    .c(_0284_),
    .y(_2664_)
  );
  al_ao21 _7197_ (
    .a(_0863_),
    .b(_2074_),
    .c(_0281_),
    .y(_2665_)
  );
  al_aoi21 _7198_ (
    .a(_2664_),
    .b(_2657_),
    .c(_2665_),
    .y(_2666_)
  );
  al_nand3 _7199_ (
    .a(\DFF_1427.Q ),
    .b(_2660_),
    .c(_2666_),
    .y(_2667_)
  );
  al_ao21ftf _7200_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_639.Q ),
    .c(_2667_),
    .y(\DFF_639.D )
  );
  al_nand3 _7201_ (
    .a(\DFF_1428.Q ),
    .b(_2660_),
    .c(_2666_),
    .y(_2668_)
  );
  al_ao21ftf _7202_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_640.Q ),
    .c(_2668_),
    .y(\DFF_640.D )
  );
  al_nand3 _7203_ (
    .a(\DFF_1429.Q ),
    .b(_2660_),
    .c(_2666_),
    .y(_2669_)
  );
  al_ao21ftf _7204_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_641.Q ),
    .c(_2669_),
    .y(\DFF_641.D )
  );
  al_ao21 _7205_ (
    .a(\DFF_1302.Q ),
    .b(_2173_),
    .c(_0304_),
    .y(_2670_)
  );
  al_aoi21 _7206_ (
    .a(_2109_),
    .b(_2147_),
    .c(_1006_),
    .y(_2671_)
  );
  al_ao21ttf _7207_ (
    .a(_0306_),
    .b(_2671_),
    .c(_0304_),
    .y(_2672_)
  );
  al_ao21 _7208_ (
    .a(_2672_),
    .b(_2670_),
    .c(_0301_),
    .y(_2673_)
  );
  al_nand3fft _7209_ (
    .a(_1102_),
    .b(_0306_),
    .c(_2148_),
    .y(_2674_)
  );
  al_nand2ft _7210_ (
    .a(_2498_),
    .b(_2674_),
    .y(_2675_)
  );
  al_aoi21ftf _7211_ (
    .a(_1000_),
    .b(\DFF_43.Q ),
    .c(_0951_),
    .y(_2676_)
  );
  al_and3 _7212_ (
    .a(_0973_),
    .b(_2676_),
    .c(_0991_),
    .y(_2677_)
  );
  al_aoi21ftf _7213_ (
    .a(_0944_),
    .b(\DFF_998.D ),
    .c(_0958_),
    .y(_2678_)
  );
  al_and3ftt _7214_ (
    .a(_0946_),
    .b(_0959_),
    .c(_2678_),
    .y(_2679_)
  );
  al_aoi21ftf _7215_ (
    .a(_0976_),
    .b(_0218_),
    .c(_1002_),
    .y(_2680_)
  );
  al_aoi21ftf _7216_ (
    .a(_0950_),
    .b(\DFF_42.Q ),
    .c(_0978_),
    .y(_2681_)
  );
  al_nand3 _7217_ (
    .a(_2680_),
    .b(_2681_),
    .c(_2679_),
    .y(_2682_)
  );
  al_nand2 _7218_ (
    .a(_0979_),
    .b(_0981_),
    .y(_2683_)
  );
  al_aoi21ftt _7219_ (
    .a(\DFF_39.Q ),
    .b(_2683_),
    .c(_1006_),
    .y(_2684_)
  );
  al_aoi21ftf _7220_ (
    .a(_2683_),
    .b(\DFF_39.Q ),
    .c(_2684_),
    .y(_2685_)
  );
  al_nand3 _7221_ (
    .a(_0965_),
    .b(_0997_),
    .c(_2685_),
    .y(_2686_)
  );
  al_nor3ftt _7222_ (
    .a(_2677_),
    .b(_2682_),
    .c(_2686_),
    .y(_2687_)
  );
  al_ao21 _7223_ (
    .a(_0941_),
    .b(_2687_),
    .c(_0298_),
    .y(_2688_)
  );
  al_aoi21 _7224_ (
    .a(_2675_),
    .b(_2670_),
    .c(_2688_),
    .y(_2689_)
  );
  al_nand3 _7225_ (
    .a(\DFF_1427.Q ),
    .b(_2673_),
    .c(_2689_),
    .y(_2690_)
  );
  al_ao21ftf _7226_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_989.Q ),
    .c(_2690_),
    .y(\DFF_989.D )
  );
  al_nand3 _7227_ (
    .a(\DFF_1428.Q ),
    .b(_2673_),
    .c(_2689_),
    .y(_2691_)
  );
  al_ao21ftf _7228_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_990.Q ),
    .c(_2691_),
    .y(\DFF_990.D )
  );
  al_nand3 _7229_ (
    .a(\DFF_1429.Q ),
    .b(_2673_),
    .c(_2689_),
    .y(_2692_)
  );
  al_ao21ftf _7230_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_991.Q ),
    .c(_2692_),
    .y(\DFF_991.D )
  );
  al_ao21 _7231_ (
    .a(\DFF_1302.Q ),
    .b(_2276_),
    .c(_0320_),
    .y(_2693_)
  );
  al_inv _7232_ (
    .a(_0320_),
    .y(_2694_)
  );
  al_ao21 _7233_ (
    .a(_1085_),
    .b(_2252_),
    .c(_2694_),
    .y(_2695_)
  );
  al_ao21 _7234_ (
    .a(_2695_),
    .b(_2693_),
    .c(_0317_),
    .y(_2696_)
  );
  al_inv _7235_ (
    .a(_0317_),
    .y(_2697_)
  );
  al_ao21 _7236_ (
    .a(_1084_),
    .b(_2252_),
    .c(_1102_),
    .y(_2698_)
  );
  al_aoi21 _7237_ (
    .a(_0320_),
    .b(_2698_),
    .c(_2697_),
    .y(_2699_)
  );
  al_ao21ttf _7238_ (
    .a(_1018_),
    .b(_1088_),
    .c(_0314_),
    .y(_2700_)
  );
  al_aoi21 _7239_ (
    .a(_2699_),
    .b(_2693_),
    .c(_2700_),
    .y(_2701_)
  );
  al_nand3 _7240_ (
    .a(\DFF_1427.Q ),
    .b(_2696_),
    .c(_2701_),
    .y(_2702_)
  );
  al_ao21ftf _7241_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_1339.Q ),
    .c(_2702_),
    .y(\DFF_1339.D )
  );
  al_nand3 _7242_ (
    .a(\DFF_1428.Q ),
    .b(_2696_),
    .c(_2701_),
    .y(_2703_)
  );
  al_ao21ftf _7243_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_1340.Q ),
    .c(_2703_),
    .y(\DFF_1340.D )
  );
  al_nand3 _7244_ (
    .a(\DFF_1429.Q ),
    .b(_2696_),
    .c(_2701_),
    .y(_2704_)
  );
  al_ao21ftf _7245_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_1341.Q ),
    .c(_2704_),
    .y(\DFF_1341.D )
  );
  al_and3 _7246_ (
    .a(_2350_),
    .b(_2296_),
    .c(_1965_),
    .y(_2705_)
  );
  al_ao21ttf _7247_ (
    .a(_2351_),
    .b(_2705_),
    .c(_2349_),
    .y(_2706_)
  );
  al_nand3 _7248_ (
    .a(_2365_),
    .b(_2367_),
    .c(_2357_),
    .y(_2707_)
  );
  al_mux2l _7249_ (
    .a(\DFF_76.Q ),
    .b(_2707_),
    .s(_2706_),
    .y(_2708_)
  );
  al_aoi21ttf _7250_ (
    .a(_2351_),
    .b(_2705_),
    .c(_2349_),
    .y(_2709_)
  );
  al_or3fft _7251_ (
    .a(_1904_),
    .b(_1906_),
    .c(_2382_),
    .y(_2710_)
  );
  al_and2 _7252_ (
    .a(_2359_),
    .b(_2382_),
    .y(_2711_)
  );
  al_nand2ft _7253_ (
    .a(_2711_),
    .b(_2710_),
    .y(_2712_)
  );
  al_nand3 _7254_ (
    .a(_2369_),
    .b(_2712_),
    .c(_2709_),
    .y(_2713_)
  );
  al_nand3 _7255_ (
    .a(\DFF_1427.Q ),
    .b(_2713_),
    .c(_2708_),
    .y(_2714_)
  );
  al_ao21ftf _7256_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_212.Q ),
    .c(_2714_),
    .y(\DFF_212.D )
  );
  al_nand3 _7257_ (
    .a(\DFF_1428.Q ),
    .b(_2713_),
    .c(_2708_),
    .y(_2715_)
  );
  al_ao21ftf _7258_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_213.Q ),
    .c(_2715_),
    .y(\DFF_213.D )
  );
  al_nand3 _7259_ (
    .a(\DFF_1429.Q ),
    .b(_2713_),
    .c(_2708_),
    .y(_2716_)
  );
  al_ao21ftf _7260_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_214.Q ),
    .c(_2716_),
    .y(\DFF_214.D )
  );
  al_mux2l _7261_ (
    .a(_0161_),
    .b(_2707_),
    .s(_2706_),
    .y(_2717_)
  );
  al_nand3ftt _7262_ (
    .a(_1900_),
    .b(_2355_),
    .c(_2295_),
    .y(_2718_)
  );
  al_ao21ftf _7263_ (
    .a(_2355_),
    .b(_2409_),
    .c(_2718_),
    .y(_2719_)
  );
  al_ao21 _7264_ (
    .a(_2719_),
    .b(_2407_),
    .c(_1912_),
    .y(_2720_)
  );
  al_and3 _7265_ (
    .a(_1912_),
    .b(_2719_),
    .c(_2407_),
    .y(_2721_)
  );
  al_nand2ft _7266_ (
    .a(_2721_),
    .b(_2720_),
    .y(_2722_)
  );
  al_nand3 _7267_ (
    .a(_2369_),
    .b(_2722_),
    .c(_2709_),
    .y(_2723_)
  );
  al_nand3 _7268_ (
    .a(\DFF_1427.Q ),
    .b(_2723_),
    .c(_2717_),
    .y(_2724_)
  );
  al_ao21ftf _7269_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_230.Q ),
    .c(_2724_),
    .y(\DFF_230.D )
  );
  al_nand3 _7270_ (
    .a(\DFF_1428.Q ),
    .b(_2723_),
    .c(_2717_),
    .y(_2725_)
  );
  al_ao21ftf _7271_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_231.Q ),
    .c(_2725_),
    .y(\DFF_231.D )
  );
  al_nand3 _7272_ (
    .a(\DFF_1429.Q ),
    .b(_2723_),
    .c(_2717_),
    .y(_2726_)
  );
  al_ao21ftf _7273_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_232.Q ),
    .c(_2726_),
    .y(\DFF_232.D )
  );
  al_mux2l _7274_ (
    .a(\DFF_78.Q ),
    .b(_2707_),
    .s(_2706_),
    .y(_2727_)
  );
  al_or3fft _7275_ (
    .a(_1934_),
    .b(_1936_),
    .c(_2379_),
    .y(_2728_)
  );
  al_inv _7276_ (
    .a(_2361_),
    .y(_2729_)
  );
  al_and2 _7277_ (
    .a(_2729_),
    .b(_2379_),
    .y(_2730_)
  );
  al_nand2ft _7278_ (
    .a(_2730_),
    .b(_2728_),
    .y(_2731_)
  );
  al_nand3 _7279_ (
    .a(_2369_),
    .b(_2731_),
    .c(_2709_),
    .y(_2732_)
  );
  al_nand3 _7280_ (
    .a(\DFF_1427.Q ),
    .b(_2732_),
    .c(_2727_),
    .y(_2733_)
  );
  al_ao21ftf _7281_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_209.Q ),
    .c(_2733_),
    .y(\DFF_209.D )
  );
  al_nand3 _7282_ (
    .a(\DFF_1428.Q ),
    .b(_2732_),
    .c(_2727_),
    .y(_2734_)
  );
  al_ao21ftf _7283_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_210.Q ),
    .c(_2734_),
    .y(\DFF_210.D )
  );
  al_nand3 _7284_ (
    .a(\DFF_1429.Q ),
    .b(_2732_),
    .c(_2727_),
    .y(_2735_)
  );
  al_ao21ftf _7285_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_211.Q ),
    .c(_2735_),
    .y(\DFF_211.D )
  );
  al_mux2l _7286_ (
    .a(\DFF_74.Q ),
    .b(_2707_),
    .s(_2706_),
    .y(_2736_)
  );
  al_ao21 _7287_ (
    .a(_2391_),
    .b(_2382_),
    .c(_2360_),
    .y(_2737_)
  );
  al_and3 _7288_ (
    .a(_2360_),
    .b(_2391_),
    .c(_2382_),
    .y(_2738_)
  );
  al_nand2ft _7289_ (
    .a(_2738_),
    .b(_2737_),
    .y(_2739_)
  );
  al_nand3 _7290_ (
    .a(_2369_),
    .b(_2739_),
    .c(_2709_),
    .y(_2740_)
  );
  al_nand3 _7291_ (
    .a(\DFF_1427.Q ),
    .b(_2740_),
    .c(_2736_),
    .y(_2741_)
  );
  al_ao21ftf _7292_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_215.Q ),
    .c(_2741_),
    .y(\DFF_215.D )
  );
  al_nand3 _7293_ (
    .a(\DFF_1428.Q ),
    .b(_2740_),
    .c(_2736_),
    .y(_2742_)
  );
  al_ao21ftf _7294_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_216.Q ),
    .c(_2742_),
    .y(\DFF_216.D )
  );
  al_nand3 _7295_ (
    .a(\DFF_1429.Q ),
    .b(_2740_),
    .c(_2736_),
    .y(_2743_)
  );
  al_ao21ftf _7296_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_217.Q ),
    .c(_2743_),
    .y(\DFF_217.D )
  );
  al_mux2l _7297_ (
    .a(_0165_),
    .b(_2707_),
    .s(_2706_),
    .y(_2744_)
  );
  al_and3 _7298_ (
    .a(_2395_),
    .b(_2719_),
    .c(_2392_),
    .y(_2745_)
  );
  al_nand2 _7299_ (
    .a(_1912_),
    .b(_2295_),
    .y(_2746_)
  );
  al_and3ftt _7300_ (
    .a(_1912_),
    .b(_0273_),
    .c(_1198_),
    .y(_2747_)
  );
  al_and2ft _7301_ (
    .a(_2747_),
    .b(_2746_),
    .y(_2748_)
  );
  al_and3 _7302_ (
    .a(_2358_),
    .b(_2748_),
    .c(_2745_),
    .y(_2749_)
  );
  al_ao21 _7303_ (
    .a(_2748_),
    .b(_2745_),
    .c(_2358_),
    .y(_2750_)
  );
  al_nand2ft _7304_ (
    .a(_2749_),
    .b(_2750_),
    .y(_2751_)
  );
  al_nand3 _7305_ (
    .a(_2369_),
    .b(_2751_),
    .c(_2709_),
    .y(_2752_)
  );
  al_nand3 _7306_ (
    .a(\DFF_1427.Q ),
    .b(_2752_),
    .c(_2744_),
    .y(_2753_)
  );
  al_ao21ftf _7307_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_233.Q ),
    .c(_2753_),
    .y(\DFF_233.D )
  );
  al_nand3 _7308_ (
    .a(\DFF_1428.Q ),
    .b(_2752_),
    .c(_2744_),
    .y(_2754_)
  );
  al_ao21ftf _7309_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_234.Q ),
    .c(_2754_),
    .y(\DFF_234.D )
  );
  al_nand3 _7310_ (
    .a(\DFF_1429.Q ),
    .b(_2752_),
    .c(_2744_),
    .y(_2755_)
  );
  al_ao21ftf _7311_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_235.Q ),
    .c(_2755_),
    .y(\DFF_235.D )
  );
  al_and3 _7312_ (
    .a(_0833_),
    .b(_0839_),
    .c(_0814_),
    .y(_2756_)
  );
  al_aoi21ftt _7313_ (
    .a(_0800_),
    .b(_0799_),
    .c(_0789_),
    .y(_2757_)
  );
  al_and3 _7314_ (
    .a(_0818_),
    .b(_0819_),
    .c(_0795_),
    .y(_2758_)
  );
  al_or2 _7315_ (
    .a(_0161_),
    .b(_0823_),
    .y(_2759_)
  );
  al_nand3ftt _7316_ (
    .a(_0805_),
    .b(_0806_),
    .c(_2759_),
    .y(_2760_)
  );
  al_aoi21 _7317_ (
    .a(_0161_),
    .b(_0823_),
    .c(_0848_),
    .y(_2761_)
  );
  al_nor3ftt _7318_ (
    .a(_2761_),
    .b(_2337_),
    .c(_2760_),
    .y(_2762_)
  );
  al_and3 _7319_ (
    .a(_2757_),
    .b(_2758_),
    .c(_2762_),
    .y(_2763_)
  );
  al_and3 _7320_ (
    .a(_2756_),
    .b(_2347_),
    .c(_2763_),
    .y(_2764_)
  );
  al_and3ftt _7321_ (
    .a(_2649_),
    .b(_2764_),
    .c(_1965_),
    .y(_2765_)
  );
  al_or3 _7322_ (
    .a(_0270_),
    .b(_1793_),
    .c(_2764_),
    .y(_2766_)
  );
  al_nand3 _7323_ (
    .a(_0270_),
    .b(_2296_),
    .c(_2650_),
    .y(_2767_)
  );
  al_ao21 _7324_ (
    .a(_2766_),
    .b(_2767_),
    .c(_2765_),
    .y(_2768_)
  );
  al_ao21 _7325_ (
    .a(_0267_),
    .b(_2768_),
    .c(_0273_),
    .y(_2769_)
  );
  al_nand2 _7326_ (
    .a(_0267_),
    .b(_0273_),
    .y(_2770_)
  );
  al_or3fft _7327_ (
    .a(_0270_),
    .b(_1955_),
    .c(_2649_),
    .y(_2771_)
  );
  al_nand3 _7328_ (
    .a(_0273_),
    .b(_1965_),
    .c(_2771_),
    .y(_2772_)
  );
  al_nand3fft _7329_ (
    .a(_1198_),
    .b(_2299_),
    .c(_2772_),
    .y(_2773_)
  );
  al_aoi21 _7330_ (
    .a(_2770_),
    .b(_2769_),
    .c(_2773_),
    .y(_2774_)
  );
  al_mux2h _7331_ (
    .a(\DFF_286.Q ),
    .b(_2774_),
    .s(\DFF_1427.Q ),
    .y(\DFF_286.D )
  );
  al_mux2h _7332_ (
    .a(\DFF_287.Q ),
    .b(_2774_),
    .s(\DFF_1428.Q ),
    .y(\DFF_287.D )
  );
  al_mux2h _7333_ (
    .a(\DFF_288.Q ),
    .b(_2774_),
    .s(\DFF_1429.Q ),
    .y(\DFF_288.D )
  );
  al_nand2 _7334_ (
    .a(_2420_),
    .b(_2429_),
    .y(_2775_)
  );
  al_and3 _7335_ (
    .a(_2450_),
    .b(_2420_),
    .c(_2429_),
    .y(_2776_)
  );
  al_ao21 _7336_ (
    .a(\DFF_58.Q ),
    .b(_2775_),
    .c(_2776_),
    .y(_2777_)
  );
  al_or2ft _7337_ (
    .a(_2441_),
    .b(_2464_),
    .y(_2778_)
  );
  al_nand2ft _7338_ (
    .a(_2441_),
    .b(_2464_),
    .y(_2779_)
  );
  al_nand3 _7339_ (
    .a(_2778_),
    .b(_2779_),
    .c(_2453_),
    .y(_2780_)
  );
  al_nand3 _7340_ (
    .a(\DFF_1427.Q ),
    .b(_2780_),
    .c(_2777_),
    .y(_2781_)
  );
  al_ao21ftf _7341_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_562.Q ),
    .c(_2781_),
    .y(\DFF_562.D )
  );
  al_nand3 _7342_ (
    .a(\DFF_1428.Q ),
    .b(_2780_),
    .c(_2777_),
    .y(_2782_)
  );
  al_ao21ftf _7343_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_563.Q ),
    .c(_2782_),
    .y(\DFF_563.D )
  );
  al_nand3 _7344_ (
    .a(\DFF_1429.Q ),
    .b(_2780_),
    .c(_2777_),
    .y(_2783_)
  );
  al_ao21ftf _7345_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_564.Q ),
    .c(_2783_),
    .y(\DFF_564.D )
  );
  al_ao21 _7346_ (
    .a(_0913_),
    .b(_2775_),
    .c(_2776_),
    .y(_2784_)
  );
  al_mux2h _7347_ (
    .a(_2490_),
    .b(_2491_),
    .s(_2435_),
    .y(_2785_)
  );
  al_ao21ttf _7348_ (
    .a(_2785_),
    .b(_2489_),
    .c(_2447_),
    .y(_2786_)
  );
  al_nand3ftt _7349_ (
    .a(_2447_),
    .b(_2785_),
    .c(_2489_),
    .y(_2787_)
  );
  al_nand3 _7350_ (
    .a(_2786_),
    .b(_2787_),
    .c(_2453_),
    .y(_2788_)
  );
  al_nand3 _7351_ (
    .a(\DFF_1427.Q ),
    .b(_2788_),
    .c(_2784_),
    .y(_2789_)
  );
  al_ao21ftf _7352_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_580.Q ),
    .c(_2789_),
    .y(\DFF_580.D )
  );
  al_nand3 _7353_ (
    .a(\DFF_1428.Q ),
    .b(_2788_),
    .c(_2784_),
    .y(_2790_)
  );
  al_ao21ftf _7354_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_581.Q ),
    .c(_2790_),
    .y(\DFF_581.D )
  );
  al_nand3 _7355_ (
    .a(\DFF_1429.Q ),
    .b(_2788_),
    .c(_2784_),
    .y(_2791_)
  );
  al_ao21ftf _7356_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_582.Q ),
    .c(_2791_),
    .y(\DFF_582.D )
  );
  al_ao21 _7357_ (
    .a(\DFF_60.Q ),
    .b(_2775_),
    .c(_2776_),
    .y(_2792_)
  );
  al_inv _7358_ (
    .a(_2440_),
    .y(_2793_)
  );
  al_nand2 _7359_ (
    .a(_2793_),
    .b(_2461_),
    .y(_2794_)
  );
  al_or3fft _7360_ (
    .a(_2006_),
    .b(_2008_),
    .c(_2461_),
    .y(_2795_)
  );
  al_nand3 _7361_ (
    .a(_2794_),
    .b(_2795_),
    .c(_2453_),
    .y(_2796_)
  );
  al_nand3 _7362_ (
    .a(\DFF_1427.Q ),
    .b(_2796_),
    .c(_2792_),
    .y(_2797_)
  );
  al_ao21ftf _7363_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_559.Q ),
    .c(_2797_),
    .y(\DFF_559.D )
  );
  al_nand3 _7364_ (
    .a(\DFF_1428.Q ),
    .b(_2796_),
    .c(_2792_),
    .y(_2798_)
  );
  al_ao21ftf _7365_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_560.Q ),
    .c(_2798_),
    .y(\DFF_560.D )
  );
  al_nand3 _7366_ (
    .a(\DFF_1429.Q ),
    .b(_2796_),
    .c(_2792_),
    .y(_2799_)
  );
  al_ao21ftf _7367_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_561.Q ),
    .c(_2799_),
    .y(\DFF_561.D )
  );
  al_ao21 _7368_ (
    .a(\DFF_56.Q ),
    .b(_2775_),
    .c(_2776_),
    .y(_2800_)
  );
  al_nand3ftt _7369_ (
    .a(_2439_),
    .b(_2473_),
    .c(_2464_),
    .y(_2801_)
  );
  al_ao21ttf _7370_ (
    .a(_2473_),
    .b(_2464_),
    .c(_2439_),
    .y(_2802_)
  );
  al_nand3 _7371_ (
    .a(_2801_),
    .b(_2802_),
    .c(_2453_),
    .y(_2803_)
  );
  al_nand3 _7372_ (
    .a(\DFF_1427.Q ),
    .b(_2803_),
    .c(_2800_),
    .y(_2804_)
  );
  al_ao21ftf _7373_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_565.Q ),
    .c(_2804_),
    .y(\DFF_565.D )
  );
  al_nand3 _7374_ (
    .a(\DFF_1428.Q ),
    .b(_2803_),
    .c(_2800_),
    .y(_2805_)
  );
  al_ao21ftf _7375_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_566.Q ),
    .c(_2805_),
    .y(\DFF_566.D )
  );
  al_nand3 _7376_ (
    .a(\DFF_1429.Q ),
    .b(_2803_),
    .c(_2800_),
    .y(_2806_)
  );
  al_ao21ftf _7377_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_567.Q ),
    .c(_2806_),
    .y(\DFF_567.D )
  );
  al_ao21 _7378_ (
    .a(_0917_),
    .b(_2775_),
    .c(_2776_),
    .y(_2807_)
  );
  al_nand2 _7379_ (
    .a(_2447_),
    .b(_2302_),
    .y(_2808_)
  );
  al_nor3fft _7380_ (
    .a(_2019_),
    .b(_2021_),
    .c(_2302_),
    .y(_2809_)
  );
  al_nor2ft _7381_ (
    .a(_2808_),
    .b(_2809_),
    .y(_2810_)
  );
  al_nand3 _7382_ (
    .a(_2785_),
    .b(_2810_),
    .c(_2489_),
    .y(_2811_)
  );
  al_or3fft _7383_ (
    .a(_2013_),
    .b(_2015_),
    .c(_2811_),
    .y(_2812_)
  );
  al_nand2 _7384_ (
    .a(_2443_),
    .b(_2811_),
    .y(_2813_)
  );
  al_nand3 _7385_ (
    .a(_2812_),
    .b(_2813_),
    .c(_2453_),
    .y(_2814_)
  );
  al_nand3 _7386_ (
    .a(\DFF_1427.Q ),
    .b(_2814_),
    .c(_2807_),
    .y(_2815_)
  );
  al_ao21ftf _7387_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_583.Q ),
    .c(_2815_),
    .y(\DFF_583.D )
  );
  al_nand3 _7388_ (
    .a(\DFF_1428.Q ),
    .b(_2814_),
    .c(_2807_),
    .y(_2816_)
  );
  al_ao21ftf _7389_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_584.Q ),
    .c(_2816_),
    .y(\DFF_584.D )
  );
  al_nand3 _7390_ (
    .a(\DFF_1429.Q ),
    .b(_2814_),
    .c(_2807_),
    .y(_2817_)
  );
  al_ao21ftf _7391_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_585.Q ),
    .c(_2817_),
    .y(\DFF_585.D )
  );
  al_nand3 _7392_ (
    .a(_0863_),
    .b(_2426_),
    .c(_2424_),
    .y(_2818_)
  );
  al_nand2 _7393_ (
    .a(\DFF_1302.Q ),
    .b(_0926_),
    .y(_2819_)
  );
  al_and3 _7394_ (
    .a(_2418_),
    .b(_0882_),
    .c(_0929_),
    .y(_2820_)
  );
  al_oa21ftf _7395_ (
    .a(_2819_),
    .b(_2820_),
    .c(_0291_),
    .y(_2821_)
  );
  al_inv _7396_ (
    .a(_0287_),
    .y(_2822_)
  );
  al_nand3 _7397_ (
    .a(_0284_),
    .b(_2658_),
    .c(_2048_),
    .y(_2823_)
  );
  al_aoi21 _7398_ (
    .a(_2061_),
    .b(_2823_),
    .c(_2822_),
    .y(_2824_)
  );
  al_oa21 _7399_ (
    .a(_2050_),
    .b(_2048_),
    .c(_2663_),
    .y(_2825_)
  );
  al_nand3 _7400_ (
    .a(_2820_),
    .b(_2658_),
    .c(_2061_),
    .y(_2826_)
  );
  al_ao21 _7401_ (
    .a(_2826_),
    .b(_2825_),
    .c(_2421_),
    .y(_2827_)
  );
  al_nand3fft _7402_ (
    .a(_2821_),
    .b(_2824_),
    .c(_2827_),
    .y(_2828_)
  );
  al_nand3fft _7403_ (
    .a(_0281_),
    .b(_0287_),
    .c(_2828_),
    .y(_2829_)
  );
  al_ao21ttf _7404_ (
    .a(_2061_),
    .b(_2823_),
    .c(_0287_),
    .y(_2830_)
  );
  al_ao21ftt _7405_ (
    .a(_2821_),
    .b(_2830_),
    .c(_0281_),
    .y(_2831_)
  );
  al_or3ftt _7406_ (
    .a(_0284_),
    .b(_0281_),
    .c(_0287_),
    .y(_2832_)
  );
  al_ao21 _7407_ (
    .a(_2826_),
    .b(_2825_),
    .c(_2832_),
    .y(_2833_)
  );
  al_ao21 _7408_ (
    .a(_0281_),
    .b(_0284_),
    .c(_0287_),
    .y(_2834_)
  );
  al_nand3 _7409_ (
    .a(_2833_),
    .b(_2834_),
    .c(_2831_),
    .y(_2835_)
  );
  al_and3 _7410_ (
    .a(_2818_),
    .b(_2835_),
    .c(_2829_),
    .y(_2836_)
  );
  al_mux2h _7411_ (
    .a(\DFF_636.Q ),
    .b(_2836_),
    .s(\DFF_1427.Q ),
    .y(\DFF_636.D )
  );
  al_mux2h _7412_ (
    .a(\DFF_637.Q ),
    .b(_2836_),
    .s(\DFF_1428.Q ),
    .y(\DFF_637.D )
  );
  al_mux2h _7413_ (
    .a(\DFF_638.Q ),
    .b(_2836_),
    .s(\DFF_1429.Q ),
    .y(\DFF_638.D )
  );
  al_nand3 _7414_ (
    .a(_2497_),
    .b(_2505_),
    .c(_2504_),
    .y(_2837_)
  );
  al_mux2l _7415_ (
    .a(\DFF_43.Q ),
    .b(_2521_),
    .s(_2837_),
    .y(_2838_)
  );
  al_and3ftt _7416_ (
    .a(_2518_),
    .b(_2535_),
    .c(_2545_),
    .y(_2839_)
  );
  al_or3fft _7417_ (
    .a(_2115_),
    .b(_2117_),
    .c(_2536_),
    .y(_2840_)
  );
  al_nand2ft _7418_ (
    .a(_2839_),
    .b(_2840_),
    .y(_2841_)
  );
  al_nand3 _7419_ (
    .a(_2527_),
    .b(_2841_),
    .c(_2506_),
    .y(_2842_)
  );
  al_nand3 _7420_ (
    .a(\DFF_1427.Q ),
    .b(_2842_),
    .c(_2838_),
    .y(_2843_)
  );
  al_ao21ftf _7421_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_912.Q ),
    .c(_2843_),
    .y(\DFF_912.D )
  );
  al_nand3 _7422_ (
    .a(\DFF_1428.Q ),
    .b(_2842_),
    .c(_2838_),
    .y(_2844_)
  );
  al_ao21ftf _7423_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_913.Q ),
    .c(_2844_),
    .y(\DFF_913.D )
  );
  al_nand3 _7424_ (
    .a(\DFF_1429.Q ),
    .b(_2842_),
    .c(_2838_),
    .y(_2845_)
  );
  al_ao21ftf _7425_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_914.Q ),
    .c(_2845_),
    .y(\DFF_914.D )
  );
  al_mux2l _7426_ (
    .a(_0953_),
    .b(_2521_),
    .s(_2837_),
    .y(_2846_)
  );
  al_ao21 _7427_ (
    .a(_2510_),
    .b(_2516_),
    .c(_2508_),
    .y(_2847_)
  );
  al_aoi21ttf _7428_ (
    .a(_2508_),
    .b(_2563_),
    .c(_2847_),
    .y(_2848_)
  );
  al_and3 _7429_ (
    .a(_2515_),
    .b(_2848_),
    .c(_2551_),
    .y(_2849_)
  );
  al_ao21 _7430_ (
    .a(_2848_),
    .b(_2551_),
    .c(_2515_),
    .y(_2850_)
  );
  al_nand2ft _7431_ (
    .a(_2849_),
    .b(_2850_),
    .y(_2851_)
  );
  al_nand3 _7432_ (
    .a(_2527_),
    .b(_2851_),
    .c(_2506_),
    .y(_2852_)
  );
  al_nand3 _7433_ (
    .a(\DFF_1427.Q ),
    .b(_2852_),
    .c(_2846_),
    .y(_2853_)
  );
  al_ao21ftf _7434_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_930.Q ),
    .c(_2853_),
    .y(\DFF_930.D )
  );
  al_nand3 _7435_ (
    .a(\DFF_1428.Q ),
    .b(_2852_),
    .c(_2846_),
    .y(_2854_)
  );
  al_ao21ftf _7436_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_931.Q ),
    .c(_2854_),
    .y(\DFF_931.D )
  );
  al_nand3 _7437_ (
    .a(\DFF_1429.Q ),
    .b(_2852_),
    .c(_2846_),
    .y(_2855_)
  );
  al_ao21ftf _7438_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_932.Q ),
    .c(_2855_),
    .y(\DFF_932.D )
  );
  al_mux2l _7439_ (
    .a(\DFF_44.Q ),
    .b(_2521_),
    .s(_2837_),
    .y(_2856_)
  );
  al_or3fft _7440_ (
    .a(_2097_),
    .b(_2099_),
    .c(_2535_),
    .y(_2857_)
  );
  al_and2 _7441_ (
    .a(_2514_),
    .b(_2535_),
    .y(_2858_)
  );
  al_nand2ft _7442_ (
    .a(_2858_),
    .b(_2857_),
    .y(_2859_)
  );
  al_nand3 _7443_ (
    .a(_2527_),
    .b(_2859_),
    .c(_2506_),
    .y(_2860_)
  );
  al_nand3 _7444_ (
    .a(\DFF_1427.Q ),
    .b(_2860_),
    .c(_2856_),
    .y(_2861_)
  );
  al_ao21ftf _7445_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_909.Q ),
    .c(_2861_),
    .y(\DFF_909.D )
  );
  al_nand3 _7446_ (
    .a(\DFF_1428.Q ),
    .b(_2860_),
    .c(_2856_),
    .y(_2862_)
  );
  al_ao21ftf _7447_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_910.Q ),
    .c(_2862_),
    .y(\DFF_910.D )
  );
  al_nand3 _7448_ (
    .a(\DFF_1429.Q ),
    .b(_2860_),
    .c(_2856_),
    .y(_2863_)
  );
  al_ao21ftf _7449_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_911.Q ),
    .c(_2863_),
    .y(\DFF_911.D )
  );
  al_mux2l _7450_ (
    .a(\DFF_42.Q ),
    .b(_2521_),
    .s(_2837_),
    .y(_2864_)
  );
  al_oai21 _7451_ (
    .a(_2537_),
    .b(_2538_),
    .c(_2536_),
    .y(_2865_)
  );
  al_or2ft _7452_ (
    .a(_2519_),
    .b(_2865_),
    .y(_2866_)
  );
  al_and2ft _7453_ (
    .a(_2519_),
    .b(_2865_),
    .y(_2867_)
  );
  al_and2ft _7454_ (
    .a(_2867_),
    .b(_2866_),
    .y(_2868_)
  );
  al_nand3 _7455_ (
    .a(_2527_),
    .b(_2868_),
    .c(_2506_),
    .y(_2869_)
  );
  al_nand3 _7456_ (
    .a(\DFF_1427.Q ),
    .b(_2869_),
    .c(_2864_),
    .y(_2870_)
  );
  al_ao21ftf _7457_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_915.Q ),
    .c(_2870_),
    .y(\DFF_915.D )
  );
  al_nand3 _7458_ (
    .a(\DFF_1428.Q ),
    .b(_2869_),
    .c(_2864_),
    .y(_2871_)
  );
  al_ao21ftf _7459_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_916.Q ),
    .c(_2871_),
    .y(\DFF_916.D )
  );
  al_nand3 _7460_ (
    .a(\DFF_1429.Q ),
    .b(_2869_),
    .c(_2864_),
    .y(_2872_)
  );
  al_ao21ftf _7461_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_917.Q ),
    .c(_2872_),
    .y(\DFF_917.D )
  );
  al_mux2l _7462_ (
    .a(_1833_),
    .b(_2521_),
    .s(_2837_),
    .y(_2873_)
  );
  al_nand2 _7463_ (
    .a(_2515_),
    .b(_2308_),
    .y(_2874_)
  );
  al_and3ftt _7464_ (
    .a(_2515_),
    .b(_0304_),
    .c(_2524_),
    .y(_2875_)
  );
  al_and2ft _7465_ (
    .a(_2875_),
    .b(_2874_),
    .y(_2876_)
  );
  al_nand3 _7466_ (
    .a(_2848_),
    .b(_2876_),
    .c(_2551_),
    .y(_2877_)
  );
  al_or2ft _7467_ (
    .a(_2143_),
    .b(_2877_),
    .y(_2878_)
  );
  al_and2ft _7468_ (
    .a(_2143_),
    .b(_2877_),
    .y(_2879_)
  );
  al_nand2ft _7469_ (
    .a(_2879_),
    .b(_2878_),
    .y(_2880_)
  );
  al_nand3 _7470_ (
    .a(_2527_),
    .b(_2880_),
    .c(_2506_),
    .y(_2881_)
  );
  al_nand3 _7471_ (
    .a(\DFF_1427.Q ),
    .b(_2881_),
    .c(_2873_),
    .y(_2882_)
  );
  al_ao21ftf _7472_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_933.Q ),
    .c(_2882_),
    .y(\DFF_933.D )
  );
  al_nand3 _7473_ (
    .a(\DFF_1428.Q ),
    .b(_2881_),
    .c(_2873_),
    .y(_2883_)
  );
  al_ao21ftf _7474_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_934.Q ),
    .c(_2883_),
    .y(\DFF_934.D )
  );
  al_nand3 _7475_ (
    .a(\DFF_1429.Q ),
    .b(_2881_),
    .c(_2873_),
    .y(_2884_)
  );
  al_ao21ftf _7476_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_935.Q ),
    .c(_2884_),
    .y(\DFF_935.D )
  );
  al_nand2 _7477_ (
    .a(_0941_),
    .b(_1010_),
    .y(_2885_)
  );
  al_nand3 _7478_ (
    .a(_0301_),
    .b(_2161_),
    .c(_2671_),
    .y(_2886_)
  );
  al_ao21ttf _7479_ (
    .a(_2172_),
    .b(_2886_),
    .c(_0304_),
    .y(_2887_)
  );
  al_oai21ftf _7480_ (
    .a(_1837_),
    .b(_2502_),
    .c(_2150_),
    .y(_2888_)
  );
  al_ao21 _7481_ (
    .a(_2888_),
    .b(_2887_),
    .c(_0298_),
    .y(_2889_)
  );
  al_or3 _7482_ (
    .a(_0298_),
    .b(_0306_),
    .c(_0304_),
    .y(_2890_)
  );
  al_aoi21ftf _7483_ (
    .a(_1102_),
    .b(_2148_),
    .c(_2162_),
    .y(_2891_)
  );
  al_and3 _7484_ (
    .a(_2501_),
    .b(_2687_),
    .c(_2671_),
    .y(_2892_)
  );
  al_nand3 _7485_ (
    .a(_2172_),
    .b(_2162_),
    .c(_2892_),
    .y(_2893_)
  );
  al_ao21 _7486_ (
    .a(_2891_),
    .b(_2893_),
    .c(_2890_),
    .y(_2894_)
  );
  al_ao21 _7487_ (
    .a(_2894_),
    .b(_2889_),
    .c(_0304_),
    .y(_2895_)
  );
  al_ao21 _7488_ (
    .a(_0298_),
    .b(_0301_),
    .c(_0304_),
    .y(_2896_)
  );
  al_nand3 _7489_ (
    .a(_2896_),
    .b(_2894_),
    .c(_2889_),
    .y(_2897_)
  );
  al_and3 _7490_ (
    .a(_2885_),
    .b(_2897_),
    .c(_2895_),
    .y(_2898_)
  );
  al_mux2h _7491_ (
    .a(\DFF_986.Q ),
    .b(_2898_),
    .s(\DFF_1427.Q ),
    .y(\DFF_986.D )
  );
  al_mux2h _7492_ (
    .a(\DFF_987.Q ),
    .b(_2898_),
    .s(\DFF_1428.Q ),
    .y(\DFF_987.D )
  );
  al_mux2h _7493_ (
    .a(\DFF_988.Q ),
    .b(_2898_),
    .s(\DFF_1429.Q ),
    .y(\DFF_988.D )
  );
  al_nand2 _7494_ (
    .a(_2576_),
    .b(_2586_),
    .y(_2899_)
  );
  al_and3 _7495_ (
    .a(_2601_),
    .b(_2576_),
    .c(_2586_),
    .y(_2900_)
  );
  al_ao21 _7496_ (
    .a(\DFF_88.Q ),
    .b(_2899_),
    .c(_2900_),
    .y(_2901_)
  );
  al_or2ft _7497_ (
    .a(_2592_),
    .b(_2615_),
    .y(_2902_)
  );
  al_nand2ft _7498_ (
    .a(_2592_),
    .b(_2615_),
    .y(_2903_)
  );
  al_nand3 _7499_ (
    .a(_2902_),
    .b(_2903_),
    .c(_2604_),
    .y(_2904_)
  );
  al_nand3 _7500_ (
    .a(\DFF_1427.Q ),
    .b(_2904_),
    .c(_2901_),
    .y(_2905_)
  );
  al_ao21ftf _7501_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_1262.Q ),
    .c(_2905_),
    .y(\DFF_1262.D )
  );
  al_nand3 _7502_ (
    .a(\DFF_1428.Q ),
    .b(_2904_),
    .c(_2901_),
    .y(_2906_)
  );
  al_ao21ftf _7503_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_1263.Q ),
    .c(_2906_),
    .y(\DFF_1263.D )
  );
  al_nand3 _7504_ (
    .a(\DFF_1429.Q ),
    .b(_2904_),
    .c(_2901_),
    .y(_2907_)
  );
  al_ao21ftf _7505_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_1264.Q ),
    .c(_2907_),
    .y(\DFF_1264.D )
  );
  al_ao21 _7506_ (
    .a(_0236_),
    .b(_2899_),
    .c(_2900_),
    .y(_2908_)
  );
  al_nand3 _7507_ (
    .a(_2588_),
    .b(_2589_),
    .c(_2321_),
    .y(_2909_)
  );
  al_ao21ftf _7508_ (
    .a(_2589_),
    .b(_2642_),
    .c(_2909_),
    .y(_2910_)
  );
  al_nand3ftt _7509_ (
    .a(_2190_),
    .b(_2910_),
    .c(_2640_),
    .y(_2911_)
  );
  al_ao21ttf _7510_ (
    .a(_2910_),
    .b(_2640_),
    .c(_2190_),
    .y(_2912_)
  );
  al_nand3 _7511_ (
    .a(_2911_),
    .b(_2912_),
    .c(_2604_),
    .y(_2913_)
  );
  al_nand3 _7512_ (
    .a(\DFF_1427.Q ),
    .b(_2913_),
    .c(_2908_),
    .y(_2914_)
  );
  al_ao21ftf _7513_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_1280.Q ),
    .c(_2914_),
    .y(\DFF_1280.D )
  );
  al_nand3 _7514_ (
    .a(\DFF_1428.Q ),
    .b(_2913_),
    .c(_2908_),
    .y(_2915_)
  );
  al_ao21ftf _7515_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_1281.Q ),
    .c(_2915_),
    .y(\DFF_1281.D )
  );
  al_nand3 _7516_ (
    .a(\DFF_1429.Q ),
    .b(_2913_),
    .c(_2908_),
    .y(_2916_)
  );
  al_ao21ftf _7517_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_1282.Q ),
    .c(_2916_),
    .y(\DFF_1282.D )
  );
  al_ao21 _7518_ (
    .a(\DFF_89.Q ),
    .b(_2899_),
    .c(_2900_),
    .y(_2917_)
  );
  al_or2 _7519_ (
    .a(_2204_),
    .b(_2612_),
    .y(_2918_)
  );
  al_nand2 _7520_ (
    .a(_2204_),
    .b(_2612_),
    .y(_2919_)
  );
  al_nand3 _7521_ (
    .a(_2918_),
    .b(_2919_),
    .c(_2604_),
    .y(_2920_)
  );
  al_nand3 _7522_ (
    .a(\DFF_1427.Q ),
    .b(_2920_),
    .c(_2917_),
    .y(_2921_)
  );
  al_ao21ftf _7523_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_1259.Q ),
    .c(_2921_),
    .y(\DFF_1259.D )
  );
  al_nand3 _7524_ (
    .a(\DFF_1428.Q ),
    .b(_2920_),
    .c(_2917_),
    .y(_2922_)
  );
  al_ao21ftf _7525_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_1260.Q ),
    .c(_2922_),
    .y(\DFF_1260.D )
  );
  al_nand3 _7526_ (
    .a(\DFF_1429.Q ),
    .b(_2920_),
    .c(_2917_),
    .y(_2923_)
  );
  al_ao21ftf _7527_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_1261.Q ),
    .c(_2923_),
    .y(\DFF_1261.D )
  );
  al_ao21 _7528_ (
    .a(\DFF_87.Q ),
    .b(_2899_),
    .c(_2900_),
    .y(_2924_)
  );
  al_nand3ftt _7529_ (
    .a(_2593_),
    .b(_2624_),
    .c(_2615_),
    .y(_2925_)
  );
  al_ao21ttf _7530_ (
    .a(_2624_),
    .b(_2615_),
    .c(_2593_),
    .y(_2926_)
  );
  al_nand3 _7531_ (
    .a(_2925_),
    .b(_2926_),
    .c(_2604_),
    .y(_2927_)
  );
  al_nand3 _7532_ (
    .a(\DFF_1427.Q ),
    .b(_2927_),
    .c(_2924_),
    .y(_2928_)
  );
  al_ao21ftf _7533_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_1265.Q ),
    .c(_2928_),
    .y(\DFF_1265.D )
  );
  al_nand3 _7534_ (
    .a(\DFF_1428.Q ),
    .b(_2927_),
    .c(_2924_),
    .y(_2929_)
  );
  al_ao21ftf _7535_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_1266.Q ),
    .c(_2929_),
    .y(\DFF_1266.D )
  );
  al_nand3 _7536_ (
    .a(\DFF_1429.Q ),
    .b(_2927_),
    .c(_2924_),
    .y(_2930_)
  );
  al_ao21ftf _7537_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_1267.Q ),
    .c(_2930_),
    .y(\DFF_1267.D )
  );
  al_ao21 _7538_ (
    .a(_0240_),
    .b(_2899_),
    .c(_2900_),
    .y(_2931_)
  );
  al_nand2 _7539_ (
    .a(_2190_),
    .b(_2321_),
    .y(_2932_)
  );
  al_and3ftt _7540_ (
    .a(_2190_),
    .b(_0320_),
    .c(_1387_),
    .y(_2933_)
  );
  al_and2ft _7541_ (
    .a(_2933_),
    .b(_2932_),
    .y(_2934_)
  );
  al_nand3 _7542_ (
    .a(_2910_),
    .b(_2934_),
    .c(_2640_),
    .y(_2935_)
  );
  al_or3fft _7543_ (
    .a(_2245_),
    .b(_2247_),
    .c(_2935_),
    .y(_2936_)
  );
  al_nand2 _7544_ (
    .a(_2594_),
    .b(_2935_),
    .y(_2937_)
  );
  al_nand3 _7545_ (
    .a(_2936_),
    .b(_2937_),
    .c(_2604_),
    .y(_2938_)
  );
  al_nand3 _7546_ (
    .a(\DFF_1427.Q ),
    .b(_2938_),
    .c(_2931_),
    .y(_2939_)
  );
  al_ao21ftf _7547_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_1283.Q ),
    .c(_2939_),
    .y(\DFF_1283.D )
  );
  al_nand3 _7548_ (
    .a(\DFF_1428.Q ),
    .b(_2938_),
    .c(_2931_),
    .y(_2940_)
  );
  al_ao21ftf _7549_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_1284.Q ),
    .c(_2940_),
    .y(\DFF_1284.D )
  );
  al_nand3 _7550_ (
    .a(\DFF_1429.Q ),
    .b(_2938_),
    .c(_2931_),
    .y(_2941_)
  );
  al_ao21ftf _7551_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_1285.Q ),
    .c(_2941_),
    .y(\DFF_1285.D )
  );
  al_and3 _7552_ (
    .a(_0317_),
    .b(_2265_),
    .c(_2263_),
    .y(_2942_)
  );
  al_nand3 _7553_ (
    .a(_1085_),
    .b(_2252_),
    .c(_2942_),
    .y(_2943_)
  );
  al_and2 _7554_ (
    .a(_0320_),
    .b(_2275_),
    .y(_2944_)
  );
  al_aoi21ftf _7555_ (
    .a(_1079_),
    .b(\DFF_88.Q ),
    .c(_1022_),
    .y(_2945_)
  );
  al_and3 _7556_ (
    .a(_2945_),
    .b(_1050_),
    .c(_1070_),
    .y(_2946_)
  );
  al_aoi21ftf _7557_ (
    .a(_1028_),
    .b(_0236_),
    .c(_1041_),
    .y(_2947_)
  );
  al_and3 _7558_ (
    .a(_1042_),
    .b(_1030_),
    .c(_2947_),
    .y(_2948_)
  );
  al_oa21 _7559_ (
    .a(_0240_),
    .b(_1053_),
    .c(_1081_),
    .y(_2949_)
  );
  al_and3ftt _7560_ (
    .a(_1023_),
    .b(_1055_),
    .c(_2949_),
    .y(_2950_)
  );
  al_nand2 _7561_ (
    .a(\DFF_84.Q ),
    .b(_1059_),
    .y(_2951_)
  );
  al_nand2 _7562_ (
    .a(\DFF_1350.D ),
    .b(_1061_),
    .y(_2952_)
  );
  al_and3ftt _7563_ (
    .a(_2256_),
    .b(_2951_),
    .c(_2952_),
    .y(_2953_)
  );
  al_and3 _7564_ (
    .a(_1036_),
    .b(_2953_),
    .c(_1076_),
    .y(_2954_)
  );
  al_and3 _7565_ (
    .a(_2948_),
    .b(_2950_),
    .c(_2954_),
    .y(_2955_)
  );
  al_nand3 _7566_ (
    .a(_1018_),
    .b(_2946_),
    .c(_2955_),
    .y(_2956_)
  );
  al_ao21ftf _7567_ (
    .a(_0314_),
    .b(_2255_),
    .c(_2956_),
    .y(_2957_)
  );
  al_ao21 _7568_ (
    .a(_2943_),
    .b(_2944_),
    .c(_2957_),
    .y(_2958_)
  );
  al_ao21 _7569_ (
    .a(_2698_),
    .b(_2266_),
    .c(_2697_),
    .y(_2959_)
  );
  al_and3 _7570_ (
    .a(_2946_),
    .b(_2574_),
    .c(_2955_),
    .y(_2960_)
  );
  al_oai21ftf _7571_ (
    .a(_1865_),
    .b(_2960_),
    .c(_0317_),
    .y(_2961_)
  );
  al_and3 _7572_ (
    .a(_1085_),
    .b(_2252_),
    .c(_2960_),
    .y(_2962_)
  );
  al_ao21ttf _7573_ (
    .a(_2275_),
    .b(_2962_),
    .c(_2961_),
    .y(_2963_)
  );
  al_ao21ttf _7574_ (
    .a(_0314_),
    .b(_2963_),
    .c(_2959_),
    .y(_2964_)
  );
  al_aoi21 _7575_ (
    .a(_2694_),
    .b(_2964_),
    .c(_2958_),
    .y(_2965_)
  );
  al_mux2h _7576_ (
    .a(\DFF_1336.Q ),
    .b(_2965_),
    .s(\DFF_1427.Q ),
    .y(\DFF_1336.D )
  );
  al_mux2h _7577_ (
    .a(\DFF_1337.Q ),
    .b(_2965_),
    .s(\DFF_1428.Q ),
    .y(\DFF_1337.D )
  );
  al_mux2h _7578_ (
    .a(\DFF_1338.Q ),
    .b(_2965_),
    .s(\DFF_1429.Q ),
    .y(\DFF_1338.D )
  );
  al_mux2h _7579_ (
    .a(\DFF_116.Q ),
    .b(\DFF_1450.D ),
    .s(\DFF_1504.Q ),
    .y(\DFF_116.D )
  );
  al_mux2h _7580_ (
    .a(\DFF_117.Q ),
    .b(\DFF_1450.D ),
    .s(\DFF_1505.Q ),
    .y(\DFF_117.D )
  );
  al_mux2h _7581_ (
    .a(\DFF_118.Q ),
    .b(\DFF_1450.D ),
    .s(\DFF_1506.Q ),
    .y(\DFF_118.D )
  );
  al_oai21ftt _7582_ (
    .a(\DFF_1611.Q ),
    .b(\DFF_1612.Q ),
    .c(\DFF_1613.Q ),
    .y(\DFF_1613.D )
  );
  al_oai21ftt _7583_ (
    .a(\DFF_17.Q ),
    .b(\DFF_18.Q ),
    .c(\DFF_19.Q ),
    .y(\DFF_19.D )
  );
  al_inv _7584_ (
    .a(\DFF_29.Q ),
    .y(_2966_)
  );
  al_ao21 _7585_ (
    .a(_0129_),
    .b(_0130_),
    .c(_2966_),
    .y(_2967_)
  );
  al_and3 _7586_ (
    .a(_2966_),
    .b(_0129_),
    .c(_0130_),
    .y(_2968_)
  );
  al_nand2ft _7587_ (
    .a(_2968_),
    .b(_2967_),
    .y(\DFF_16.D )
  );
  al_inv _7588_ (
    .a(\DFF_20.Q ),
    .y(_2969_)
  );
  al_ao21 _7589_ (
    .a(_0150_),
    .b(_0151_),
    .c(_2969_),
    .y(_2970_)
  );
  al_and3 _7590_ (
    .a(_2969_),
    .b(_0150_),
    .c(_0151_),
    .y(_2971_)
  );
  al_nand2ft _7591_ (
    .a(_2971_),
    .b(_2970_),
    .y(\DFF_15.D )
  );
  al_and2ft _7592_ (
    .a(\DFF_1620.Q ),
    .b(\DFF_1621.Q ),
    .y(_2972_)
  );
  al_nand2ft _7593_ (
    .a(\DFF_1621.Q ),
    .b(\DFF_1620.Q ),
    .y(_2973_)
  );
  al_and2ft _7594_ (
    .a(\DFF_1619.Q ),
    .b(\DFF_1618.Q ),
    .y(_2974_)
  );
  al_nand2ft _7595_ (
    .a(\DFF_1618.Q ),
    .b(\DFF_1619.Q ),
    .y(_2975_)
  );
  al_nand2ft _7596_ (
    .a(_2974_),
    .b(_2975_),
    .y(_2976_)
  );
  al_aoi21ftf _7597_ (
    .a(_2972_),
    .b(_2973_),
    .c(_2976_),
    .y(_2977_)
  );
  al_and3fft _7598_ (
    .a(_2972_),
    .b(_2976_),
    .c(_2973_),
    .y(_2978_)
  );
  al_and2ft _7599_ (
    .a(\DFF_1615.Q ),
    .b(\DFF_1614.Q ),
    .y(_2979_)
  );
  al_nand2ft _7600_ (
    .a(\DFF_1614.Q ),
    .b(\DFF_1615.Q ),
    .y(_2980_)
  );
  al_and2ft _7601_ (
    .a(\DFF_1616.Q ),
    .b(\DFF_1617.Q ),
    .y(_2981_)
  );
  al_nand2ft _7602_ (
    .a(\DFF_1617.Q ),
    .b(\DFF_1616.Q ),
    .y(_2982_)
  );
  al_nand2ft _7603_ (
    .a(_2981_),
    .b(_2982_),
    .y(_2983_)
  );
  al_and3ftt _7604_ (
    .a(_2979_),
    .b(_2980_),
    .c(_2983_),
    .y(_2984_)
  );
  al_ao21ftt _7605_ (
    .a(_2979_),
    .b(_2980_),
    .c(_2983_),
    .y(_2985_)
  );
  al_nand2ft _7606_ (
    .a(_2984_),
    .b(_2985_),
    .y(_2986_)
  );
  al_or3 _7607_ (
    .a(_2977_),
    .b(_2978_),
    .c(_2986_),
    .y(_2987_)
  );
  al_oa21 _7608_ (
    .a(_2977_),
    .b(_2978_),
    .c(_2986_),
    .y(_2988_)
  );
  al_nand2ft _7609_ (
    .a(_2988_),
    .b(_2987_),
    .y(_2989_)
  );
  al_or3fft _7610_ (
    .a(\DFF_158.Q ),
    .b(_0113_),
    .c(_2989_),
    .y(_2990_)
  );
  al_inv _7611_ (
    .a(\DFF_158.Q ),
    .y(_2991_)
  );
  al_aoi21ftf _7612_ (
    .a(_2991_),
    .b(_0113_),
    .c(_2989_),
    .y(_2992_)
  );
  al_nand2ft _7613_ (
    .a(_2992_),
    .b(_2990_),
    .y(\DFF_1623.D )
  );
  al_and2ft _7614_ (
    .a(\DFF_1631.Q ),
    .b(\DFF_1629.Q ),
    .y(_2993_)
  );
  al_nand2ft _7615_ (
    .a(\DFF_1629.Q ),
    .b(\DFF_1631.Q ),
    .y(_2994_)
  );
  al_and2ft _7616_ (
    .a(\DFF_1630.Q ),
    .b(\DFF_1632.Q ),
    .y(_2995_)
  );
  al_nand2ft _7617_ (
    .a(\DFF_1632.Q ),
    .b(\DFF_1630.Q ),
    .y(_2996_)
  );
  al_nand2ft _7618_ (
    .a(_2995_),
    .b(_2996_),
    .y(_2997_)
  );
  al_aoi21ftf _7619_ (
    .a(_2993_),
    .b(_2994_),
    .c(_2997_),
    .y(_2998_)
  );
  al_and3fft _7620_ (
    .a(_2993_),
    .b(_2997_),
    .c(_2994_),
    .y(_2999_)
  );
  al_and2ft _7621_ (
    .a(\DFF_1626.Q ),
    .b(\DFF_1625.Q ),
    .y(_3000_)
  );
  al_nand2ft _7622_ (
    .a(\DFF_1625.Q ),
    .b(\DFF_1626.Q ),
    .y(_3001_)
  );
  al_and2ft _7623_ (
    .a(\DFF_1627.Q ),
    .b(\DFF_1628.Q ),
    .y(_3002_)
  );
  al_nand2ft _7624_ (
    .a(\DFF_1628.Q ),
    .b(\DFF_1627.Q ),
    .y(_3003_)
  );
  al_nand2ft _7625_ (
    .a(_3002_),
    .b(_3003_),
    .y(_3004_)
  );
  al_and3ftt _7626_ (
    .a(_3000_),
    .b(_3001_),
    .c(_3004_),
    .y(_3005_)
  );
  al_ao21ftt _7627_ (
    .a(_3000_),
    .b(_3001_),
    .c(_3004_),
    .y(_3006_)
  );
  al_nand2ft _7628_ (
    .a(_3005_),
    .b(_3006_),
    .y(_3007_)
  );
  al_or3 _7629_ (
    .a(_2998_),
    .b(_2999_),
    .c(_3007_),
    .y(_3008_)
  );
  al_oa21 _7630_ (
    .a(_2998_),
    .b(_2999_),
    .c(_3007_),
    .y(_3009_)
  );
  al_nand2ft _7631_ (
    .a(_3009_),
    .b(_3008_),
    .y(_3010_)
  );
  al_or3fft _7632_ (
    .a(\DFF_158.Q ),
    .b(_0113_),
    .c(_3010_),
    .y(_3011_)
  );
  al_aoi21ftf _7633_ (
    .a(_2991_),
    .b(_0113_),
    .c(_3010_),
    .y(_3012_)
  );
  al_nand2ft _7634_ (
    .a(_3012_),
    .b(_3011_),
    .y(\DFF_1635.D )
  );
  al_or2 _7635_ (
    .a(\DFF_2.Q ),
    .b(g51),
    .y(\DFF_3.D )
  );
  al_or2 _7636_ (
    .a(\DFF_1562.Q ),
    .b(g3234),
    .y(\DFF_1563.D )
  );
  al_nand2 _7637_ (
    .a(\DFF_4.Q ),
    .b(\DFF_3.Q ),
    .y(_3013_)
  );
  al_nor2 _7638_ (
    .a(\DFF_4.Q ),
    .b(\DFF_3.Q ),
    .y(_3014_)
  );
  al_ao21ftf _7639_ (
    .a(_3014_),
    .b(_3013_),
    .c(_0261_),
    .y(\DFF_4.D )
  );
  al_nand2 _7640_ (
    .a(_0326_),
    .b(_0260_),
    .y(_3015_)
  );
  al_ao21ftf _7641_ (
    .a(_0327_),
    .b(_3015_),
    .c(_0329_),
    .y(\DFF_11.D )
  );
  al_ao21 _7642_ (
    .a(\DFF_1563.Q ),
    .b(_0006_),
    .c(\DFF_1607.Q ),
    .y(_3016_)
  );
  al_ao21ftf _7643_ (
    .a(_0334_),
    .b(_3016_),
    .c(_0336_),
    .y(\DFF_1607.D )
  );
  al_nand2 _7644_ (
    .a(_1877_),
    .b(_1912_),
    .y(_3017_)
  );
  al_aoi21ftf _7645_ (
    .a(_1900_),
    .b(\DFF_242.Q ),
    .c(_3017_),
    .y(_3018_)
  );
  al_ao21 _7646_ (
    .a(_1934_),
    .b(_1936_),
    .c(\DFF_237.Q ),
    .y(_3019_)
  );
  al_aoi21ftf _7647_ (
    .a(\DFF_238.Q ),
    .b(_2359_),
    .c(_3019_),
    .y(_3020_)
  );
  al_nand2 _7648_ (
    .a(_1783_),
    .b(_1900_),
    .y(_3021_)
  );
  al_nor3fft _7649_ (
    .a(_0393_),
    .b(_3021_),
    .c(_0274_),
    .y(_3022_)
  );
  al_and3 _7650_ (
    .a(_3020_),
    .b(_3018_),
    .c(_3022_),
    .y(_3023_)
  );
  al_or2 _7651_ (
    .a(_1877_),
    .b(_1912_),
    .y(_3024_)
  );
  al_nand3 _7652_ (
    .a(\DFF_236.Q ),
    .b(_1892_),
    .c(_1894_),
    .y(_3025_)
  );
  al_and3 _7653_ (
    .a(\DFF_245.Q ),
    .b(_1923_),
    .c(_1925_),
    .y(_3026_)
  );
  al_aoi21 _7654_ (
    .a(\DFF_237.Q ),
    .b(_2361_),
    .c(_3026_),
    .y(_3027_)
  );
  al_and3 _7655_ (
    .a(_3025_),
    .b(_3024_),
    .c(_3027_),
    .y(_3028_)
  );
  al_ao21 _7656_ (
    .a(_1885_),
    .b(_1887_),
    .c(\DFF_243.Q ),
    .y(_3029_)
  );
  al_nand3 _7657_ (
    .a(\DFF_243.Q ),
    .b(_1885_),
    .c(_1887_),
    .y(_3030_)
  );
  al_ao21 _7658_ (
    .a(_1892_),
    .b(_1894_),
    .c(\DFF_236.Q ),
    .y(_3031_)
  );
  al_aoi21ftf _7659_ (
    .a(\DFF_245.Q ),
    .b(_2358_),
    .c(_3031_),
    .y(_3032_)
  );
  al_and3 _7660_ (
    .a(_3029_),
    .b(_3030_),
    .c(_3032_),
    .y(_3033_)
  );
  al_and3 _7661_ (
    .a(\DFF_239.Q ),
    .b(_1917_),
    .c(_1919_),
    .y(_3034_)
  );
  al_aoi21 _7662_ (
    .a(_1195_),
    .b(_1931_),
    .c(_3034_),
    .y(_3035_)
  );
  al_aoi21ftf _7663_ (
    .a(_1931_),
    .b(\DFF_240.Q ),
    .c(_3035_),
    .y(_3036_)
  );
  al_and3 _7664_ (
    .a(\DFF_238.Q ),
    .b(_1904_),
    .c(_1906_),
    .y(_3037_)
  );
  al_oa21ttf _7665_ (
    .a(\DFF_241.Q ),
    .b(_1882_),
    .c(_3037_),
    .y(_3038_)
  );
  al_ao21 _7666_ (
    .a(_1917_),
    .b(_1919_),
    .c(\DFF_239.Q ),
    .y(_3039_)
  );
  al_aoi21ttf _7667_ (
    .a(\DFF_241.Q ),
    .b(_1882_),
    .c(_3039_),
    .y(_3040_)
  );
  al_and3 _7668_ (
    .a(_3038_),
    .b(_3040_),
    .c(_3036_),
    .y(_3041_)
  );
  al_and3 _7669_ (
    .a(_3028_),
    .b(_3033_),
    .c(_3041_),
    .y(_3042_)
  );
  al_aoi21 _7670_ (
    .a(_3023_),
    .b(_3042_),
    .c(_2364_),
    .y(\DFF_328.D )
  );
  al_and3fft _7671_ (
    .a(_0287_),
    .b(_2445_),
    .c(_2431_),
    .y(_3043_)
  );
  al_aoi21ttf _7672_ (
    .a(\DFF_587.Q ),
    .b(_2440_),
    .c(_0393_),
    .y(_3044_)
  );
  al_ao21 _7673_ (
    .a(_2006_),
    .b(_2008_),
    .c(\DFF_587.Q ),
    .y(_3045_)
  );
  al_oa21ftt _7674_ (
    .a(\DFF_590.Q ),
    .b(_2433_),
    .c(_3045_),
    .y(_3046_)
  );
  al_ao21 _7675_ (
    .a(_1976_),
    .b(_1978_),
    .c(_0370_),
    .y(_3047_)
  );
  al_and3 _7676_ (
    .a(_0370_),
    .b(_1976_),
    .c(_1978_),
    .y(_3048_)
  );
  al_aoi21ftt _7677_ (
    .a(_3048_),
    .b(_3047_),
    .c(_0288_),
    .y(_3049_)
  );
  al_and3 _7678_ (
    .a(_3044_),
    .b(_3046_),
    .c(_3049_),
    .y(_3050_)
  );
  al_and3 _7679_ (
    .a(\DFF_592.Q ),
    .b(_2031_),
    .c(_2033_),
    .y(_3051_)
  );
  al_aoi21 _7680_ (
    .a(_1804_),
    .b(_2435_),
    .c(_3051_),
    .y(_3052_)
  );
  al_ao21 _7681_ (
    .a(_1988_),
    .b(_1990_),
    .c(\DFF_591.Q ),
    .y(_3053_)
  );
  al_nand3 _7682_ (
    .a(\DFF_593.Q ),
    .b(_1994_),
    .c(_1996_),
    .y(_3054_)
  );
  al_and3 _7683_ (
    .a(_3053_),
    .b(_3054_),
    .c(_3052_),
    .y(_3055_)
  );
  al_ao21 _7684_ (
    .a(_2025_),
    .b(_2027_),
    .c(\DFF_590.Q ),
    .y(_3056_)
  );
  al_nand3 _7685_ (
    .a(\DFF_594.Q ),
    .b(_2019_),
    .c(_2021_),
    .y(_3057_)
  );
  al_nand3 _7686_ (
    .a(\DFF_595.Q ),
    .b(_2013_),
    .c(_2015_),
    .y(_3058_)
  );
  al_aoi21ftf _7687_ (
    .a(\DFF_589.Q ),
    .b(_2439_),
    .c(_3058_),
    .y(_3059_)
  );
  al_and3 _7688_ (
    .a(_3056_),
    .b(_3057_),
    .c(_3059_),
    .y(_3060_)
  );
  al_ao21 _7689_ (
    .a(_2013_),
    .b(_2015_),
    .c(\DFF_595.Q ),
    .y(_3061_)
  );
  al_aoi21ftf _7690_ (
    .a(\DFF_588.Q ),
    .b(_2441_),
    .c(_3061_),
    .y(_3062_)
  );
  al_aoi21ftf _7691_ (
    .a(_2441_),
    .b(\DFF_588.Q ),
    .c(_3062_),
    .y(_3063_)
  );
  al_nand3 _7692_ (
    .a(\DFF_591.Q ),
    .b(_1988_),
    .c(_1990_),
    .y(_3064_)
  );
  al_aoi21ftf _7693_ (
    .a(\DFF_592.Q ),
    .b(_2436_),
    .c(_3064_),
    .y(_3065_)
  );
  al_nand3 _7694_ (
    .a(\DFF_589.Q ),
    .b(_2000_),
    .c(_2002_),
    .y(_3066_)
  );
  al_aoi21ftf _7695_ (
    .a(\DFF_594.Q ),
    .b(_2447_),
    .c(_3066_),
    .y(_3067_)
  );
  al_and3 _7696_ (
    .a(_3065_),
    .b(_3067_),
    .c(_3063_),
    .y(_3068_)
  );
  al_and3 _7697_ (
    .a(_3055_),
    .b(_3060_),
    .c(_3068_),
    .y(_3069_)
  );
  al_aoi21 _7698_ (
    .a(_3050_),
    .b(_3069_),
    .c(_3043_),
    .y(\DFF_678.D )
  );
  al_and3 _7699_ (
    .a(\DFF_942.Q ),
    .b(_2090_),
    .c(_2092_),
    .y(_3070_)
  );
  al_aoi21 _7700_ (
    .a(\DFF_940.Q ),
    .b(_2509_),
    .c(_3070_),
    .y(_3071_)
  );
  al_and3 _7701_ (
    .a(\DFF_939.Q ),
    .b(_2127_),
    .c(_2129_),
    .y(_3072_)
  );
  al_aoi21 _7702_ (
    .a(\DFF_938.Q ),
    .b(_2518_),
    .c(_3072_),
    .y(_3073_)
  );
  al_and3 _7703_ (
    .a(\DFF_936.Q ),
    .b(_2103_),
    .c(_2105_),
    .y(_3074_)
  );
  al_and3fft _7704_ (
    .a(_3074_),
    .b(_0305_),
    .c(_0393_),
    .y(_3075_)
  );
  al_and3 _7705_ (
    .a(_3071_),
    .b(_3073_),
    .c(_3075_),
    .y(_3076_)
  );
  al_ao21 _7706_ (
    .a(_2097_),
    .b(_2099_),
    .c(\DFF_937.Q ),
    .y(_3077_)
  );
  al_and3 _7707_ (
    .a(\DFF_937.Q ),
    .b(_2097_),
    .c(_2099_),
    .y(_3078_)
  );
  al_ao21 _7708_ (
    .a(_2122_),
    .b(_2124_),
    .c(\DFF_941.Q ),
    .y(_3079_)
  );
  al_oa21ftt _7709_ (
    .a(\DFF_944.Q ),
    .b(_2515_),
    .c(_3079_),
    .y(_3080_)
  );
  al_and3ftt _7710_ (
    .a(_3078_),
    .b(_3077_),
    .c(_3080_),
    .y(_3081_)
  );
  al_ao21 _7711_ (
    .a(_2127_),
    .b(_2129_),
    .c(\DFF_939.Q ),
    .y(_3082_)
  );
  al_oa21ftt _7712_ (
    .a(\DFF_945.Q ),
    .b(_2143_),
    .c(_3082_),
    .y(_3083_)
  );
  al_nand3 _7713_ (
    .a(\DFF_941.Q ),
    .b(_2122_),
    .c(_2124_),
    .y(_3084_)
  );
  al_aoi21ftf _7714_ (
    .a(\DFF_944.Q ),
    .b(_2515_),
    .c(_3084_),
    .y(_3085_)
  );
  al_and3 _7715_ (
    .a(_3083_),
    .b(_3085_),
    .c(_3081_),
    .y(_3086_)
  );
  al_ao21 _7716_ (
    .a(_2085_),
    .b(_2087_),
    .c(\DFF_940.Q ),
    .y(_3087_)
  );
  al_aoi21ftf _7717_ (
    .a(\DFF_936.Q ),
    .b(_2511_),
    .c(_3087_),
    .y(_3088_)
  );
  al_aoi21ftf _7718_ (
    .a(\DFF_945.Q ),
    .b(_2143_),
    .c(_3088_),
    .y(_3089_)
  );
  al_ao21 _7719_ (
    .a(_2134_),
    .b(_2136_),
    .c(\DFF_943.Q ),
    .y(_3090_)
  );
  al_nand3 _7720_ (
    .a(\DFF_943.Q ),
    .b(_2134_),
    .c(_2136_),
    .y(_3091_)
  );
  al_ao21 _7721_ (
    .a(_2115_),
    .b(_2117_),
    .c(\DFF_938.Q ),
    .y(_3092_)
  );
  al_aoi21ftf _7722_ (
    .a(\DFF_942.Q ),
    .b(_2510_),
    .c(_3092_),
    .y(_3093_)
  );
  al_and3 _7723_ (
    .a(_3090_),
    .b(_3091_),
    .c(_3093_),
    .y(_3094_)
  );
  al_and3 _7724_ (
    .a(_3089_),
    .b(_3094_),
    .c(_3086_),
    .y(_3095_)
  );
  al_aoi21 _7725_ (
    .a(_3076_),
    .b(_3095_),
    .c(_2526_),
    .y(\DFF_1028.D )
  );
  al_aoi21ftf _7726_ (
    .a(\DFF_1295.Q ),
    .b(_2594_),
    .c(_0393_),
    .y(_3096_)
  );
  al_ao21ttf _7727_ (
    .a(_2193_),
    .b(_2195_),
    .c(\DFF_1292.Q ),
    .y(_3097_)
  );
  al_and3ftt _7728_ (
    .a(\DFF_1292.Q ),
    .b(_2193_),
    .c(_2195_),
    .y(_3098_)
  );
  al_nand2ft _7729_ (
    .a(_3098_),
    .b(_3097_),
    .y(_3099_)
  );
  al_ao21ttf _7730_ (
    .a(_2227_),
    .b(_2229_),
    .c(\DFF_1289.Q ),
    .y(_3100_)
  );
  al_and3ftt _7731_ (
    .a(\DFF_1289.Q ),
    .b(_2227_),
    .c(_2229_),
    .y(_3101_)
  );
  al_aoi21ftf _7732_ (
    .a(_3101_),
    .b(_3100_),
    .c(_3099_),
    .y(_3102_)
  );
  al_and3ftt _7733_ (
    .a(_0321_),
    .b(_3096_),
    .c(_3102_),
    .y(_3103_)
  );
  al_and3 _7734_ (
    .a(\DFF_1295.Q ),
    .b(_2245_),
    .c(_2247_),
    .y(_3104_)
  );
  al_aoi21ftt _7735_ (
    .a(\DFF_1294.Q ),
    .b(_2190_),
    .c(_3104_),
    .y(_3105_)
  );
  al_ao21 _7736_ (
    .a(_2239_),
    .b(_2241_),
    .c(\DFF_1293.Q ),
    .y(_3106_)
  );
  al_nand3 _7737_ (
    .a(\DFF_1288.Q ),
    .b(_2220_),
    .c(_2222_),
    .y(_3107_)
  );
  al_and3 _7738_ (
    .a(_3106_),
    .b(_3107_),
    .c(_3105_),
    .y(_3108_)
  );
  al_and3 _7739_ (
    .a(\DFF_1293.Q ),
    .b(_2239_),
    .c(_2241_),
    .y(_3109_)
  );
  al_oa21ftf _7740_ (
    .a(\DFF_1290.Q ),
    .b(_2217_),
    .c(_3109_),
    .y(_3110_)
  );
  al_and2 _7741_ (
    .a(\DFF_1287.Q ),
    .b(_2204_),
    .y(_3111_)
  );
  al_oa21ttf _7742_ (
    .a(\DFF_1291.Q ),
    .b(_2235_),
    .c(_3111_),
    .y(_3112_)
  );
  al_and3 _7743_ (
    .a(_3110_),
    .b(_3112_),
    .c(_3108_),
    .y(_3113_)
  );
  al_ao21 _7744_ (
    .a(_2220_),
    .b(_2222_),
    .c(\DFF_1288.Q ),
    .y(_3114_)
  );
  al_aoi21ttf _7745_ (
    .a(\DFF_1291.Q ),
    .b(_2235_),
    .c(_3114_),
    .y(_3115_)
  );
  al_aoi21ftf _7746_ (
    .a(_2190_),
    .b(\DFF_1294.Q ),
    .c(_3115_),
    .y(_3116_)
  );
  al_nand2ft _7747_ (
    .a(\DFF_1287.Q ),
    .b(_2202_),
    .y(_3117_)
  );
  al_aoi21ftf _7748_ (
    .a(\DFF_1286.Q ),
    .b(_2209_),
    .c(_3117_),
    .y(_3118_)
  );
  al_nand2ft _7749_ (
    .a(\DFF_1290.Q ),
    .b(_2217_),
    .y(_3119_)
  );
  al_ao21ftf _7750_ (
    .a(_2209_),
    .b(\DFF_1286.Q ),
    .c(_3119_),
    .y(_3120_)
  );
  al_and3ftt _7751_ (
    .a(_3120_),
    .b(_3118_),
    .c(_3116_),
    .y(_3121_)
  );
  al_nand3 _7752_ (
    .a(_3121_),
    .b(_3103_),
    .c(_3113_),
    .y(_3122_)
  );
  al_aoi21ttf _7753_ (
    .a(_0322_),
    .b(_2597_),
    .c(_3122_),
    .y(\DFF_1378.D )
  );
  al_inv _7754_ (
    .a(_0170_),
    .y(\DFF_316.D )
  );
  al_inv _7755_ (
    .a(_0362_),
    .y(\DFF_395.D )
  );
  al_inv _7756_ (
    .a(_0385_),
    .y(\DFF_745.D )
  );
  al_inv _7757_ (
    .a(_0409_),
    .y(\DFF_1095.D )
  );
  al_inv _7758_ (
    .a(_0351_),
    .y(\DFF_362.D )
  );
  al_inv _7759_ (
    .a(_0432_),
    .y(\DFF_1445.D )
  );
  al_inv _7760_ (
    .a(_0375_),
    .y(\DFF_712.D )
  );
  al_inv _7761_ (
    .a(_0399_),
    .y(\DFF_1062.D )
  );
  al_inv _7762_ (
    .a(_0422_),
    .y(\DFF_1412.D )
  );
  al_nand2ft _7763_ (
    .a(\DFF_389.Q ),
    .b(\DFF_1505.Q ),
    .y(_3123_)
  );
  al_aoi21ftf _7764_ (
    .a(\DFF_391.Q ),
    .b(\DFF_1504.Q ),
    .c(_3123_),
    .y(_3124_)
  );
  al_aoi21ftf _7765_ (
    .a(\DFF_390.Q ),
    .b(\DFF_1506.Q ),
    .c(_3124_),
    .y(\DFF_401.D )
  );
  al_nand2ft _7766_ (
    .a(\DFF_739.Q ),
    .b(\DFF_1505.Q ),
    .y(_3125_)
  );
  al_aoi21ftf _7767_ (
    .a(\DFF_741.Q ),
    .b(\DFF_1504.Q ),
    .c(_3125_),
    .y(_3126_)
  );
  al_aoi21ftf _7768_ (
    .a(\DFF_740.Q ),
    .b(\DFF_1506.Q ),
    .c(_3126_),
    .y(\DFF_751.D )
  );
  al_nand2ft _7769_ (
    .a(\DFF_1089.Q ),
    .b(\DFF_1505.Q ),
    .y(_3127_)
  );
  al_aoi21ftf _7770_ (
    .a(\DFF_1091.Q ),
    .b(\DFF_1504.Q ),
    .c(_3127_),
    .y(_3128_)
  );
  al_aoi21ftf _7771_ (
    .a(\DFF_1090.Q ),
    .b(\DFF_1506.Q ),
    .c(_3128_),
    .y(\DFF_1101.D )
  );
  al_nand2ft _7772_ (
    .a(\DFF_1439.Q ),
    .b(\DFF_1505.Q ),
    .y(_3129_)
  );
  al_aoi21ftf _7773_ (
    .a(\DFF_1441.Q ),
    .b(\DFF_1504.Q ),
    .c(_3129_),
    .y(_3130_)
  );
  al_aoi21ftf _7774_ (
    .a(\DFF_1440.Q ),
    .b(\DFF_1506.Q ),
    .c(_3130_),
    .y(\DFF_1451.D )
  );
  al_nand2ft _7775_ (
    .a(\DFF_386.Q ),
    .b(\DFF_1505.Q ),
    .y(_3131_)
  );
  al_aoi21ftf _7776_ (
    .a(\DFF_388.Q ),
    .b(\DFF_1504.Q ),
    .c(_3131_),
    .y(_3132_)
  );
  al_aoi21ftf _7777_ (
    .a(\DFF_387.Q ),
    .b(\DFF_1506.Q ),
    .c(_3132_),
    .y(\DFF_398.D )
  );
  al_nand2ft _7778_ (
    .a(\DFF_736.Q ),
    .b(\DFF_1505.Q ),
    .y(_3133_)
  );
  al_aoi21ftf _7779_ (
    .a(\DFF_738.Q ),
    .b(\DFF_1504.Q ),
    .c(_3133_),
    .y(_3134_)
  );
  al_aoi21ftf _7780_ (
    .a(\DFF_737.Q ),
    .b(\DFF_1506.Q ),
    .c(_3134_),
    .y(\DFF_748.D )
  );
  al_nand2ft _7781_ (
    .a(\DFF_380.Q ),
    .b(\DFF_1505.Q ),
    .y(_3135_)
  );
  al_aoi21ftf _7782_ (
    .a(\DFF_382.Q ),
    .b(\DFF_1504.Q ),
    .c(_3135_),
    .y(_3136_)
  );
  al_aoi21ftf _7783_ (
    .a(\DFF_381.Q ),
    .b(\DFF_1506.Q ),
    .c(_3136_),
    .y(\DFF_403.D )
  );
  al_nand2ft _7784_ (
    .a(\DFF_1086.Q ),
    .b(\DFF_1505.Q ),
    .y(_3137_)
  );
  al_aoi21ftf _7785_ (
    .a(\DFF_1088.Q ),
    .b(\DFF_1504.Q ),
    .c(_3137_),
    .y(_3138_)
  );
  al_aoi21ftf _7786_ (
    .a(\DFF_1087.Q ),
    .b(\DFF_1506.Q ),
    .c(_3138_),
    .y(\DFF_1098.D )
  );
  al_nand2ft _7787_ (
    .a(\DFF_730.Q ),
    .b(\DFF_1505.Q ),
    .y(_3139_)
  );
  al_aoi21ftf _7788_ (
    .a(\DFF_732.Q ),
    .b(\DFF_1504.Q ),
    .c(_3139_),
    .y(_3140_)
  );
  al_aoi21ftf _7789_ (
    .a(\DFF_731.Q ),
    .b(\DFF_1506.Q ),
    .c(_3140_),
    .y(\DFF_753.D )
  );
  al_nand2ft _7790_ (
    .a(\DFF_1436.Q ),
    .b(\DFF_1505.Q ),
    .y(_3141_)
  );
  al_aoi21ftf _7791_ (
    .a(\DFF_1438.Q ),
    .b(\DFF_1504.Q ),
    .c(_3141_),
    .y(_3142_)
  );
  al_aoi21ftf _7792_ (
    .a(\DFF_1437.Q ),
    .b(\DFF_1506.Q ),
    .c(_3142_),
    .y(\DFF_1448.D )
  );
  al_nand2ft _7793_ (
    .a(\DFF_1080.Q ),
    .b(\DFF_1505.Q ),
    .y(_3143_)
  );
  al_aoi21ftf _7794_ (
    .a(\DFF_1082.Q ),
    .b(\DFF_1504.Q ),
    .c(_3143_),
    .y(_3144_)
  );
  al_aoi21ftf _7795_ (
    .a(\DFF_1081.Q ),
    .b(\DFF_1506.Q ),
    .c(_3144_),
    .y(\DFF_1103.D )
  );
  al_nand2ft _7796_ (
    .a(\DFF_1430.Q ),
    .b(\DFF_1505.Q ),
    .y(_3145_)
  );
  al_aoi21ftf _7797_ (
    .a(\DFF_1432.Q ),
    .b(\DFF_1504.Q ),
    .c(_3145_),
    .y(_3146_)
  );
  al_aoi21ftf _7798_ (
    .a(\DFF_1431.Q ),
    .b(\DFF_1506.Q ),
    .c(_3146_),
    .y(\DFF_1453.D )
  );
  al_mux2l _7799_ (
    .a(\DFF_361.Q ),
    .b(\DFF_457.Q ),
    .s(\DFF_1506.Q ),
    .y(\DFF_457.D )
  );
  al_mux2l _7800_ (
    .a(\DFF_711.Q ),
    .b(\DFF_807.Q ),
    .s(\DFF_1506.Q ),
    .y(\DFF_807.D )
  );
  al_mux2l _7801_ (
    .a(\DFF_1061.Q ),
    .b(\DFF_1157.Q ),
    .s(\DFF_1506.Q ),
    .y(\DFF_1157.D )
  );
  al_mux2l _7802_ (
    .a(\DFF_1411.Q ),
    .b(\DFF_1507.Q ),
    .s(\DFF_1506.Q ),
    .y(\DFF_1507.D )
  );
  al_and2ft _7803_ (
    .a(g51),
    .b(\DFF_3.Q ),
    .y(\DFF_1.D )
  );
  al_mux2l _7804_ (
    .a(\DFF_1586.Q ),
    .b(\DFF_1568.Q ),
    .s(\DFF_1613.Q ),
    .y(\DFF_1618.D )
  );
  al_and2ft _7805_ (
    .a(g51),
    .b(\DFF_1.Q ),
    .y(\DFF_2.D )
  );
  al_mux2l _7806_ (
    .a(\DFF_1582.Q ),
    .b(\DFF_1564.Q ),
    .s(\DFF_1613.Q ),
    .y(\DFF_1614.D )
  );
  al_mux2l _7807_ (
    .a(\DFF_1587.Q ),
    .b(\DFF_1569.Q ),
    .s(\DFF_1613.Q ),
    .y(\DFF_1619.D )
  );
  al_mux2l _7808_ (
    .a(\DFF_1583.Q ),
    .b(\DFF_1565.Q ),
    .s(\DFF_1613.Q ),
    .y(\DFF_1615.D )
  );
  al_mux2l _7809_ (
    .a(\DFF_1591.Q ),
    .b(\DFF_1573.Q ),
    .s(\DFF_1613.Q ),
    .y(\DFF_1625.D )
  );
  al_mux2l _7810_ (
    .a(\DFF_1588.Q ),
    .b(\DFF_1570.Q ),
    .s(\DFF_1613.Q ),
    .y(\DFF_1620.D )
  );
  al_mux2l _7811_ (
    .a(\DFF_1584.Q ),
    .b(\DFF_1566.Q ),
    .s(\DFF_1613.Q ),
    .y(\DFF_1616.D )
  );
  al_mux2l _7812_ (
    .a(\DFF_1592.Q ),
    .b(\DFF_1574.Q ),
    .s(\DFF_1613.Q ),
    .y(\DFF_1626.D )
  );
  al_mux2l _7813_ (
    .a(\DFF_1589.Q ),
    .b(\DFF_1571.Q ),
    .s(\DFF_1613.Q ),
    .y(\DFF_1621.D )
  );
  al_mux2l _7814_ (
    .a(\DFF_1585.Q ),
    .b(\DFF_1567.Q ),
    .s(\DFF_1613.Q ),
    .y(\DFF_1617.D )
  );
  al_mux2l _7815_ (
    .a(\DFF_1593.Q ),
    .b(\DFF_1575.Q ),
    .s(\DFF_1613.Q ),
    .y(\DFF_1627.D )
  );
  al_mux2l _7816_ (
    .a(\DFF_1590.Q ),
    .b(\DFF_1572.Q ),
    .s(\DFF_1613.Q ),
    .y(\DFF_1622.D )
  );
  al_mux2l _7817_ (
    .a(\DFF_1594.Q ),
    .b(\DFF_1576.Q ),
    .s(\DFF_1613.Q ),
    .y(\DFF_1628.D )
  );
  al_mux2l _7818_ (
    .a(\DFF_754.Q ),
    .b(\DFF_98.Q ),
    .s(\DFF_1504.Q ),
    .y(\DFF_98.D )
  );
  al_mux2l _7819_ (
    .a(\DFF_1104.Q ),
    .b(\DFF_101.Q ),
    .s(\DFF_1504.Q ),
    .y(\DFF_101.D )
  );
  al_mux2l _7820_ (
    .a(\DFF_754.Q ),
    .b(\DFF_99.Q ),
    .s(\DFF_1505.Q ),
    .y(\DFF_99.D )
  );
  al_mux2l _7821_ (
    .a(\DFF_1454.Q ),
    .b(\DFF_104.Q ),
    .s(\DFF_1504.Q ),
    .y(\DFF_104.D )
  );
  al_mux2l _7822_ (
    .a(\DFF_1104.Q ),
    .b(\DFF_102.Q ),
    .s(\DFF_1505.Q ),
    .y(\DFF_102.D )
  );
  al_mux2l _7823_ (
    .a(\DFF_402.Q ),
    .b(\DFF_119.Q ),
    .s(\DFF_1504.Q ),
    .y(\DFF_119.D )
  );
  al_mux2l _7824_ (
    .a(\DFF_754.Q ),
    .b(\DFF_100.Q ),
    .s(\DFF_1506.Q ),
    .y(\DFF_100.D )
  );
  al_mux2l _7825_ (
    .a(\DFF_1454.Q ),
    .b(\DFF_105.Q ),
    .s(\DFF_1505.Q ),
    .y(\DFF_105.D )
  );
  al_mux2l _7826_ (
    .a(\DFF_752.Q ),
    .b(\DFF_122.Q ),
    .s(\DFF_1504.Q ),
    .y(\DFF_122.D )
  );
  al_mux2l _7827_ (
    .a(\DFF_1104.Q ),
    .b(\DFF_103.Q ),
    .s(\DFF_1506.Q ),
    .y(\DFF_103.D )
  );
  al_mux2l _7828_ (
    .a(\DFF_402.Q ),
    .b(\DFF_120.Q ),
    .s(\DFF_1505.Q ),
    .y(\DFF_120.D )
  );
  al_mux2l _7829_ (
    .a(\DFF_1102.Q ),
    .b(\DFF_125.Q ),
    .s(\DFF_1504.Q ),
    .y(\DFF_125.D )
  );
  al_mux2l _7830_ (
    .a(\DFF_1454.Q ),
    .b(\DFF_106.Q ),
    .s(\DFF_1506.Q ),
    .y(\DFF_106.D )
  );
  al_mux2l _7831_ (
    .a(\DFF_752.Q ),
    .b(\DFF_123.Q ),
    .s(\DFF_1505.Q ),
    .y(\DFF_123.D )
  );
  al_mux2l _7832_ (
    .a(\DFF_1452.Q ),
    .b(\DFF_128.Q ),
    .s(\DFF_1504.Q ),
    .y(\DFF_128.D )
  );
  al_mux2l _7833_ (
    .a(\DFF_402.Q ),
    .b(\DFF_121.Q ),
    .s(\DFF_1506.Q ),
    .y(\DFF_121.D )
  );
  al_mux2l _7834_ (
    .a(\DFF_1102.Q ),
    .b(\DFF_126.Q ),
    .s(\DFF_1505.Q ),
    .y(\DFF_126.D )
  );
  al_mux2l _7835_ (
    .a(\DFF_752.Q ),
    .b(\DFF_124.Q ),
    .s(\DFF_1506.Q ),
    .y(\DFF_124.D )
  );
  al_mux2l _7836_ (
    .a(\DFF_1452.Q ),
    .b(\DFF_129.Q ),
    .s(\DFF_1505.Q ),
    .y(\DFF_129.D )
  );
  al_mux2l _7837_ (
    .a(\DFF_1102.Q ),
    .b(\DFF_127.Q ),
    .s(\DFF_1506.Q ),
    .y(\DFF_127.D )
  );
  al_mux2l _7838_ (
    .a(\DFF_1452.Q ),
    .b(\DFF_130.Q ),
    .s(\DFF_1506.Q ),
    .y(\DFF_130.D )
  );
  al_mux2l _7839_ (
    .a(\DFF_404.Q ),
    .b(\DFF_95.Q ),
    .s(\DFF_1504.Q ),
    .y(\DFF_95.D )
  );
  al_nand2ft _7840_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_360.Q ),
    .y(_3147_)
  );
  al_ao21ftf _7841_ (
    .a(\DFF_359.Q ),
    .b(\DFF_1506.Q ),
    .c(_3147_),
    .y(\DFF_360.D )
  );
  al_nand2ft _7842_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_710.Q ),
    .y(_3148_)
  );
  al_ao21ftf _7843_ (
    .a(\DFF_709.Q ),
    .b(\DFF_1506.Q ),
    .c(_3148_),
    .y(\DFF_710.D )
  );
  al_mux2l _7844_ (
    .a(\DFF_404.Q ),
    .b(\DFF_96.Q ),
    .s(\DFF_1505.Q ),
    .y(\DFF_96.D )
  );
  al_mux2l _7845_ (
    .a(\DFF_360.Q ),
    .b(\DFF_361.Q ),
    .s(\DFF_1506.Q ),
    .y(\DFF_361.D )
  );
  al_nand2ft _7846_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_1060.Q ),
    .y(_3149_)
  );
  al_ao21ftf _7847_ (
    .a(\DFF_1059.Q ),
    .b(\DFF_1506.Q ),
    .c(_3149_),
    .y(\DFF_1060.D )
  );
  al_mux2l _7848_ (
    .a(\DFF_28.Q ),
    .b(\DFF_38.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_38.D )
  );
  al_mux2l _7849_ (
    .a(\DFF_1595.Q ),
    .b(\DFF_1577.Q ),
    .s(\DFF_1613.Q ),
    .y(\DFF_1629.D )
  );
  al_mux2l _7850_ (
    .a(\DFF_710.Q ),
    .b(\DFF_711.Q ),
    .s(\DFF_1506.Q ),
    .y(\DFF_711.D )
  );
  al_nand2ft _7851_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_1410.Q ),
    .y(_3150_)
  );
  al_ao21ftf _7852_ (
    .a(\DFF_1409.Q ),
    .b(\DFF_1506.Q ),
    .c(_3150_),
    .y(\DFF_1410.D )
  );
  al_mux2l _7853_ (
    .a(\DFF_27.Q ),
    .b(\DFF_39.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_39.D )
  );
  al_mux2l _7854_ (
    .a(\DFF_404.Q ),
    .b(\DFF_97.Q ),
    .s(\DFF_1506.Q ),
    .y(\DFF_97.D )
  );
  al_mux2l _7855_ (
    .a(\DFF_1060.Q ),
    .b(\DFF_1061.Q ),
    .s(\DFF_1506.Q ),
    .y(\DFF_1061.D )
  );
  al_mux2l _7856_ (
    .a(\DFF_26.Q ),
    .b(\DFF_40.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_40.D )
  );
  al_mux2l _7857_ (
    .a(\DFF_1596.Q ),
    .b(\DFF_1578.Q ),
    .s(\DFF_1613.Q ),
    .y(\DFF_1630.D )
  );
  al_mux2l _7858_ (
    .a(\DFF_1410.Q ),
    .b(\DFF_1411.Q ),
    .s(\DFF_1506.Q ),
    .y(\DFF_1411.D )
  );
  al_mux2l _7859_ (
    .a(\DFF_25.Q ),
    .b(\DFF_41.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_41.D )
  );
  al_mux2l _7860_ (
    .a(\DFF_24.Q ),
    .b(\DFF_42.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_42.D )
  );
  al_mux2l _7861_ (
    .a(\DFF_31.Q ),
    .b(\DFF_89.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_89.D )
  );
  al_mux2l _7862_ (
    .a(\DFF_1597.Q ),
    .b(\DFF_1579.Q ),
    .s(\DFF_1613.Q ),
    .y(\DFF_1631.D )
  );
  al_mux2l _7863_ (
    .a(\DFF_23.Q ),
    .b(\DFF_43.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_43.D )
  );
  al_mux2l _7864_ (
    .a(\DFF_22.Q ),
    .b(\DFF_44.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_44.D )
  );
  al_mux2l _7865_ (
    .a(\DFF_32.Q ),
    .b(\DFF_88.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_88.D )
  );
  al_mux2l _7866_ (
    .a(\DFF_1598.Q ),
    .b(\DFF_1580.Q ),
    .s(\DFF_1613.Q ),
    .y(\DFF_1632.D )
  );
  al_mux2l _7867_ (
    .a(\DFF_21.Q ),
    .b(\DFF_45.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_45.D )
  );
  al_mux2l _7868_ (
    .a(\DFF_37.Q ),
    .b(\DFF_83.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_83.D )
  );
  al_mux2l _7869_ (
    .a(\DFF_33.Q ),
    .b(\DFF_87.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_87.D )
  );
  al_mux2l _7870_ (
    .a(\DFF_1599.Q ),
    .b(\DFF_1581.Q ),
    .s(\DFF_1613.Q ),
    .y(\DFF_1633.D )
  );
  al_mux2l _7871_ (
    .a(\DFF_34.Q ),
    .b(\DFF_86.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_86.D )
  );
  al_mux2l _7872_ (
    .a(\DFF_30.Q ),
    .b(\DFF_90.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_90.D )
  );
  al_mux2l _7873_ (
    .a(\DFF_35.Q ),
    .b(\DFF_85.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_85.D )
  );
  al_mux2l _7874_ (
    .a(\DFF_36.Q ),
    .b(\DFF_84.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_84.D )
  );
  al_mux2l _7875_ (
    .a(\DFF_71.Q ),
    .b(\DFF_25.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_71.D )
  );
  al_mux2l _7876_ (
    .a(\DFF_73.Q ),
    .b(\DFF_24.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_73.D )
  );
  al_mux2l _7877_ (
    .a(\DFF_65.Q ),
    .b(\DFF_28.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_65.D )
  );
  al_mux2l _7878_ (
    .a(\DFF_47.Q ),
    .b(\DFF_37.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_47.D )
  );
  al_mux2l _7879_ (
    .a(\DFF_75.Q ),
    .b(\DFF_23.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_75.D )
  );
  al_mux2l _7880_ (
    .a(\DFF_67.Q ),
    .b(\DFF_27.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_67.D )
  );
  al_mux2l _7881_ (
    .a(\DFF_49.Q ),
    .b(\DFF_36.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_49.D )
  );
  al_mux2l _7882_ (
    .a(\DFF_77.Q ),
    .b(\DFF_22.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_77.D )
  );
  al_mux2l _7883_ (
    .a(\DFF_69.Q ),
    .b(\DFF_26.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_69.D )
  );
  al_mux2l _7884_ (
    .a(\DFF_51.Q ),
    .b(\DFF_35.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_51.D )
  );
  al_mux2l _7885_ (
    .a(\DFF_79.Q ),
    .b(\DFF_21.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_79.D )
  );
  al_mux2l _7886_ (
    .a(\DFF_53.Q ),
    .b(\DFF_34.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_53.D )
  );
  al_mux2l _7887_ (
    .a(\DFF_55.Q ),
    .b(\DFF_33.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_55.D )
  );
  al_mux2h _7888_ (
    .a(\DFF_458.Q ),
    .b(_0178_),
    .s(\DFF_1506.Q ),
    .y(\DFF_458.D )
  );
  al_mux2h _7889_ (
    .a(\DFF_808.Q ),
    .b(_0178_),
    .s(\DFF_1506.Q ),
    .y(\DFF_808.D )
  );
  al_mux2l _7890_ (
    .a(\DFF_57.Q ),
    .b(\DFF_32.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_57.D )
  );
  al_mux2h _7891_ (
    .a(\DFF_1158.Q ),
    .b(_0178_),
    .s(\DFF_1506.Q ),
    .y(\DFF_1158.D )
  );
  al_mux2h _7892_ (
    .a(\DFF_1508.Q ),
    .b(_0178_),
    .s(\DFF_1506.Q ),
    .y(\DFF_1508.D )
  );
  al_mux2l _7893_ (
    .a(\DFF_59.Q ),
    .b(\DFF_31.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_59.D )
  );
  al_mux2l _7894_ (
    .a(\DFF_61.Q ),
    .b(\DFF_30.Q ),
    .s(\DFF_19.Q ),
    .y(\DFF_61.D )
  );
  al_oai21ftf _7895_ (
    .a(\DFF_1506.Q ),
    .b(\DFF_458.Q ),
    .c(\DFF_459.Q ),
    .y(_3151_)
  );
  al_and3fft _7896_ (
    .a(_0186_),
    .b(_0029_),
    .c(_3151_),
    .y(\DFF_459.D )
  );
  al_mux2l _7897_ (
    .a(\DFF_469.Q ),
    .b(_0010_),
    .s(_0015_),
    .y(\DFF_469.D )
  );
  al_oai21 _7898_ (
    .a(\DFF_15.Q ),
    .b(\DFF_16.Q ),
    .c(_1751_),
    .y(_3152_)
  );
  al_and3fft _7899_ (
    .a(\DFF_1624.Q ),
    .b(\DFF_1634.Q ),
    .c(\DFF_158.Q ),
    .y(_3153_)
  );
  al_or3 _7900_ (
    .a(\DFF_159.Q ),
    .b(\DFF_157.Q ),
    .c(_3153_),
    .y(_3154_)
  );
  al_aoi21ttf _7901_ (
    .a(\DFF_107.Q ),
    .b(_1777_),
    .c(_3154_),
    .y(_3155_)
  );
  al_nand3 _7902_ (
    .a(_1748_),
    .b(_3152_),
    .c(_3155_),
    .y(g25489)
  );
  al_oai21ftf _7903_ (
    .a(_1453_),
    .b(_1761_),
    .c(_2991_),
    .y(_3156_)
  );
  al_and2 _7904_ (
    .a(_1756_),
    .b(_1747_),
    .y(_3157_)
  );
  al_and3ftt _7905_ (
    .a(_1748_),
    .b(\DFF_95.Q ),
    .c(_1747_),
    .y(_3158_)
  );
  al_aoi21 _7906_ (
    .a(\DFF_96.Q ),
    .b(_3157_),
    .c(_3158_),
    .y(_3159_)
  );
  al_oai21 _7907_ (
    .a(\DFF_15.Q ),
    .b(\DFF_16.Q ),
    .c(_1752_),
    .y(_3160_)
  );
  al_aoi21ttf _7908_ (
    .a(\DFF_97.Q ),
    .b(_1755_),
    .c(_3160_),
    .y(_3161_)
  );
  al_and3 _7909_ (
    .a(_3156_),
    .b(_3159_),
    .c(_3161_),
    .y(_3162_)
  );
  al_nand3 _7910_ (
    .a(\DFF_100.Q ),
    .b(_1764_),
    .c(_1747_),
    .y(_3163_)
  );
  al_and2 _7911_ (
    .a(_1773_),
    .b(_1769_),
    .y(_3164_)
  );
  al_and3 _7912_ (
    .a(\DFF_104.Q ),
    .b(_1756_),
    .c(_1769_),
    .y(_3165_)
  );
  al_aoi21 _7913_ (
    .a(\DFF_106.Q ),
    .b(_3164_),
    .c(_3165_),
    .y(_3166_)
  );
  al_nand2 _7914_ (
    .a(\DFF_101.Q ),
    .b(_1767_),
    .y(_3167_)
  );
  al_and3 _7915_ (
    .a(_3163_),
    .b(_3167_),
    .c(_3166_),
    .y(_3168_)
  );
  al_nand3 _7916_ (
    .a(\DFF_105.Q ),
    .b(_1450_),
    .c(_1769_),
    .y(_3169_)
  );
  al_and2 _7917_ (
    .a(_1762_),
    .b(_1747_),
    .y(_3170_)
  );
  al_and3 _7918_ (
    .a(\DFF_98.Q ),
    .b(_1773_),
    .c(_1747_),
    .y(_3171_)
  );
  al_ao21 _7919_ (
    .a(\DFF_99.Q ),
    .b(_3170_),
    .c(_3171_),
    .y(_3172_)
  );
  al_nand3 _7920_ (
    .a(\DFF_102.Q ),
    .b(_1777_),
    .c(_1747_),
    .y(_3173_)
  );
  al_nand3ftt _7921_ (
    .a(_1748_),
    .b(\DFF_103.Q ),
    .c(_1769_),
    .y(_3174_)
  );
  al_nand3 _7922_ (
    .a(_1449_),
    .b(_3173_),
    .c(_3174_),
    .y(_3175_)
  );
  al_nor3ftt _7923_ (
    .a(_3169_),
    .b(_3175_),
    .c(_3172_),
    .y(_3176_)
  );
  al_nand3 _7924_ (
    .a(_3168_),
    .b(_3176_),
    .c(_3162_),
    .y(\DFF_158.D )
  );
  al_and3ftt _7925_ (
    .a(_1748_),
    .b(\DFF_119.Q ),
    .c(_1747_),
    .y(_3177_)
  );
  al_and3 _7926_ (
    .a(\DFF_129.Q ),
    .b(_1450_),
    .c(_1769_),
    .y(_3178_)
  );
  al_and3 _7927_ (
    .a(\DFF_126.Q ),
    .b(_1777_),
    .c(_1747_),
    .y(_3179_)
  );
  al_aoi21 _7928_ (
    .a(\DFF_125.Q ),
    .b(_1767_),
    .c(_3179_),
    .y(_3180_)
  );
  al_nand3fft _7929_ (
    .a(_3177_),
    .b(_3178_),
    .c(_3180_),
    .y(_3181_)
  );
  al_and3 _7930_ (
    .a(\DFF_122.Q ),
    .b(_1773_),
    .c(_1747_),
    .y(_3182_)
  );
  al_and3 _7931_ (
    .a(\DFF_124.Q ),
    .b(_1764_),
    .c(_1747_),
    .y(_3183_)
  );
  al_and3ftt _7932_ (
    .a(_1748_),
    .b(\DFF_127.Q ),
    .c(_1769_),
    .y(_3184_)
  );
  al_aoi21 _7933_ (
    .a(\DFF_130.Q ),
    .b(_3164_),
    .c(_3184_),
    .y(_3185_)
  );
  al_nand3fft _7934_ (
    .a(_3182_),
    .b(_3183_),
    .c(_3185_),
    .y(_3186_)
  );
  al_nand3 _7935_ (
    .a(\DFF_128.Q ),
    .b(_1756_),
    .c(_1769_),
    .y(_3187_)
  );
  al_and3 _7936_ (
    .a(\DFF_121.Q ),
    .b(_1450_),
    .c(_1747_),
    .y(_3188_)
  );
  al_aoi21 _7937_ (
    .a(\DFF_123.Q ),
    .b(_3170_),
    .c(_3188_),
    .y(_3189_)
  );
  al_aoi21ttf _7938_ (
    .a(\DFF_120.Q ),
    .b(_3157_),
    .c(_3189_),
    .y(_3190_)
  );
  al_and2 _7939_ (
    .a(_1762_),
    .b(_1452_),
    .y(_3191_)
  );
  al_nor3fft _7940_ (
    .a(_1449_),
    .b(_1453_),
    .c(_3191_),
    .y(_3192_)
  );
  al_and3 _7941_ (
    .a(_3187_),
    .b(_3192_),
    .c(_3190_),
    .y(_3193_)
  );
  al_nand3fft _7942_ (
    .a(_3181_),
    .b(_3186_),
    .c(_3193_),
    .y(\DFF_156.D )
  );
  al_and3fft _7943_ (
    .a(\DFF_1633.Q ),
    .b(_3009_),
    .c(_3008_),
    .y(_3194_)
  );
  al_oai21ftt _7944_ (
    .a(_3008_),
    .b(_3009_),
    .c(\DFF_1633.Q ),
    .y(_3195_)
  );
  al_and2ft _7945_ (
    .a(_3194_),
    .b(_3195_),
    .y(\DFF_1634.D )
  );
  al_and3fft _7946_ (
    .a(\DFF_1622.Q ),
    .b(_2988_),
    .c(_2987_),
    .y(_3196_)
  );
  al_oai21ftt _7947_ (
    .a(_2987_),
    .b(_2988_),
    .c(\DFF_1622.Q ),
    .y(_3197_)
  );
  al_and2ft _7948_ (
    .a(_3196_),
    .b(_3197_),
    .y(\DFF_1624.D )
  );
  al_and2ft _7949_ (
    .a(\DFF_361.Q ),
    .b(\DFF_360.Q ),
    .y(_3198_)
  );
  al_and2ft _7950_ (
    .a(\DFF_402.Q ),
    .b(\DFF_1504.Q ),
    .y(_3199_)
  );
  al_nor2 _7951_ (
    .a(\DFF_404.Q ),
    .b(g563),
    .y(_3200_)
  );
  al_and3fft _7952_ (
    .a(_3199_),
    .b(\DFF_400.D ),
    .c(_3200_),
    .y(_3201_)
  );
  al_and2ft _7953_ (
    .a(\DFF_506.Q ),
    .b(\DFF_1505.Q ),
    .y(_3202_)
  );
  al_nand2ft _7954_ (
    .a(\DFF_507.Q ),
    .b(\DFF_1506.Q ),
    .y(_3203_)
  );
  al_ao21ftf _7955_ (
    .a(\DFF_505.Q ),
    .b(\DFF_1504.Q ),
    .c(_3203_),
    .y(_3204_)
  );
  al_nor2 _7956_ (
    .a(_0484_),
    .b(_0517_),
    .y(_3205_)
  );
  al_nand3 _7957_ (
    .a(_0480_),
    .b(_0506_),
    .c(_3205_),
    .y(_3206_)
  );
  al_nand2 _7958_ (
    .a(_0494_),
    .b(_0500_),
    .y(_3207_)
  );
  al_nand2ft _7959_ (
    .a(_0527_),
    .b(_0489_),
    .y(_3208_)
  );
  al_nand2ft _7960_ (
    .a(_0474_),
    .b(_0511_),
    .y(_3209_)
  );
  al_nand2ft _7961_ (
    .a(\DFF_508.Q ),
    .b(\DFF_1504.Q ),
    .y(_3210_)
  );
  al_nand2ft _7962_ (
    .a(\DFF_510.Q ),
    .b(\DFF_1506.Q ),
    .y(_3211_)
  );
  al_ao21ftf _7963_ (
    .a(\DFF_509.Q ),
    .b(\DFF_1505.Q ),
    .c(_3211_),
    .y(_3212_)
  );
  al_aoi21ftf _7964_ (
    .a(_3212_),
    .b(_3210_),
    .c(_0468_),
    .y(_3213_)
  );
  al_nor3ftt _7965_ (
    .a(_3213_),
    .b(_3209_),
    .c(_3208_),
    .y(_3214_)
  );
  al_nand3fft _7966_ (
    .a(_3207_),
    .b(_3206_),
    .c(_3214_),
    .y(_3215_)
  );
  al_nand3fft _7967_ (
    .a(_3202_),
    .b(_3204_),
    .c(_3215_),
    .y(_3216_)
  );
  al_nand2 _7968_ (
    .a(\DFF_402.Q ),
    .b(_3216_),
    .y(_3217_)
  );
  al_ao21ttf _7969_ (
    .a(_3201_),
    .b(_3217_),
    .c(_3198_),
    .y(_3218_)
  );
  al_oai21ttf _7970_ (
    .a(\DFF_360.Q ),
    .b(\DFF_443.Q ),
    .c(\DFF_361.Q ),
    .y(_3219_)
  );
  al_and3ftt _7971_ (
    .a(\DFF_399.Q ),
    .b(\DFF_402.Q ),
    .c(_3200_),
    .y(_3220_)
  );
  al_nand2ft _7972_ (
    .a(_0474_),
    .b(_0033_),
    .y(_3221_)
  );
  al_nor2ft _7973_ (
    .a(_0474_),
    .b(_0033_),
    .y(_3222_)
  );
  al_oa21ftt _7974_ (
    .a(_3221_),
    .b(_3222_),
    .c(_3220_),
    .y(_3223_)
  );
  al_and2ft _7975_ (
    .a(_3219_),
    .b(_3201_),
    .y(_3224_)
  );
  al_oai21ttf _7976_ (
    .a(\DFF_361.Q ),
    .b(\DFF_443.Q ),
    .c(\DFF_360.Q ),
    .y(_3225_)
  );
  al_ao21ftt _7977_ (
    .a(\DFF_446.Q ),
    .b(_3224_),
    .c(_3225_),
    .y(_3226_)
  );
  al_ao21 _7978_ (
    .a(_3219_),
    .b(_3223_),
    .c(_3226_),
    .y(_3227_)
  );
  al_nand2 _7979_ (
    .a(_3227_),
    .b(_3218_),
    .y(\DFF_1566.D )
  );
  al_inv _7980_ (
    .a(\DFF_361.Q ),
    .y(_3228_)
  );
  al_or3fft _7981_ (
    .a(\DFF_360.Q ),
    .b(_3228_),
    .c(_3201_),
    .y(_3229_)
  );
  al_aoi21ttf _7982_ (
    .a(_3198_),
    .b(_3217_),
    .c(_3229_),
    .y(_3230_)
  );
  al_oa21ftt _7983_ (
    .a(_0468_),
    .b(_0033_),
    .c(_3220_),
    .y(_3231_)
  );
  al_ao21ftf _7984_ (
    .a(_0468_),
    .b(_0033_),
    .c(_3231_),
    .y(_3232_)
  );
  al_ao21ftt _7985_ (
    .a(\DFF_444.Q ),
    .b(_3224_),
    .c(_3225_),
    .y(_3233_)
  );
  al_oai21ftf _7986_ (
    .a(_3219_),
    .b(_3232_),
    .c(_3233_),
    .y(_3234_)
  );
  al_nand2 _7987_ (
    .a(_3234_),
    .b(_3230_),
    .y(\DFF_1564.D )
  );
  al_nand2ft _7988_ (
    .a(_0511_),
    .b(_0180_),
    .y(_3235_)
  );
  al_nand2ft _7989_ (
    .a(_0520_),
    .b(_0028_),
    .y(_3236_)
  );
  al_aoi21ttf _7990_ (
    .a(_3236_),
    .b(_3235_),
    .c(_3220_),
    .y(_3237_)
  );
  al_ao21ftt _7991_ (
    .a(\DFF_447.Q ),
    .b(_3224_),
    .c(_3225_),
    .y(_3238_)
  );
  al_ao21 _7992_ (
    .a(_3219_),
    .b(_3237_),
    .c(_3238_),
    .y(_3239_)
  );
  al_nand2 _7993_ (
    .a(_3239_),
    .b(_3230_),
    .y(\DFF_1567.D )
  );
  al_nand3 _7994_ (
    .a(_0033_),
    .b(_0506_),
    .c(_3215_),
    .y(_3240_)
  );
  al_ao21 _7995_ (
    .a(_0506_),
    .b(_3215_),
    .c(_0033_),
    .y(_3241_)
  );
  al_nand3 _7996_ (
    .a(_3220_),
    .b(_3240_),
    .c(_3241_),
    .y(_3242_)
  );
  al_nand3 _7997_ (
    .a(_0033_),
    .b(_0500_),
    .c(_3215_),
    .y(_3243_)
  );
  al_ao21 _7998_ (
    .a(_0500_),
    .b(_3215_),
    .c(_0033_),
    .y(_3244_)
  );
  al_and3 _7999_ (
    .a(_3220_),
    .b(_3243_),
    .c(_3244_),
    .y(_3245_)
  );
  al_aoi21ftt _8000_ (
    .a(\DFF_450.Q ),
    .b(_3224_),
    .c(_3225_),
    .y(_3246_)
  );
  al_ao21ttf _8001_ (
    .a(\DFF_361.Q ),
    .b(_3245_),
    .c(_3246_),
    .y(_3247_)
  );
  al_ao21ttf _8002_ (
    .a(_3198_),
    .b(_3242_),
    .c(_3247_),
    .y(\DFF_1570.D )
  );
  al_ao21 _8003_ (
    .a(_0489_),
    .b(_3215_),
    .c(_0028_),
    .y(_3248_)
  );
  al_nand3 _8004_ (
    .a(_0028_),
    .b(_0489_),
    .c(_3215_),
    .y(_3249_)
  );
  al_nand3 _8005_ (
    .a(_3220_),
    .b(_3249_),
    .c(_3248_),
    .y(_3250_)
  );
  al_aoi21ftf _8006_ (
    .a(_0484_),
    .b(_0180_),
    .c(_3220_),
    .y(_3251_)
  );
  al_aoi21ftf _8007_ (
    .a(_0180_),
    .b(_0484_),
    .c(_3251_),
    .y(_3252_)
  );
  al_ao21ftt _8008_ (
    .a(\DFF_451.Q ),
    .b(_3224_),
    .c(_3225_),
    .y(_3253_)
  );
  al_aoi21 _8009_ (
    .a(_3219_),
    .b(_3252_),
    .c(_3253_),
    .y(_3254_)
  );
  al_ao21 _8010_ (
    .a(_3198_),
    .b(_3250_),
    .c(_3254_),
    .y(\DFF_1571.D )
  );
  al_and3fft _8011_ (
    .a(\DFF_448.Q ),
    .b(_3219_),
    .c(_3201_),
    .y(_3255_)
  );
  al_aoi21 _8012_ (
    .a(_0494_),
    .b(_3215_),
    .c(_0033_),
    .y(_3256_)
  );
  al_nand3 _8013_ (
    .a(_0033_),
    .b(_0494_),
    .c(_3215_),
    .y(_3257_)
  );
  al_nor3fft _8014_ (
    .a(_3220_),
    .b(_3257_),
    .c(_3256_),
    .y(_3258_)
  );
  al_ao21 _8015_ (
    .a(\DFF_361.Q ),
    .b(_3258_),
    .c(_3225_),
    .y(_3259_)
  );
  al_aoi21 _8016_ (
    .a(_3229_),
    .b(_3259_),
    .c(_3255_),
    .y(\DFF_1568.D )
  );
  al_or2ft _8017_ (
    .a(_0517_),
    .b(_0180_),
    .y(_3260_)
  );
  al_nand2ft _8018_ (
    .a(_0517_),
    .b(_0180_),
    .y(_3261_)
  );
  al_and3 _8019_ (
    .a(_3220_),
    .b(_3261_),
    .c(_3260_),
    .y(_3262_)
  );
  al_ao21ftt _8020_ (
    .a(\DFF_445.Q ),
    .b(_3224_),
    .c(_3225_),
    .y(_3263_)
  );
  al_ao21 _8021_ (
    .a(\DFF_361.Q ),
    .b(_3262_),
    .c(_3263_),
    .y(_3264_)
  );
  al_nand2 _8022_ (
    .a(_3264_),
    .b(_3218_),
    .y(\DFF_1565.D )
  );
  al_and3fft _8023_ (
    .a(\DFF_449.Q ),
    .b(_3219_),
    .c(_3201_),
    .y(_3265_)
  );
  al_nand3 _8024_ (
    .a(_0028_),
    .b(_0480_),
    .c(_3215_),
    .y(_3266_)
  );
  al_ao21ttf _8025_ (
    .a(_0480_),
    .b(_3215_),
    .c(_0180_),
    .y(_3267_)
  );
  al_and3 _8026_ (
    .a(_3220_),
    .b(_3266_),
    .c(_3267_),
    .y(_3268_)
  );
  al_ao21 _8027_ (
    .a(\DFF_361.Q ),
    .b(_3268_),
    .c(_3225_),
    .y(_3269_)
  );
  al_aoi21 _8028_ (
    .a(_3229_),
    .b(_3269_),
    .c(_3265_),
    .y(\DFF_1569.D )
  );
  al_nand3 _8029_ (
    .a(_3235_),
    .b(_3236_),
    .c(_3223_),
    .y(_3270_)
  );
  al_nand3ftt _8030_ (
    .a(_3222_),
    .b(_3221_),
    .c(_3237_),
    .y(_3271_)
  );
  al_ao21 _8031_ (
    .a(_3271_),
    .b(_3270_),
    .c(_3232_),
    .y(_3272_)
  );
  al_and3 _8032_ (
    .a(_3232_),
    .b(_3271_),
    .c(_3270_),
    .y(_3273_)
  );
  al_nand2ft _8033_ (
    .a(_3273_),
    .b(_3272_),
    .y(_3274_)
  );
  al_nand2 _8034_ (
    .a(_3220_),
    .b(_3257_),
    .y(_3275_)
  );
  al_or3 _8035_ (
    .a(_3256_),
    .b(_3275_),
    .c(_3268_),
    .y(_3276_)
  );
  al_ao21ftf _8036_ (
    .a(_3256_),
    .b(_3257_),
    .c(_3268_),
    .y(_3277_)
  );
  al_ao21ttf _8037_ (
    .a(_3277_),
    .b(_3276_),
    .c(_3274_),
    .y(_3278_)
  );
  al_and3ftt _8038_ (
    .a(_3274_),
    .b(_3277_),
    .c(_3276_),
    .y(_3279_)
  );
  al_nand2ft _8039_ (
    .a(_3279_),
    .b(_3278_),
    .y(_3280_)
  );
  al_nand2ft _8040_ (
    .a(_3252_),
    .b(_3245_),
    .y(_3281_)
  );
  al_ao21ttf _8041_ (
    .a(_3243_),
    .b(_3244_),
    .c(_3252_),
    .y(_3282_)
  );
  al_ao21 _8042_ (
    .a(_3282_),
    .b(_3281_),
    .c(_3262_),
    .y(_3283_)
  );
  al_and3 _8043_ (
    .a(_3262_),
    .b(_3282_),
    .c(_3281_),
    .y(_3284_)
  );
  al_or3ftt _8044_ (
    .a(_3283_),
    .b(_3284_),
    .c(_3280_),
    .y(_3285_)
  );
  al_nand2ft _8045_ (
    .a(_3284_),
    .b(_3283_),
    .y(_3286_)
  );
  al_aoi21 _8046_ (
    .a(_3286_),
    .b(_3280_),
    .c(_3228_),
    .y(_3287_)
  );
  al_mux2l _8047_ (
    .a(\DFF_452.Q ),
    .b(\DFF_453.Q ),
    .s(g3229),
    .y(_3288_)
  );
  al_and3fft _8048_ (
    .a(\DFF_360.Q ),
    .b(\DFF_361.Q ),
    .c(\DFF_443.Q ),
    .y(_3289_)
  );
  al_and3 _8049_ (
    .a(_3288_),
    .b(_3289_),
    .c(_3201_),
    .y(_3290_)
  );
  al_or3fft _8050_ (
    .a(_3240_),
    .b(_3241_),
    .c(_3250_),
    .y(_3291_)
  );
  al_aoi21ttf _8051_ (
    .a(_3242_),
    .b(_3250_),
    .c(\DFF_360.Q ),
    .y(_3292_)
  );
  al_ao21 _8052_ (
    .a(_3291_),
    .b(_3292_),
    .c(_3290_),
    .y(_3293_)
  );
  al_ao21 _8053_ (
    .a(_3285_),
    .b(_3287_),
    .c(_3293_),
    .y(\DFF_1572.D )
  );
  al_inv _8054_ (
    .a(\DFF_711.Q ),
    .y(_3294_)
  );
  al_inv _8055_ (
    .a(\DFF_754.Q ),
    .y(_3295_)
  );
  al_and3fft _8056_ (
    .a(g1249),
    .b(\DFF_750.D ),
    .c(_3295_),
    .y(_3296_)
  );
  al_or3fft _8057_ (
    .a(\DFF_710.Q ),
    .b(_3294_),
    .c(_3296_),
    .y(_3297_)
  );
  al_nand2ft _8058_ (
    .a(\DFF_855.Q ),
    .b(\DFF_1504.Q ),
    .y(_3298_)
  );
  al_aoi21ftf _8059_ (
    .a(\DFF_857.Q ),
    .b(\DFF_1506.Q ),
    .c(_3298_),
    .y(_3299_)
  );
  al_ao21ftf _8060_ (
    .a(\DFF_856.Q ),
    .b(\DFF_1505.Q ),
    .c(_3299_),
    .y(_3300_)
  );
  al_and2ft _8061_ (
    .a(_0564_),
    .b(_0573_),
    .y(_3301_)
  );
  al_nor2 _8062_ (
    .a(_0546_),
    .b(_0590_),
    .y(_3302_)
  );
  al_or2 _8063_ (
    .a(_0552_),
    .b(_0569_),
    .y(_3303_)
  );
  al_and3ftt _8064_ (
    .a(_3303_),
    .b(_3301_),
    .c(_3302_),
    .y(_3304_)
  );
  al_and2ft _8065_ (
    .a(\DFF_859.Q ),
    .b(\DFF_1505.Q ),
    .y(_3305_)
  );
  al_nand2ft _8066_ (
    .a(\DFF_860.Q ),
    .b(\DFF_1506.Q ),
    .y(_3306_)
  );
  al_aoi21ftf _8067_ (
    .a(\DFF_858.Q ),
    .b(\DFF_1504.Q ),
    .c(_3306_),
    .y(_3307_)
  );
  al_aoi21ftt _8068_ (
    .a(_3305_),
    .b(_3307_),
    .c(_0579_),
    .y(_3308_)
  );
  al_and3ftt _8069_ (
    .a(_0605_),
    .b(_0585_),
    .c(_3308_),
    .y(_3309_)
  );
  al_and3 _8070_ (
    .a(_0557_),
    .b(_0596_),
    .c(_3309_),
    .y(_3310_)
  );
  al_ao21 _8071_ (
    .a(_3304_),
    .b(_3310_),
    .c(_3300_),
    .y(_3311_)
  );
  al_and3ftt _8072_ (
    .a(\DFF_711.Q ),
    .b(\DFF_752.Q ),
    .c(\DFF_710.Q ),
    .y(_3312_)
  );
  al_aoi21ttf _8073_ (
    .a(_3312_),
    .b(_3311_),
    .c(_3297_),
    .y(_3313_)
  );
  al_nand2 _8074_ (
    .a(\DFF_752.Q ),
    .b(_3296_),
    .y(_3314_)
  );
  al_nor2ft _8075_ (
    .a(_0569_),
    .b(_0059_),
    .y(_3315_)
  );
  al_nand2ft _8076_ (
    .a(_0569_),
    .b(_0059_),
    .y(_3316_)
  );
  al_nor3ftt _8077_ (
    .a(_3316_),
    .b(_3314_),
    .c(_3315_),
    .y(_3317_)
  );
  al_oa21ttf _8078_ (
    .a(\DFF_710.Q ),
    .b(\DFF_793.Q ),
    .c(\DFF_711.Q ),
    .y(_3318_)
  );
  al_and2 _8079_ (
    .a(_3318_),
    .b(_3296_),
    .y(_3319_)
  );
  al_oai21ttf _8080_ (
    .a(\DFF_711.Q ),
    .b(\DFF_793.Q ),
    .c(\DFF_710.Q ),
    .y(_3320_)
  );
  al_ao21ftt _8081_ (
    .a(\DFF_796.Q ),
    .b(_3319_),
    .c(_3320_),
    .y(_3321_)
  );
  al_ao21 _8082_ (
    .a(\DFF_711.Q ),
    .b(_3317_),
    .c(_3321_),
    .y(_3322_)
  );
  al_nand2 _8083_ (
    .a(_3322_),
    .b(_3313_),
    .y(\DFF_1575.D )
  );
  al_and2ft _8084_ (
    .a(\DFF_711.Q ),
    .b(\DFF_710.Q ),
    .y(_3323_)
  );
  al_ao21ftf _8085_ (
    .a(_3314_),
    .b(_3311_),
    .c(_3323_),
    .y(_3324_)
  );
  al_nor2ft _8086_ (
    .a(_0579_),
    .b(_0059_),
    .y(_3325_)
  );
  al_nand2ft _8087_ (
    .a(_0579_),
    .b(_0059_),
    .y(_3326_)
  );
  al_or3ftt _8088_ (
    .a(_3326_),
    .b(_3314_),
    .c(_3325_),
    .y(_3327_)
  );
  al_ao21ftt _8089_ (
    .a(\DFF_794.Q ),
    .b(_3319_),
    .c(_3320_),
    .y(_3328_)
  );
  al_oai21ftf _8090_ (
    .a(\DFF_711.Q ),
    .b(_3327_),
    .c(_3328_),
    .y(_3329_)
  );
  al_nand2 _8091_ (
    .a(_3329_),
    .b(_3324_),
    .y(\DFF_1573.D )
  );
  al_nand2 _8092_ (
    .a(_0552_),
    .b(_0054_),
    .y(_3330_)
  );
  al_or2 _8093_ (
    .a(_0552_),
    .b(_0054_),
    .y(_3331_)
  );
  al_aoi21 _8094_ (
    .a(_3331_),
    .b(_3330_),
    .c(_3314_),
    .y(_3332_)
  );
  al_aoi21ftt _8095_ (
    .a(\DFF_797.Q ),
    .b(_3319_),
    .c(_3320_),
    .y(_3333_)
  );
  al_ao21ftf _8096_ (
    .a(_3318_),
    .b(_3332_),
    .c(_3333_),
    .y(_3334_)
  );
  al_nand2 _8097_ (
    .a(_3334_),
    .b(_3324_),
    .y(\DFF_1576.D )
  );
  al_nand3fft _8098_ (
    .a(_0564_),
    .b(_0552_),
    .c(_3308_),
    .y(_3335_)
  );
  al_and2ft _8099_ (
    .a(_0590_),
    .b(_0557_),
    .y(_3336_)
  );
  al_nand3fft _8100_ (
    .a(_0546_),
    .b(_0569_),
    .c(_3336_),
    .y(_3337_)
  );
  al_and2ft _8101_ (
    .a(_0605_),
    .b(_0573_),
    .y(_3338_)
  );
  al_and3 _8102_ (
    .a(_0585_),
    .b(_0596_),
    .c(_3338_),
    .y(_3339_)
  );
  al_nand3fft _8103_ (
    .a(_3335_),
    .b(_3337_),
    .c(_3339_),
    .y(_3340_)
  );
  al_nand3fft _8104_ (
    .a(_0059_),
    .b(_0564_),
    .c(_3340_),
    .y(_3341_)
  );
  al_ao21ftf _8105_ (
    .a(_0564_),
    .b(_3340_),
    .c(_0059_),
    .y(_3342_)
  );
  al_nand3ftt _8106_ (
    .a(_3314_),
    .b(_3341_),
    .c(_3342_),
    .y(_3343_)
  );
  al_nand2 _8107_ (
    .a(_3323_),
    .b(_3343_),
    .y(_3344_)
  );
  al_and3 _8108_ (
    .a(_0060_),
    .b(_0596_),
    .c(_3340_),
    .y(_3345_)
  );
  al_ao21ttf _8109_ (
    .a(_3304_),
    .b(_3310_),
    .c(_0596_),
    .y(_3346_)
  );
  al_aoi21 _8110_ (
    .a(_0059_),
    .b(_3346_),
    .c(_3314_),
    .y(_3347_)
  );
  al_nand3fft _8111_ (
    .a(_3294_),
    .b(_3345_),
    .c(_3347_),
    .y(_3348_)
  );
  al_aoi21ftt _8112_ (
    .a(\DFF_800.Q ),
    .b(_3319_),
    .c(_3320_),
    .y(_3349_)
  );
  al_ao21ttf _8113_ (
    .a(_3349_),
    .b(_3348_),
    .c(_3344_),
    .y(\DFF_1579.D )
  );
  al_ao21 _8114_ (
    .a(_0585_),
    .b(_3340_),
    .c(_0055_),
    .y(_3350_)
  );
  al_nand3 _8115_ (
    .a(_0055_),
    .b(_0585_),
    .c(_3340_),
    .y(_3351_)
  );
  al_nand3ftt _8116_ (
    .a(_3314_),
    .b(_3351_),
    .c(_3350_),
    .y(_3352_)
  );
  al_or2ft _8117_ (
    .a(_0590_),
    .b(_0054_),
    .y(_3353_)
  );
  al_and2ft _8118_ (
    .a(_0590_),
    .b(_0054_),
    .y(_3354_)
  );
  al_and3fft _8119_ (
    .a(_3354_),
    .b(_3314_),
    .c(_3353_),
    .y(_3355_)
  );
  al_ao21ftt _8120_ (
    .a(\DFF_801.Q ),
    .b(_3319_),
    .c(_3320_),
    .y(_3356_)
  );
  al_aoi21 _8121_ (
    .a(\DFF_711.Q ),
    .b(_3355_),
    .c(_3356_),
    .y(_3357_)
  );
  al_ao21 _8122_ (
    .a(_3323_),
    .b(_3352_),
    .c(_3357_),
    .y(\DFF_1580.D )
  );
  al_and3ftt _8123_ (
    .a(\DFF_798.Q ),
    .b(_3318_),
    .c(_3296_),
    .y(_3358_)
  );
  al_nand3 _8124_ (
    .a(_0060_),
    .b(_0557_),
    .c(_3340_),
    .y(_3359_)
  );
  al_ao21ttf _8125_ (
    .a(_0557_),
    .b(_3340_),
    .c(_0059_),
    .y(_3360_)
  );
  al_and3ftt _8126_ (
    .a(_3314_),
    .b(_3359_),
    .c(_3360_),
    .y(_3361_)
  );
  al_ao21 _8127_ (
    .a(\DFF_711.Q ),
    .b(_3361_),
    .c(_3320_),
    .y(_3362_)
  );
  al_aoi21 _8128_ (
    .a(_3297_),
    .b(_3362_),
    .c(_3358_),
    .y(\DFF_1577.D )
  );
  al_or2ft _8129_ (
    .a(_0546_),
    .b(_0054_),
    .y(_3363_)
  );
  al_and2ft _8130_ (
    .a(_0546_),
    .b(_0054_),
    .y(_3364_)
  );
  al_and3fft _8131_ (
    .a(_3364_),
    .b(_3314_),
    .c(_3363_),
    .y(_3365_)
  );
  al_ao21ftt _8132_ (
    .a(\DFF_795.Q ),
    .b(_3319_),
    .c(_3320_),
    .y(_3366_)
  );
  al_ao21 _8133_ (
    .a(\DFF_711.Q ),
    .b(_3365_),
    .c(_3366_),
    .y(_3367_)
  );
  al_nand2 _8134_ (
    .a(_3367_),
    .b(_3313_),
    .y(\DFF_1574.D )
  );
  al_and3ftt _8135_ (
    .a(\DFF_799.Q ),
    .b(_3318_),
    .c(_3296_),
    .y(_3368_)
  );
  al_nand3 _8136_ (
    .a(_0055_),
    .b(_0573_),
    .c(_3340_),
    .y(_3369_)
  );
  al_ao21ttf _8137_ (
    .a(_0573_),
    .b(_3340_),
    .c(_0054_),
    .y(_3370_)
  );
  al_and3ftt _8138_ (
    .a(_3314_),
    .b(_3369_),
    .c(_3370_),
    .y(_3371_)
  );
  al_ao21 _8139_ (
    .a(\DFF_711.Q ),
    .b(_3371_),
    .c(_3320_),
    .y(_3372_)
  );
  al_aoi21 _8140_ (
    .a(_3297_),
    .b(_3372_),
    .c(_3368_),
    .y(\DFF_1578.D )
  );
  al_or2ft _8141_ (
    .a(_3316_),
    .b(_3315_),
    .y(_3373_)
  );
  al_mux2l _8142_ (
    .a(_3373_),
    .b(_3317_),
    .s(_3332_),
    .y(_3374_)
  );
  al_nand2ft _8143_ (
    .a(_3354_),
    .b(_3353_),
    .y(_3375_)
  );
  al_nand3ftt _8144_ (
    .a(_3345_),
    .b(_3375_),
    .c(_3347_),
    .y(_3376_)
  );
  al_ao21 _8145_ (
    .a(_0596_),
    .b(_3340_),
    .c(_0060_),
    .y(_3377_)
  );
  al_ao21ftf _8146_ (
    .a(_3345_),
    .b(_3377_),
    .c(_3355_),
    .y(_3378_)
  );
  al_ao21 _8147_ (
    .a(_3378_),
    .b(_3376_),
    .c(_3374_),
    .y(_3379_)
  );
  al_and3 _8148_ (
    .a(_3374_),
    .b(_3378_),
    .c(_3376_),
    .y(_3380_)
  );
  al_nand2ft _8149_ (
    .a(_3380_),
    .b(_3379_),
    .y(_3381_)
  );
  al_ao21ttf _8150_ (
    .a(_3359_),
    .b(_3360_),
    .c(_3371_),
    .y(_3382_)
  );
  al_ao21ttf _8151_ (
    .a(_3369_),
    .b(_3370_),
    .c(_3361_),
    .y(_3383_)
  );
  al_nand2ft _8152_ (
    .a(_3364_),
    .b(_3363_),
    .y(_3384_)
  );
  al_ao21ftf _8153_ (
    .a(_3325_),
    .b(_3326_),
    .c(_3365_),
    .y(_3385_)
  );
  al_aoi21ftf _8154_ (
    .a(_3327_),
    .b(_3384_),
    .c(_3385_),
    .y(_3386_)
  );
  al_ao21 _8155_ (
    .a(_3382_),
    .b(_3383_),
    .c(_3386_),
    .y(_3387_)
  );
  al_nand3 _8156_ (
    .a(_3386_),
    .b(_3382_),
    .c(_3383_),
    .y(_3388_)
  );
  al_ao21 _8157_ (
    .a(_3387_),
    .b(_3388_),
    .c(_3381_),
    .y(_3389_)
  );
  al_nand3 _8158_ (
    .a(_3387_),
    .b(_3388_),
    .c(_3381_),
    .y(_3390_)
  );
  al_nand3 _8159_ (
    .a(\DFF_711.Q ),
    .b(_3390_),
    .c(_3389_),
    .y(_3391_)
  );
  al_mux2l _8160_ (
    .a(\DFF_802.Q ),
    .b(\DFF_803.Q ),
    .s(g3229),
    .y(_3392_)
  );
  al_and3fft _8161_ (
    .a(\DFF_710.Q ),
    .b(\DFF_711.Q ),
    .c(\DFF_793.Q ),
    .y(_3393_)
  );
  al_and3 _8162_ (
    .a(_3392_),
    .b(_3393_),
    .c(_3296_),
    .y(_3394_)
  );
  al_or3fft _8163_ (
    .a(_3341_),
    .b(_3342_),
    .c(_3352_),
    .y(_3395_)
  );
  al_aoi21ttf _8164_ (
    .a(_3352_),
    .b(_3343_),
    .c(\DFF_710.Q ),
    .y(_3396_)
  );
  al_aoi21 _8165_ (
    .a(_3395_),
    .b(_3396_),
    .c(_3394_),
    .y(_3397_)
  );
  al_nand2 _8166_ (
    .a(_3397_),
    .b(_3391_),
    .y(\DFF_1581.D )
  );
  al_inv _8167_ (
    .a(\DFF_1061.Q ),
    .y(_3398_)
  );
  al_and3fft _8168_ (
    .a(\DFF_1104.Q ),
    .b(g1943),
    .c(_1854_),
    .y(_3399_)
  );
  al_or3fft _8169_ (
    .a(\DFF_1060.Q ),
    .b(_3398_),
    .c(_3399_),
    .y(_3400_)
  );
  al_and2ft _8170_ (
    .a(\DFF_1061.Q ),
    .b(\DFF_1060.Q ),
    .y(_3401_)
  );
  al_nand2ft _8171_ (
    .a(\DFF_1205.Q ),
    .b(\DFF_1504.Q ),
    .y(_3402_)
  );
  al_aoi21ftf _8172_ (
    .a(\DFF_1207.Q ),
    .b(\DFF_1506.Q ),
    .c(_3402_),
    .y(_3403_)
  );
  al_aoi21ftf _8173_ (
    .a(\DFF_1206.Q ),
    .b(\DFF_1505.Q ),
    .c(_3403_),
    .y(_3404_)
  );
  al_and2ft _8174_ (
    .a(\DFF_1208.Q ),
    .b(\DFF_1504.Q ),
    .y(_3405_)
  );
  al_nand2ft _8175_ (
    .a(\DFF_1209.Q ),
    .b(\DFF_1505.Q ),
    .y(_3406_)
  );
  al_aoi21ftf _8176_ (
    .a(\DFF_1210.Q ),
    .b(\DFF_1506.Q ),
    .c(_3406_),
    .y(_3407_)
  );
  al_aoi21ftf _8177_ (
    .a(_3405_),
    .b(_3407_),
    .c(_0654_),
    .y(_3408_)
  );
  al_and3ftt _8178_ (
    .a(_0667_),
    .b(_0632_),
    .c(_3408_),
    .y(_3409_)
  );
  al_and2ft _8179_ (
    .a(_0659_),
    .b(_0627_),
    .y(_3410_)
  );
  al_and3 _8180_ (
    .a(_0647_),
    .b(_0637_),
    .c(_3410_),
    .y(_3411_)
  );
  al_and2ft _8181_ (
    .a(_0686_),
    .b(_0678_),
    .y(_3412_)
  );
  al_nand3ftt _8182_ (
    .a(_0644_),
    .b(_0671_),
    .c(_3412_),
    .y(_3413_)
  );
  al_nand3ftt _8183_ (
    .a(_3413_),
    .b(_3409_),
    .c(_3411_),
    .y(_3414_)
  );
  al_nand2 _8184_ (
    .a(_3404_),
    .b(_3414_),
    .y(_3415_)
  );
  al_nand3 _8185_ (
    .a(\DFF_1102.Q ),
    .b(_3401_),
    .c(_3415_),
    .y(_3416_)
  );
  al_and2 _8186_ (
    .a(\DFF_1102.Q ),
    .b(_3399_),
    .y(_3417_)
  );
  al_nand2ft _8187_ (
    .a(_0632_),
    .b(_0086_),
    .y(_3418_)
  );
  al_nor2ft _8188_ (
    .a(_0632_),
    .b(_0086_),
    .y(_3419_)
  );
  al_nand3ftt _8189_ (
    .a(_3419_),
    .b(_3418_),
    .c(_3417_),
    .y(_3420_)
  );
  al_oa21ttf _8190_ (
    .a(\DFF_1060.Q ),
    .b(\DFF_1143.Q ),
    .c(\DFF_1061.Q ),
    .y(_3421_)
  );
  al_and2 _8191_ (
    .a(_3421_),
    .b(_3399_),
    .y(_3422_)
  );
  al_oa21ttf _8192_ (
    .a(\DFF_1061.Q ),
    .b(\DFF_1143.Q ),
    .c(\DFF_1060.Q ),
    .y(_3423_)
  );
  al_aoi21ftf _8193_ (
    .a(\DFF_1146.Q ),
    .b(_3422_),
    .c(_3423_),
    .y(_3424_)
  );
  al_oai21 _8194_ (
    .a(_3398_),
    .b(_3420_),
    .c(_3424_),
    .y(_3425_)
  );
  al_nand3 _8195_ (
    .a(_3400_),
    .b(_3416_),
    .c(_3425_),
    .y(\DFF_1584.D )
  );
  al_aoi21ttf _8196_ (
    .a(_3417_),
    .b(_3415_),
    .c(_3401_),
    .y(_3426_)
  );
  al_or2 _8197_ (
    .a(_0627_),
    .b(_0086_),
    .y(_3427_)
  );
  al_and2ft _8198_ (
    .a(_0625_),
    .b(_0086_),
    .y(_3428_)
  );
  al_nand2ft _8199_ (
    .a(_3428_),
    .b(_3427_),
    .y(_3429_)
  );
  al_and3 _8200_ (
    .a(\DFF_1061.Q ),
    .b(_3429_),
    .c(_3417_),
    .y(_3430_)
  );
  al_aoi21ftf _8201_ (
    .a(\DFF_1144.Q ),
    .b(_3422_),
    .c(_3423_),
    .y(_3431_)
  );
  al_ao21ftt _8202_ (
    .a(_3430_),
    .b(_3431_),
    .c(_3426_),
    .y(\DFF_1582.D )
  );
  al_nand2 _8203_ (
    .a(_0659_),
    .b(_0081_),
    .y(_3432_)
  );
  al_nor2 _8204_ (
    .a(_0659_),
    .b(_0081_),
    .y(_3433_)
  );
  al_nand2ft _8205_ (
    .a(_3433_),
    .b(_3432_),
    .y(_3434_)
  );
  al_and3 _8206_ (
    .a(\DFF_1061.Q ),
    .b(_3434_),
    .c(_3417_),
    .y(_3435_)
  );
  al_aoi21ftf _8207_ (
    .a(\DFF_1147.Q ),
    .b(_3422_),
    .c(_3423_),
    .y(_3436_)
  );
  al_ao21ftt _8208_ (
    .a(_3435_),
    .b(_3436_),
    .c(_3426_),
    .y(\DFF_1585.D )
  );
  al_nand3 _8209_ (
    .a(_0086_),
    .b(_0647_),
    .c(_3414_),
    .y(_3437_)
  );
  al_ao21 _8210_ (
    .a(_0647_),
    .b(_3414_),
    .c(_0086_),
    .y(_3438_)
  );
  al_nand3 _8211_ (
    .a(_3417_),
    .b(_3437_),
    .c(_3438_),
    .y(_3439_)
  );
  al_nand3 _8212_ (
    .a(_0086_),
    .b(_0678_),
    .c(_3414_),
    .y(_3440_)
  );
  al_ao21 _8213_ (
    .a(_0678_),
    .b(_3414_),
    .c(_0086_),
    .y(_3441_)
  );
  al_and3 _8214_ (
    .a(_3417_),
    .b(_3440_),
    .c(_3441_),
    .y(_3442_)
  );
  al_aoi21ftf _8215_ (
    .a(\DFF_1150.Q ),
    .b(_3422_),
    .c(_3423_),
    .y(_3443_)
  );
  al_ao21ftf _8216_ (
    .a(_3421_),
    .b(_3442_),
    .c(_3443_),
    .y(_3444_)
  );
  al_ao21ttf _8217_ (
    .a(_3401_),
    .b(_3439_),
    .c(_3444_),
    .y(\DFF_1588.D )
  );
  al_nand3 _8218_ (
    .a(_0082_),
    .b(_0637_),
    .c(_3414_),
    .y(_3445_)
  );
  al_ao21 _8219_ (
    .a(_0637_),
    .b(_3414_),
    .c(_0082_),
    .y(_3446_)
  );
  al_nand3 _8220_ (
    .a(_3417_),
    .b(_3445_),
    .c(_3446_),
    .y(_3447_)
  );
  al_or2ft _8221_ (
    .a(_0667_),
    .b(_0081_),
    .y(_3448_)
  );
  al_and2ft _8222_ (
    .a(_0667_),
    .b(_0081_),
    .y(_3449_)
  );
  al_nand2ft _8223_ (
    .a(_3449_),
    .b(_3448_),
    .y(_3450_)
  );
  al_nor3fft _8224_ (
    .a(\DFF_1102.Q ),
    .b(_3399_),
    .c(_3450_),
    .y(_3451_)
  );
  al_aoi21ftf _8225_ (
    .a(\DFF_1151.Q ),
    .b(_3422_),
    .c(_3423_),
    .y(_3452_)
  );
  al_aoi21ftf _8226_ (
    .a(_3398_),
    .b(_3451_),
    .c(_3452_),
    .y(_3453_)
  );
  al_ao21 _8227_ (
    .a(_3401_),
    .b(_3447_),
    .c(_3453_),
    .y(\DFF_1589.D )
  );
  al_and3ftt _8228_ (
    .a(\DFF_1148.Q ),
    .b(_3421_),
    .c(_3399_),
    .y(_3454_)
  );
  al_inv _8229_ (
    .a(_0086_),
    .y(_3455_)
  );
  al_and3 _8230_ (
    .a(_3455_),
    .b(_0654_),
    .c(_3414_),
    .y(_3456_)
  );
  al_aoi21 _8231_ (
    .a(_0654_),
    .b(_3414_),
    .c(_3455_),
    .y(_3457_)
  );
  al_oa21 _8232_ (
    .a(_3456_),
    .b(_3457_),
    .c(_3417_),
    .y(_3458_)
  );
  al_ao21ttf _8233_ (
    .a(\DFF_1061.Q ),
    .b(_3458_),
    .c(_3423_),
    .y(_3459_)
  );
  al_aoi21 _8234_ (
    .a(_3400_),
    .b(_3459_),
    .c(_3454_),
    .y(\DFF_1586.D )
  );
  al_or2ft _8235_ (
    .a(_0644_),
    .b(_0081_),
    .y(_3460_)
  );
  al_and2ft _8236_ (
    .a(_0644_),
    .b(_0081_),
    .y(_3461_)
  );
  al_nand2ft _8237_ (
    .a(_3461_),
    .b(_3460_),
    .y(_3462_)
  );
  al_nor3fft _8238_ (
    .a(\DFF_1102.Q ),
    .b(_3399_),
    .c(_3462_),
    .y(_3463_)
  );
  al_ao21ftf _8239_ (
    .a(\DFF_1145.Q ),
    .b(_3422_),
    .c(_3423_),
    .y(_3464_)
  );
  al_ao21ftt _8240_ (
    .a(_3398_),
    .b(_3463_),
    .c(_3464_),
    .y(_3465_)
  );
  al_nand3 _8241_ (
    .a(_3400_),
    .b(_3416_),
    .c(_3465_),
    .y(\DFF_1583.D )
  );
  al_and3ftt _8242_ (
    .a(\DFF_1149.Q ),
    .b(_3421_),
    .c(_3399_),
    .y(_3466_)
  );
  al_nand3 _8243_ (
    .a(_0082_),
    .b(_0671_),
    .c(_3414_),
    .y(_3467_)
  );
  al_ao21ttf _8244_ (
    .a(_0671_),
    .b(_3414_),
    .c(_0081_),
    .y(_3468_)
  );
  al_and3 _8245_ (
    .a(_3417_),
    .b(_3467_),
    .c(_3468_),
    .y(_3469_)
  );
  al_ao21ttf _8246_ (
    .a(\DFF_1061.Q ),
    .b(_3469_),
    .c(_3423_),
    .y(_3470_)
  );
  al_aoi21 _8247_ (
    .a(_3400_),
    .b(_3470_),
    .c(_3466_),
    .y(\DFF_1587.D )
  );
  al_ao21ttf _8248_ (
    .a(_3440_),
    .b(_3441_),
    .c(_3451_),
    .y(_3471_)
  );
  al_nand2 _8249_ (
    .a(_3450_),
    .b(_3442_),
    .y(_3472_)
  );
  al_nand3 _8250_ (
    .a(\DFF_1102.Q ),
    .b(_3434_),
    .c(_3399_),
    .y(_3473_)
  );
  al_mux2l _8251_ (
    .a(_3473_),
    .b(_3434_),
    .s(_3420_),
    .y(_3474_)
  );
  al_and3 _8252_ (
    .a(_3471_),
    .b(_3474_),
    .c(_3472_),
    .y(_3475_)
  );
  al_ao21 _8253_ (
    .a(_3471_),
    .b(_3472_),
    .c(_3474_),
    .y(_3476_)
  );
  al_nand2ft _8254_ (
    .a(_3475_),
    .b(_3476_),
    .y(_3477_)
  );
  al_nand3fft _8255_ (
    .a(_3457_),
    .b(_3456_),
    .c(_3469_),
    .y(_3478_)
  );
  al_ao21ttf _8256_ (
    .a(_3467_),
    .b(_3468_),
    .c(_3458_),
    .y(_3479_)
  );
  al_nand3 _8257_ (
    .a(_3429_),
    .b(_3462_),
    .c(_3417_),
    .y(_3480_)
  );
  al_aoi21ftf _8258_ (
    .a(_3429_),
    .b(_3463_),
    .c(_3480_),
    .y(_3481_)
  );
  al_nand3 _8259_ (
    .a(_3481_),
    .b(_3478_),
    .c(_3479_),
    .y(_3482_)
  );
  al_aoi21 _8260_ (
    .a(_3478_),
    .b(_3479_),
    .c(_3481_),
    .y(_3483_)
  );
  al_or3ftt _8261_ (
    .a(_3482_),
    .b(_3483_),
    .c(_3477_),
    .y(_3484_)
  );
  al_or2ft _8262_ (
    .a(_3482_),
    .b(_3483_),
    .y(_3485_)
  );
  al_aoi21 _8263_ (
    .a(_3477_),
    .b(_3485_),
    .c(_3398_),
    .y(_3486_)
  );
  al_mux2l _8264_ (
    .a(\DFF_1152.Q ),
    .b(\DFF_1153.Q ),
    .s(g3229),
    .y(_3487_)
  );
  al_and3fft _8265_ (
    .a(\DFF_1060.Q ),
    .b(\DFF_1061.Q ),
    .c(\DFF_1143.Q ),
    .y(_3488_)
  );
  al_and3 _8266_ (
    .a(_3487_),
    .b(_3488_),
    .c(_3399_),
    .y(_3489_)
  );
  al_or3fft _8267_ (
    .a(_3445_),
    .b(_3446_),
    .c(_3439_),
    .y(_3490_)
  );
  al_aoi21ttf _8268_ (
    .a(_3439_),
    .b(_3447_),
    .c(\DFF_1060.Q ),
    .y(_3491_)
  );
  al_ao21 _8269_ (
    .a(_3490_),
    .b(_3491_),
    .c(_3489_),
    .y(_3492_)
  );
  al_ao21 _8270_ (
    .a(_3484_),
    .b(_3486_),
    .c(_3492_),
    .y(\DFF_1590.D )
  );
  al_nor2 _8271_ (
    .a(\DFF_1454.Q ),
    .b(g2637),
    .y(_3493_)
  );
  al_and2ft _8272_ (
    .a(\DFF_1411.Q ),
    .b(\DFF_1410.Q ),
    .y(_3494_)
  );
  al_ao21ttf _8273_ (
    .a(_3493_),
    .b(_2334_),
    .c(_3494_),
    .y(_3495_)
  );
  al_nand2ft _8274_ (
    .a(\DFF_1555.Q ),
    .b(\DFF_1504.Q ),
    .y(_3496_)
  );
  al_aoi21ftf _8275_ (
    .a(\DFF_1557.Q ),
    .b(\DFF_1506.Q ),
    .c(_3496_),
    .y(_3497_)
  );
  al_aoi21ftf _8276_ (
    .a(\DFF_1556.Q ),
    .b(\DFF_1505.Q ),
    .c(_3497_),
    .y(_3498_)
  );
  al_aoi21ftf _8277_ (
    .a(_0744_),
    .b(_0746_),
    .c(_0736_),
    .y(_3499_)
  );
  al_and3 _8278_ (
    .a(_0721_),
    .b(_0723_),
    .c(_0740_),
    .y(_3500_)
  );
  al_nand3 _8279_ (
    .a(_0714_),
    .b(_3500_),
    .c(_3499_),
    .y(_3501_)
  );
  al_nand2ft _8280_ (
    .a(\DFF_1560.Q ),
    .b(\DFF_1506.Q ),
    .y(_3502_)
  );
  al_aoi21ftf _8281_ (
    .a(\DFF_1558.Q ),
    .b(\DFF_1504.Q ),
    .c(_3502_),
    .y(_3503_)
  );
  al_ao21ftf _8282_ (
    .a(\DFF_1559.Q ),
    .b(\DFF_1505.Q ),
    .c(_3503_),
    .y(_3504_)
  );
  al_and3 _8283_ (
    .a(_0704_),
    .b(_0706_),
    .c(_3504_),
    .y(_3505_)
  );
  al_nand3ftt _8284_ (
    .a(_0764_),
    .b(_0731_),
    .c(_3505_),
    .y(_3506_)
  );
  al_nor3ftt _8285_ (
    .a(_0753_),
    .b(_0711_),
    .c(_0720_),
    .y(_3507_)
  );
  al_or3ftt _8286_ (
    .a(_3507_),
    .b(_3506_),
    .c(_3501_),
    .y(_3508_)
  );
  al_nand2 _8287_ (
    .a(_3498_),
    .b(_3508_),
    .y(_3509_)
  );
  al_nand3ftt _8288_ (
    .a(\DFF_1411.Q ),
    .b(\DFF_1452.Q ),
    .c(\DFF_1410.Q ),
    .y(_3510_)
  );
  al_ao21ftf _8289_ (
    .a(_3510_),
    .b(_3509_),
    .c(_3495_),
    .y(_3511_)
  );
  al_inv _8290_ (
    .a(\DFF_1411.Q ),
    .y(_3512_)
  );
  al_and3 _8291_ (
    .a(\DFF_1452.Q ),
    .b(_3493_),
    .c(_2334_),
    .y(_3513_)
  );
  al_nand2 _8292_ (
    .a(_0720_),
    .b(_0111_),
    .y(_3514_)
  );
  al_or2 _8293_ (
    .a(_0720_),
    .b(_0111_),
    .y(_3515_)
  );
  al_nand3 _8294_ (
    .a(_3514_),
    .b(_3515_),
    .c(_3513_),
    .y(_3516_)
  );
  al_or2 _8295_ (
    .a(_3512_),
    .b(_3516_),
    .y(_3517_)
  );
  al_and2 _8296_ (
    .a(_3493_),
    .b(_2334_),
    .y(_3518_)
  );
  al_nand2ft _8297_ (
    .a(\DFF_1411.Q ),
    .b(\DFF_1493.Q ),
    .y(_3519_)
  );
  al_aoi21ftf _8298_ (
    .a(_3494_),
    .b(_3519_),
    .c(_3518_),
    .y(_3520_)
  );
  al_oai21ttf _8299_ (
    .a(\DFF_1411.Q ),
    .b(\DFF_1493.Q ),
    .c(\DFF_1410.Q ),
    .y(_3521_)
  );
  al_aoi21ftt _8300_ (
    .a(\DFF_1496.Q ),
    .b(_3520_),
    .c(_3521_),
    .y(_3522_)
  );
  al_ao21 _8301_ (
    .a(_3517_),
    .b(_3522_),
    .c(_3511_),
    .y(\DFF_1593.D )
  );
  al_aoi21ttf _8302_ (
    .a(_3509_),
    .b(_3513_),
    .c(_3494_),
    .y(_3523_)
  );
  al_or2ft _8303_ (
    .a(_0711_),
    .b(_0111_),
    .y(_3524_)
  );
  al_and2ft _8304_ (
    .a(_0711_),
    .b(_0111_),
    .y(_3525_)
  );
  al_nand2ft _8305_ (
    .a(_3525_),
    .b(_3524_),
    .y(_3526_)
  );
  al_nand3 _8306_ (
    .a(\DFF_1411.Q ),
    .b(_3526_),
    .c(_3513_),
    .y(_3527_)
  );
  al_aoi21ftt _8307_ (
    .a(\DFF_1494.Q ),
    .b(_3520_),
    .c(_3521_),
    .y(_3528_)
  );
  al_ao21 _8308_ (
    .a(_3527_),
    .b(_3528_),
    .c(_3523_),
    .y(\DFF_1591.D )
  );
  al_ao21 _8309_ (
    .a(_0704_),
    .b(_0706_),
    .c(_0107_),
    .y(_3529_)
  );
  al_and3 _8310_ (
    .a(_0704_),
    .b(_0706_),
    .c(_0107_),
    .y(_3530_)
  );
  al_nand2ft _8311_ (
    .a(_3530_),
    .b(_3529_),
    .y(_3531_)
  );
  al_nand3 _8312_ (
    .a(\DFF_1411.Q ),
    .b(_3531_),
    .c(_3513_),
    .y(_3532_)
  );
  al_aoi21ftt _8313_ (
    .a(\DFF_1497.Q ),
    .b(_3520_),
    .c(_3521_),
    .y(_3533_)
  );
  al_ao21 _8314_ (
    .a(_3532_),
    .b(_3533_),
    .c(_3523_),
    .y(\DFF_1594.D )
  );
  al_nand2ft _8315_ (
    .a(_0744_),
    .b(_0746_),
    .y(_3534_)
  );
  al_nand3 _8316_ (
    .a(_0111_),
    .b(_3534_),
    .c(_3508_),
    .y(_3535_)
  );
  al_ao21 _8317_ (
    .a(_3534_),
    .b(_3508_),
    .c(_0111_),
    .y(_3536_)
  );
  al_nand3 _8318_ (
    .a(_3535_),
    .b(_3536_),
    .c(_3513_),
    .y(_3537_)
  );
  al_and2 _8319_ (
    .a(_3494_),
    .b(_3537_),
    .y(_3538_)
  );
  al_inv _8320_ (
    .a(_0111_),
    .y(_3539_)
  );
  al_and3 _8321_ (
    .a(_3539_),
    .b(_0740_),
    .c(_3508_),
    .y(_3540_)
  );
  al_ao21 _8322_ (
    .a(_0740_),
    .b(_3508_),
    .c(_3539_),
    .y(_3541_)
  );
  al_nand2ft _8323_ (
    .a(_3540_),
    .b(_3541_),
    .y(_3542_)
  );
  al_nand3 _8324_ (
    .a(\DFF_1411.Q ),
    .b(_3513_),
    .c(_3542_),
    .y(_3543_)
  );
  al_aoi21ftt _8325_ (
    .a(\DFF_1500.Q ),
    .b(_3520_),
    .c(_3521_),
    .y(_3544_)
  );
  al_ao21 _8326_ (
    .a(_3543_),
    .b(_3544_),
    .c(_3538_),
    .y(\DFF_1597.D )
  );
  al_and3 _8327_ (
    .a(_0107_),
    .b(_0731_),
    .c(_3508_),
    .y(_3545_)
  );
  al_ao21 _8328_ (
    .a(_0731_),
    .b(_3508_),
    .c(_0107_),
    .y(_3546_)
  );
  al_nand3ftt _8329_ (
    .a(_3545_),
    .b(_3546_),
    .c(_3513_),
    .y(_3547_)
  );
  al_and2 _8330_ (
    .a(_3494_),
    .b(_3547_),
    .y(_3548_)
  );
  al_and2 _8331_ (
    .a(_0753_),
    .b(_0107_),
    .y(_3549_)
  );
  al_or2 _8332_ (
    .a(_0753_),
    .b(_0107_),
    .y(_3550_)
  );
  al_nand2ft _8333_ (
    .a(_3549_),
    .b(_3550_),
    .y(_3551_)
  );
  al_nand3 _8334_ (
    .a(\DFF_1411.Q ),
    .b(_3551_),
    .c(_3513_),
    .y(_3552_)
  );
  al_aoi21ftt _8335_ (
    .a(\DFF_1501.Q ),
    .b(_3520_),
    .c(_3521_),
    .y(_3553_)
  );
  al_ao21 _8336_ (
    .a(_3552_),
    .b(_3553_),
    .c(_3548_),
    .y(\DFF_1598.D )
  );
  al_and2ft _8337_ (
    .a(\DFF_1498.Q ),
    .b(_3520_),
    .y(_3554_)
  );
  al_and3 _8338_ (
    .a(_3539_),
    .b(_0714_),
    .c(_3508_),
    .y(_3555_)
  );
  al_aoi21 _8339_ (
    .a(_0714_),
    .b(_3508_),
    .c(_3539_),
    .y(_3556_)
  );
  al_oa21 _8340_ (
    .a(_3555_),
    .b(_3556_),
    .c(_3513_),
    .y(_3557_)
  );
  al_ao21 _8341_ (
    .a(\DFF_1411.Q ),
    .b(_3557_),
    .c(_3521_),
    .y(_3558_)
  );
  al_aoi21 _8342_ (
    .a(_3495_),
    .b(_3558_),
    .c(_3554_),
    .y(\DFF_1595.D )
  );
  al_ao21 _8343_ (
    .a(_0721_),
    .b(_0723_),
    .c(_0107_),
    .y(_3559_)
  );
  al_and3 _8344_ (
    .a(_0721_),
    .b(_0723_),
    .c(_0107_),
    .y(_3560_)
  );
  al_nand2ft _8345_ (
    .a(_3560_),
    .b(_3559_),
    .y(_3561_)
  );
  al_nand3 _8346_ (
    .a(\DFF_1411.Q ),
    .b(_3561_),
    .c(_3513_),
    .y(_3562_)
  );
  al_aoi21ftt _8347_ (
    .a(\DFF_1495.Q ),
    .b(_3520_),
    .c(_3521_),
    .y(_3563_)
  );
  al_ao21 _8348_ (
    .a(_3562_),
    .b(_3563_),
    .c(_3511_),
    .y(\DFF_1592.D )
  );
  al_and2ft _8349_ (
    .a(\DFF_1499.Q ),
    .b(_3520_),
    .y(_3564_)
  );
  al_and3 _8350_ (
    .a(_0107_),
    .b(_0736_),
    .c(_3508_),
    .y(_3565_)
  );
  al_ao21 _8351_ (
    .a(_0736_),
    .b(_3508_),
    .c(_0107_),
    .y(_3566_)
  );
  al_and3ftt _8352_ (
    .a(_3565_),
    .b(_3566_),
    .c(_3513_),
    .y(_3567_)
  );
  al_ao21 _8353_ (
    .a(\DFF_1411.Q ),
    .b(_3567_),
    .c(_3521_),
    .y(_3568_)
  );
  al_aoi21 _8354_ (
    .a(_3495_),
    .b(_3568_),
    .c(_3564_),
    .y(\DFF_1596.D )
  );
  al_or3fft _8355_ (
    .a(_3513_),
    .b(_3551_),
    .c(_3542_),
    .y(_3569_)
  );
  al_nand3ftt _8356_ (
    .a(_3551_),
    .b(_3513_),
    .c(_3542_),
    .y(_3570_)
  );
  al_nand3 _8357_ (
    .a(\DFF_1452.Q ),
    .b(_3531_),
    .c(_3518_),
    .y(_3571_)
  );
  al_mux2h _8358_ (
    .a(_3531_),
    .b(_3571_),
    .s(_3516_),
    .y(_3572_)
  );
  al_nand3 _8359_ (
    .a(_3570_),
    .b(_3569_),
    .c(_3572_),
    .y(_3573_)
  );
  al_aoi21 _8360_ (
    .a(_3570_),
    .b(_3569_),
    .c(_3572_),
    .y(_3574_)
  );
  al_nand2ft _8361_ (
    .a(_3574_),
    .b(_3573_),
    .y(_3575_)
  );
  al_nand3fft _8362_ (
    .a(_3555_),
    .b(_3556_),
    .c(_3567_),
    .y(_3576_)
  );
  al_ao21ftf _8363_ (
    .a(_3565_),
    .b(_3566_),
    .c(_3557_),
    .y(_3577_)
  );
  al_and2 _8364_ (
    .a(_3526_),
    .b(_3513_),
    .y(_3578_)
  );
  al_nand3ftt _8365_ (
    .a(_3526_),
    .b(_3561_),
    .c(_3513_),
    .y(_3579_)
  );
  al_aoi21ftf _8366_ (
    .a(_3561_),
    .b(_3578_),
    .c(_3579_),
    .y(_3580_)
  );
  al_ao21 _8367_ (
    .a(_3576_),
    .b(_3577_),
    .c(_3580_),
    .y(_3581_)
  );
  al_and3 _8368_ (
    .a(_3576_),
    .b(_3577_),
    .c(_3580_),
    .y(_3582_)
  );
  al_or3ftt _8369_ (
    .a(_3581_),
    .b(_3582_),
    .c(_3575_),
    .y(_3583_)
  );
  al_or2ft _8370_ (
    .a(_3581_),
    .b(_3582_),
    .y(_3584_)
  );
  al_aoi21 _8371_ (
    .a(_3575_),
    .b(_3584_),
    .c(_3512_),
    .y(_3585_)
  );
  al_mux2l _8372_ (
    .a(\DFF_1502.Q ),
    .b(\DFF_1503.Q ),
    .s(g3229),
    .y(_3586_)
  );
  al_and3fft _8373_ (
    .a(\DFF_1410.Q ),
    .b(_3519_),
    .c(_3586_),
    .y(_3587_)
  );
  al_and3 _8374_ (
    .a(_3493_),
    .b(_3587_),
    .c(_2334_),
    .y(_3588_)
  );
  al_or3fft _8375_ (
    .a(_3535_),
    .b(_3536_),
    .c(_3547_),
    .y(_3589_)
  );
  al_aoi21ttf _8376_ (
    .a(_3547_),
    .b(_3537_),
    .c(\DFF_1410.Q ),
    .y(_3590_)
  );
  al_ao21 _8377_ (
    .a(_3589_),
    .b(_3590_),
    .c(_3588_),
    .y(_3591_)
  );
  al_ao21 _8378_ (
    .a(_3583_),
    .b(_3585_),
    .c(_3591_),
    .y(\DFF_1599.D )
  );
  al_inv _8379_ (
    .a(_1449_),
    .y(\DFF_152.D )
  );
  al_dffl _8380_ (
    .clk(CK),
    .d(\DFF_1.D ),
    .q(\DFF_1.Q )
  );
  al_dffl _8381_ (
    .clk(CK),
    .d(\DFF_2.D ),
    .q(\DFF_2.Q )
  );
  al_dffl _8382_ (
    .clk(CK),
    .d(\DFF_3.D ),
    .q(\DFF_3.Q )
  );
  al_dffl _8383_ (
    .clk(CK),
    .d(\DFF_4.D ),
    .q(\DFF_4.Q )
  );
  al_dffl _8384_ (
    .clk(CK),
    .d(\DFF_5.D ),
    .q(\DFF_5.Q )
  );
  al_dffl _8385_ (
    .clk(CK),
    .d(\DFF_6.D ),
    .q(\DFF_6.Q )
  );
  al_dffl _8386_ (
    .clk(CK),
    .d(\DFF_7.D ),
    .q(\DFF_7.Q )
  );
  al_dffl _8387_ (
    .clk(CK),
    .d(\DFF_8.D ),
    .q(\DFF_8.Q )
  );
  al_dffl _8388_ (
    .clk(CK),
    .d(\DFF_9.D ),
    .q(\DFF_9.Q )
  );
  al_dffl _8389_ (
    .clk(CK),
    .d(\DFF_10.D ),
    .q(\DFF_10.Q )
  );
  al_dffl _8390_ (
    .clk(CK),
    .d(\DFF_11.D ),
    .q(\DFF_11.Q )
  );
  al_dffl _8391_ (
    .clk(CK),
    .d(\DFF_12.D ),
    .q(\DFF_12.Q )
  );
  al_dffl _8392_ (
    .clk(CK),
    .d(\DFF_13.D ),
    .q(\DFF_13.Q )
  );
  al_dffl _8393_ (
    .clk(CK),
    .d(\DFF_14.D ),
    .q(\DFF_14.Q )
  );
  al_dffl _8394_ (
    .clk(CK),
    .d(\DFF_15.D ),
    .q(\DFF_15.Q )
  );
  al_dffl _8395_ (
    .clk(CK),
    .d(\DFF_16.D ),
    .q(\DFF_16.Q )
  );
  al_dffl _8396_ (
    .clk(CK),
    .d(g51),
    .q(\DFF_17.Q )
  );
  al_dffl _8397_ (
    .clk(CK),
    .d(\DFF_17.Q ),
    .q(\DFF_18.Q )
  );
  al_dffl _8398_ (
    .clk(CK),
    .d(\DFF_19.D ),
    .q(\DFF_19.Q )
  );
  al_dffl _8399_ (
    .clk(CK),
    .d(g3212),
    .q(\DFF_20.Q )
  );
  al_dffl _8400_ (
    .clk(CK),
    .d(g3228),
    .q(\DFF_21.Q )
  );
  al_dffl _8401_ (
    .clk(CK),
    .d(g3227),
    .q(\DFF_22.Q )
  );
  al_dffl _8402_ (
    .clk(CK),
    .d(g3226),
    .q(\DFF_23.Q )
  );
  al_dffl _8403_ (
    .clk(CK),
    .d(g3225),
    .q(\DFF_24.Q )
  );
  al_dffl _8404_ (
    .clk(CK),
    .d(g3224),
    .q(\DFF_25.Q )
  );
  al_dffl _8405_ (
    .clk(CK),
    .d(g3223),
    .q(\DFF_26.Q )
  );
  al_dffl _8406_ (
    .clk(CK),
    .d(g3222),
    .q(\DFF_27.Q )
  );
  al_dffl _8407_ (
    .clk(CK),
    .d(g3221),
    .q(\DFF_28.Q )
  );
  al_dffl _8408_ (
    .clk(CK),
    .d(g3232),
    .q(\DFF_29.Q )
  );
  al_dffl _8409_ (
    .clk(CK),
    .d(g3220),
    .q(\DFF_30.Q )
  );
  al_dffl _8410_ (
    .clk(CK),
    .d(g3219),
    .q(\DFF_31.Q )
  );
  al_dffl _8411_ (
    .clk(CK),
    .d(g3218),
    .q(\DFF_32.Q )
  );
  al_dffl _8412_ (
    .clk(CK),
    .d(g3217),
    .q(\DFF_33.Q )
  );
  al_dffl _8413_ (
    .clk(CK),
    .d(g3216),
    .q(\DFF_34.Q )
  );
  al_dffl _8414_ (
    .clk(CK),
    .d(g3215),
    .q(\DFF_35.Q )
  );
  al_dffl _8415_ (
    .clk(CK),
    .d(g3214),
    .q(\DFF_36.Q )
  );
  al_dffl _8416_ (
    .clk(CK),
    .d(g3213),
    .q(\DFF_37.Q )
  );
  al_dffl _8417_ (
    .clk(CK),
    .d(\DFF_38.D ),
    .q(\DFF_38.Q )
  );
  al_dffl _8418_ (
    .clk(CK),
    .d(\DFF_39.D ),
    .q(\DFF_39.Q )
  );
  al_dffl _8419_ (
    .clk(CK),
    .d(\DFF_40.D ),
    .q(\DFF_40.Q )
  );
  al_dffl _8420_ (
    .clk(CK),
    .d(\DFF_41.D ),
    .q(\DFF_41.Q )
  );
  al_dffl _8421_ (
    .clk(CK),
    .d(\DFF_42.D ),
    .q(\DFF_42.Q )
  );
  al_dffl _8422_ (
    .clk(CK),
    .d(\DFF_43.D ),
    .q(\DFF_43.Q )
  );
  al_dffl _8423_ (
    .clk(CK),
    .d(\DFF_44.D ),
    .q(\DFF_44.Q )
  );
  al_dffl _8424_ (
    .clk(CK),
    .d(\DFF_45.D ),
    .q(\DFF_45.Q )
  );
  al_dffl _8425_ (
    .clk(CK),
    .d(\DFF_46.D ),
    .q(\DFF_46.Q )
  );
  al_dffl _8426_ (
    .clk(CK),
    .d(\DFF_47.D ),
    .q(\DFF_47.Q )
  );
  al_dffl _8427_ (
    .clk(CK),
    .d(\DFF_47.Q ),
    .q(\DFF_48.Q )
  );
  al_dffl _8428_ (
    .clk(CK),
    .d(\DFF_49.D ),
    .q(\DFF_49.Q )
  );
  al_dffl _8429_ (
    .clk(CK),
    .d(\DFF_49.Q ),
    .q(\DFF_50.Q )
  );
  al_dffl _8430_ (
    .clk(CK),
    .d(\DFF_51.D ),
    .q(\DFF_51.Q )
  );
  al_dffl _8431_ (
    .clk(CK),
    .d(\DFF_51.Q ),
    .q(\DFF_52.Q )
  );
  al_dffl _8432_ (
    .clk(CK),
    .d(\DFF_53.D ),
    .q(\DFF_53.Q )
  );
  al_dffl _8433_ (
    .clk(CK),
    .d(\DFF_53.Q ),
    .q(\DFF_54.Q )
  );
  al_dffl _8434_ (
    .clk(CK),
    .d(\DFF_55.D ),
    .q(\DFF_55.Q )
  );
  al_dffl _8435_ (
    .clk(CK),
    .d(\DFF_55.Q ),
    .q(\DFF_56.Q )
  );
  al_dffl _8436_ (
    .clk(CK),
    .d(\DFF_57.D ),
    .q(\DFF_57.Q )
  );
  al_dffl _8437_ (
    .clk(CK),
    .d(\DFF_57.Q ),
    .q(\DFF_58.Q )
  );
  al_dffl _8438_ (
    .clk(CK),
    .d(\DFF_59.D ),
    .q(\DFF_59.Q )
  );
  al_dffl _8439_ (
    .clk(CK),
    .d(\DFF_59.Q ),
    .q(\DFF_60.Q )
  );
  al_dffl _8440_ (
    .clk(CK),
    .d(\DFF_61.D ),
    .q(\DFF_61.Q )
  );
  al_dffl _8441_ (
    .clk(CK),
    .d(\DFF_61.Q ),
    .q(\DFF_62.Q )
  );
  al_dffl _8442_ (
    .clk(CK),
    .d(\DFF_63.D ),
    .q(\DFF_63.Q )
  );
  al_dffl _8443_ (
    .clk(CK),
    .d(\DFF_63.Q ),
    .q(\DFF_64.Q )
  );
  al_dffl _8444_ (
    .clk(CK),
    .d(\DFF_65.D ),
    .q(\DFF_65.Q )
  );
  al_dffl _8445_ (
    .clk(CK),
    .d(\DFF_65.Q ),
    .q(\DFF_66.Q )
  );
  al_dffl _8446_ (
    .clk(CK),
    .d(\DFF_67.D ),
    .q(\DFF_67.Q )
  );
  al_dffl _8447_ (
    .clk(CK),
    .d(\DFF_67.Q ),
    .q(\DFF_68.Q )
  );
  al_dffl _8448_ (
    .clk(CK),
    .d(\DFF_69.D ),
    .q(\DFF_69.Q )
  );
  al_dffl _8449_ (
    .clk(CK),
    .d(\DFF_69.Q ),
    .q(\DFF_70.Q )
  );
  al_dffl _8450_ (
    .clk(CK),
    .d(\DFF_71.D ),
    .q(\DFF_71.Q )
  );
  al_dffl _8451_ (
    .clk(CK),
    .d(\DFF_71.Q ),
    .q(\DFF_72.Q )
  );
  al_dffl _8452_ (
    .clk(CK),
    .d(\DFF_73.D ),
    .q(\DFF_73.Q )
  );
  al_dffl _8453_ (
    .clk(CK),
    .d(\DFF_73.Q ),
    .q(\DFF_74.Q )
  );
  al_dffl _8454_ (
    .clk(CK),
    .d(\DFF_75.D ),
    .q(\DFF_75.Q )
  );
  al_dffl _8455_ (
    .clk(CK),
    .d(\DFF_75.Q ),
    .q(\DFF_76.Q )
  );
  al_dffl _8456_ (
    .clk(CK),
    .d(\DFF_77.D ),
    .q(\DFF_77.Q )
  );
  al_dffl _8457_ (
    .clk(CK),
    .d(\DFF_77.Q ),
    .q(\DFF_78.Q )
  );
  al_dffl _8458_ (
    .clk(CK),
    .d(\DFF_79.D ),
    .q(\DFF_79.Q )
  );
  al_dffl _8459_ (
    .clk(CK),
    .d(\DFF_79.Q ),
    .q(\DFF_80.Q )
  );
  al_dffl _8460_ (
    .clk(CK),
    .d(\DFF_81.D ),
    .q(\DFF_81.Q )
  );
  al_dffl _8461_ (
    .clk(CK),
    .d(\DFF_81.Q ),
    .q(\DFF_82.Q )
  );
  al_dffl _8462_ (
    .clk(CK),
    .d(\DFF_83.D ),
    .q(\DFF_83.Q )
  );
  al_dffl _8463_ (
    .clk(CK),
    .d(\DFF_84.D ),
    .q(\DFF_84.Q )
  );
  al_dffl _8464_ (
    .clk(CK),
    .d(\DFF_85.D ),
    .q(\DFF_85.Q )
  );
  al_dffl _8465_ (
    .clk(CK),
    .d(\DFF_86.D ),
    .q(\DFF_86.Q )
  );
  al_dffl _8466_ (
    .clk(CK),
    .d(\DFF_87.D ),
    .q(\DFF_87.Q )
  );
  al_dffl _8467_ (
    .clk(CK),
    .d(\DFF_88.D ),
    .q(\DFF_88.Q )
  );
  al_dffl _8468_ (
    .clk(CK),
    .d(\DFF_89.D ),
    .q(\DFF_89.Q )
  );
  al_dffl _8469_ (
    .clk(CK),
    .d(\DFF_90.D ),
    .q(\DFF_90.Q )
  );
  al_dffl _8470_ (
    .clk(CK),
    .d(\DFF_91.D ),
    .q(\DFF_91.Q )
  );
  al_dffl _8471_ (
    .clk(CK),
    .d(\DFF_95.D ),
    .q(\DFF_95.Q )
  );
  al_dffl _8472_ (
    .clk(CK),
    .d(\DFF_96.D ),
    .q(\DFF_96.Q )
  );
  al_dffl _8473_ (
    .clk(CK),
    .d(\DFF_97.D ),
    .q(\DFF_97.Q )
  );
  al_dffl _8474_ (
    .clk(CK),
    .d(\DFF_98.D ),
    .q(\DFF_98.Q )
  );
  al_dffl _8475_ (
    .clk(CK),
    .d(\DFF_99.D ),
    .q(\DFF_99.Q )
  );
  al_dffl _8476_ (
    .clk(CK),
    .d(\DFF_100.D ),
    .q(\DFF_100.Q )
  );
  al_dffl _8477_ (
    .clk(CK),
    .d(\DFF_101.D ),
    .q(\DFF_101.Q )
  );
  al_dffl _8478_ (
    .clk(CK),
    .d(\DFF_102.D ),
    .q(\DFF_102.Q )
  );
  al_dffl _8479_ (
    .clk(CK),
    .d(\DFF_103.D ),
    .q(\DFF_103.Q )
  );
  al_dffl _8480_ (
    .clk(CK),
    .d(\DFF_104.D ),
    .q(\DFF_104.Q )
  );
  al_dffl _8481_ (
    .clk(CK),
    .d(\DFF_105.D ),
    .q(\DFF_105.Q )
  );
  al_dffl _8482_ (
    .clk(CK),
    .d(\DFF_106.D ),
    .q(\DFF_106.Q )
  );
  al_dffl _8483_ (
    .clk(CK),
    .d(\DFF_107.D ),
    .q(\DFF_107.Q )
  );
  al_dffl _8484_ (
    .clk(CK),
    .d(\DFF_108.D ),
    .q(\DFF_108.Q )
  );
  al_dffl _8485_ (
    .clk(CK),
    .d(\DFF_109.D ),
    .q(\DFF_109.Q )
  );
  al_dffl _8486_ (
    .clk(CK),
    .d(\DFF_110.D ),
    .q(\DFF_110.Q )
  );
  al_dffl _8487_ (
    .clk(CK),
    .d(\DFF_111.D ),
    .q(\DFF_111.Q )
  );
  al_dffl _8488_ (
    .clk(CK),
    .d(\DFF_112.D ),
    .q(\DFF_112.Q )
  );
  al_dffl _8489_ (
    .clk(CK),
    .d(\DFF_113.D ),
    .q(\DFF_113.Q )
  );
  al_dffl _8490_ (
    .clk(CK),
    .d(\DFF_114.D ),
    .q(\DFF_114.Q )
  );
  al_dffl _8491_ (
    .clk(CK),
    .d(\DFF_115.D ),
    .q(\DFF_115.Q )
  );
  al_dffl _8492_ (
    .clk(CK),
    .d(\DFF_116.D ),
    .q(\DFF_116.Q )
  );
  al_dffl _8493_ (
    .clk(CK),
    .d(\DFF_117.D ),
    .q(\DFF_117.Q )
  );
  al_dffl _8494_ (
    .clk(CK),
    .d(\DFF_118.D ),
    .q(\DFF_118.Q )
  );
  al_dffl _8495_ (
    .clk(CK),
    .d(\DFF_119.D ),
    .q(\DFF_119.Q )
  );
  al_dffl _8496_ (
    .clk(CK),
    .d(\DFF_120.D ),
    .q(\DFF_120.Q )
  );
  al_dffl _8497_ (
    .clk(CK),
    .d(\DFF_121.D ),
    .q(\DFF_121.Q )
  );
  al_dffl _8498_ (
    .clk(CK),
    .d(\DFF_122.D ),
    .q(\DFF_122.Q )
  );
  al_dffl _8499_ (
    .clk(CK),
    .d(\DFF_123.D ),
    .q(\DFF_123.Q )
  );
  al_dffl _8500_ (
    .clk(CK),
    .d(\DFF_124.D ),
    .q(\DFF_124.Q )
  );
  al_dffl _8501_ (
    .clk(CK),
    .d(\DFF_125.D ),
    .q(\DFF_125.Q )
  );
  al_dffl _8502_ (
    .clk(CK),
    .d(\DFF_126.D ),
    .q(\DFF_126.Q )
  );
  al_dffl _8503_ (
    .clk(CK),
    .d(\DFF_127.D ),
    .q(\DFF_127.Q )
  );
  al_dffl _8504_ (
    .clk(CK),
    .d(\DFF_128.D ),
    .q(\DFF_128.Q )
  );
  al_dffl _8505_ (
    .clk(CK),
    .d(\DFF_129.D ),
    .q(\DFF_129.Q )
  );
  al_dffl _8506_ (
    .clk(CK),
    .d(\DFF_130.D ),
    .q(\DFF_130.Q )
  );
  al_dffl _8507_ (
    .clk(CK),
    .d(\DFF_131.D ),
    .q(\DFF_131.Q )
  );
  al_dffl _8508_ (
    .clk(CK),
    .d(\DFF_141.D ),
    .q(\DFF_141.Q )
  );
  al_dffl _8509_ (
    .clk(CK),
    .d(\DFF_144.D ),
    .q(\DFF_144.Q )
  );
  al_dffl _8510_ (
    .clk(CK),
    .d(\DFF_146.D ),
    .q(\DFF_146.Q )
  );
  al_dffl _8511_ (
    .clk(CK),
    .d(\DFF_150.D ),
    .q(\DFF_150.Q )
  );
  al_dffl _8512_ (
    .clk(CK),
    .d(\DFF_151.D ),
    .q(\DFF_151.Q )
  );
  al_dffl _8513_ (
    .clk(CK),
    .d(\DFF_152.D ),
    .q(\DFF_152.Q )
  );
  al_dffl _8514_ (
    .clk(CK),
    .d(\DFF_156.D ),
    .q(\DFF_156.Q )
  );
  al_dffl _8515_ (
    .clk(CK),
    .d(\DFF_157.D ),
    .q(\DFF_157.Q )
  );
  al_dffl _8516_ (
    .clk(CK),
    .d(\DFF_158.D ),
    .q(\DFF_158.Q )
  );
  al_dffl _8517_ (
    .clk(CK),
    .d(\DFF_159.D ),
    .q(\DFF_159.Q )
  );
  al_dffl _8518_ (
    .clk(CK),
    .d(\DFF_160.D ),
    .q(\DFF_160.Q )
  );
  al_dffl _8519_ (
    .clk(CK),
    .d(\DFF_164.D ),
    .q(\DFF_164.Q )
  );
  al_dffl _8520_ (
    .clk(CK),
    .d(\DFF_165.D ),
    .q(\DFF_165.Q )
  );
  al_dffl _8521_ (
    .clk(CK),
    .d(\DFF_166.D ),
    .q(\DFF_166.Q )
  );
  al_dffl _8522_ (
    .clk(CK),
    .d(\DFF_167.D ),
    .q(\DFF_167.Q )
  );
  al_dffl _8523_ (
    .clk(CK),
    .d(\DFF_168.D ),
    .q(\DFF_168.Q )
  );
  al_dffl _8524_ (
    .clk(CK),
    .d(\DFF_169.D ),
    .q(\DFF_169.Q )
  );
  al_dffl _8525_ (
    .clk(CK),
    .d(\DFF_170.D ),
    .q(\DFF_170.Q )
  );
  al_dffl _8526_ (
    .clk(CK),
    .d(\DFF_171.D ),
    .q(\DFF_171.Q )
  );
  al_dffl _8527_ (
    .clk(CK),
    .d(\DFF_172.D ),
    .q(\DFF_172.Q )
  );
  al_dffl _8528_ (
    .clk(CK),
    .d(\DFF_173.D ),
    .q(\DFF_173.Q )
  );
  al_dffl _8529_ (
    .clk(CK),
    .d(\DFF_174.D ),
    .q(\DFF_174.Q )
  );
  al_dffl _8530_ (
    .clk(CK),
    .d(\DFF_175.D ),
    .q(\DFF_175.Q )
  );
  al_dffl _8531_ (
    .clk(CK),
    .d(\DFF_176.D ),
    .q(\DFF_176.Q )
  );
  al_dffl _8532_ (
    .clk(CK),
    .d(\DFF_177.D ),
    .q(\DFF_177.Q )
  );
  al_dffl _8533_ (
    .clk(CK),
    .d(\DFF_178.D ),
    .q(\DFF_178.Q )
  );
  al_dffl _8534_ (
    .clk(CK),
    .d(\DFF_179.D ),
    .q(\DFF_179.Q )
  );
  al_dffl _8535_ (
    .clk(CK),
    .d(\DFF_180.D ),
    .q(\DFF_180.Q )
  );
  al_dffl _8536_ (
    .clk(CK),
    .d(\DFF_181.D ),
    .q(\DFF_181.Q )
  );
  al_dffl _8537_ (
    .clk(CK),
    .d(\DFF_182.D ),
    .q(\DFF_182.Q )
  );
  al_dffl _8538_ (
    .clk(CK),
    .d(\DFF_183.D ),
    .q(\DFF_183.Q )
  );
  al_dffl _8539_ (
    .clk(CK),
    .d(\DFF_184.D ),
    .q(\DFF_184.Q )
  );
  al_dffl _8540_ (
    .clk(CK),
    .d(\DFF_185.D ),
    .q(\DFF_185.Q )
  );
  al_dffl _8541_ (
    .clk(CK),
    .d(\DFF_186.D ),
    .q(\DFF_186.Q )
  );
  al_dffl _8542_ (
    .clk(CK),
    .d(\DFF_187.D ),
    .q(\DFF_187.Q )
  );
  al_dffl _8543_ (
    .clk(CK),
    .d(\DFF_188.D ),
    .q(\DFF_188.Q )
  );
  al_dffl _8544_ (
    .clk(CK),
    .d(\DFF_189.D ),
    .q(\DFF_189.Q )
  );
  al_dffl _8545_ (
    .clk(CK),
    .d(\DFF_190.D ),
    .q(\DFF_190.Q )
  );
  al_dffl _8546_ (
    .clk(CK),
    .d(\DFF_191.D ),
    .q(\DFF_191.Q )
  );
  al_dffl _8547_ (
    .clk(CK),
    .d(\DFF_192.D ),
    .q(\DFF_192.Q )
  );
  al_dffl _8548_ (
    .clk(CK),
    .d(\DFF_193.D ),
    .q(\DFF_193.Q )
  );
  al_dffl _8549_ (
    .clk(CK),
    .d(\DFF_194.D ),
    .q(\DFF_194.Q )
  );
  al_dffl _8550_ (
    .clk(CK),
    .d(\DFF_195.D ),
    .q(\DFF_195.Q )
  );
  al_dffl _8551_ (
    .clk(CK),
    .d(\DFF_196.D ),
    .q(\DFF_196.Q )
  );
  al_dffl _8552_ (
    .clk(CK),
    .d(\DFF_197.D ),
    .q(\DFF_197.Q )
  );
  al_dffl _8553_ (
    .clk(CK),
    .d(\DFF_198.D ),
    .q(\DFF_198.Q )
  );
  al_dffl _8554_ (
    .clk(CK),
    .d(\DFF_199.D ),
    .q(\DFF_199.Q )
  );
  al_dffl _8555_ (
    .clk(CK),
    .d(\DFF_200.D ),
    .q(\DFF_200.Q )
  );
  al_dffl _8556_ (
    .clk(CK),
    .d(\DFF_201.D ),
    .q(\DFF_201.Q )
  );
  al_dffl _8557_ (
    .clk(CK),
    .d(\DFF_202.D ),
    .q(\DFF_202.Q )
  );
  al_dffl _8558_ (
    .clk(CK),
    .d(\DFF_203.D ),
    .q(\DFF_203.Q )
  );
  al_dffl _8559_ (
    .clk(CK),
    .d(\DFF_204.D ),
    .q(\DFF_204.Q )
  );
  al_dffl _8560_ (
    .clk(CK),
    .d(\DFF_205.D ),
    .q(\DFF_205.Q )
  );
  al_dffl _8561_ (
    .clk(CK),
    .d(\DFF_206.D ),
    .q(\DFF_206.Q )
  );
  al_dffl _8562_ (
    .clk(CK),
    .d(\DFF_207.D ),
    .q(\DFF_207.Q )
  );
  al_dffl _8563_ (
    .clk(CK),
    .d(\DFF_208.D ),
    .q(\DFF_208.Q )
  );
  al_dffl _8564_ (
    .clk(CK),
    .d(\DFF_209.D ),
    .q(\DFF_209.Q )
  );
  al_dffl _8565_ (
    .clk(CK),
    .d(\DFF_210.D ),
    .q(\DFF_210.Q )
  );
  al_dffl _8566_ (
    .clk(CK),
    .d(\DFF_211.D ),
    .q(\DFF_211.Q )
  );
  al_dffl _8567_ (
    .clk(CK),
    .d(\DFF_212.D ),
    .q(\DFF_212.Q )
  );
  al_dffl _8568_ (
    .clk(CK),
    .d(\DFF_213.D ),
    .q(\DFF_213.Q )
  );
  al_dffl _8569_ (
    .clk(CK),
    .d(\DFF_214.D ),
    .q(\DFF_214.Q )
  );
  al_dffl _8570_ (
    .clk(CK),
    .d(\DFF_215.D ),
    .q(\DFF_215.Q )
  );
  al_dffl _8571_ (
    .clk(CK),
    .d(\DFF_216.D ),
    .q(\DFF_216.Q )
  );
  al_dffl _8572_ (
    .clk(CK),
    .d(\DFF_217.D ),
    .q(\DFF_217.Q )
  );
  al_dffl _8573_ (
    .clk(CK),
    .d(\DFF_218.D ),
    .q(\DFF_218.Q )
  );
  al_dffl _8574_ (
    .clk(CK),
    .d(\DFF_219.D ),
    .q(\DFF_219.Q )
  );
  al_dffl _8575_ (
    .clk(CK),
    .d(\DFF_220.D ),
    .q(\DFF_220.Q )
  );
  al_dffl _8576_ (
    .clk(CK),
    .d(\DFF_221.D ),
    .q(\DFF_221.Q )
  );
  al_dffl _8577_ (
    .clk(CK),
    .d(\DFF_222.D ),
    .q(\DFF_222.Q )
  );
  al_dffl _8578_ (
    .clk(CK),
    .d(\DFF_223.D ),
    .q(\DFF_223.Q )
  );
  al_dffl _8579_ (
    .clk(CK),
    .d(\DFF_224.D ),
    .q(\DFF_224.Q )
  );
  al_dffl _8580_ (
    .clk(CK),
    .d(\DFF_225.D ),
    .q(\DFF_225.Q )
  );
  al_dffl _8581_ (
    .clk(CK),
    .d(\DFF_226.D ),
    .q(\DFF_226.Q )
  );
  al_dffl _8582_ (
    .clk(CK),
    .d(\DFF_227.D ),
    .q(\DFF_227.Q )
  );
  al_dffl _8583_ (
    .clk(CK),
    .d(\DFF_228.D ),
    .q(\DFF_228.Q )
  );
  al_dffl _8584_ (
    .clk(CK),
    .d(\DFF_229.D ),
    .q(\DFF_229.Q )
  );
  al_dffl _8585_ (
    .clk(CK),
    .d(\DFF_230.D ),
    .q(\DFF_230.Q )
  );
  al_dffl _8586_ (
    .clk(CK),
    .d(\DFF_231.D ),
    .q(\DFF_231.Q )
  );
  al_dffl _8587_ (
    .clk(CK),
    .d(\DFF_232.D ),
    .q(\DFF_232.Q )
  );
  al_dffl _8588_ (
    .clk(CK),
    .d(\DFF_233.D ),
    .q(\DFF_233.Q )
  );
  al_dffl _8589_ (
    .clk(CK),
    .d(\DFF_234.D ),
    .q(\DFF_234.Q )
  );
  al_dffl _8590_ (
    .clk(CK),
    .d(\DFF_235.D ),
    .q(\DFF_235.Q )
  );
  al_dffl _8591_ (
    .clk(CK),
    .d(\DFF_236.D ),
    .q(\DFF_236.Q )
  );
  al_dffl _8592_ (
    .clk(CK),
    .d(\DFF_237.D ),
    .q(\DFF_237.Q )
  );
  al_dffl _8593_ (
    .clk(CK),
    .d(\DFF_238.D ),
    .q(\DFF_238.Q )
  );
  al_dffl _8594_ (
    .clk(CK),
    .d(\DFF_239.D ),
    .q(\DFF_239.Q )
  );
  al_dffl _8595_ (
    .clk(CK),
    .d(\DFF_240.D ),
    .q(\DFF_240.Q )
  );
  al_dffl _8596_ (
    .clk(CK),
    .d(\DFF_241.D ),
    .q(\DFF_241.Q )
  );
  al_dffl _8597_ (
    .clk(CK),
    .d(\DFF_242.D ),
    .q(\DFF_242.Q )
  );
  al_dffl _8598_ (
    .clk(CK),
    .d(\DFF_243.D ),
    .q(\DFF_243.Q )
  );
  al_dffl _8599_ (
    .clk(CK),
    .d(\DFF_244.D ),
    .q(\DFF_244.Q )
  );
  al_dffl _8600_ (
    .clk(CK),
    .d(\DFF_245.D ),
    .q(\DFF_245.Q )
  );
  al_dffl _8601_ (
    .clk(CK),
    .d(\DFF_253.D ),
    .q(\DFF_253.Q )
  );
  al_dffl _8602_ (
    .clk(CK),
    .d(\DFF_254.D ),
    .q(\DFF_254.Q )
  );
  al_dffl _8603_ (
    .clk(CK),
    .d(\DFF_255.D ),
    .q(\DFF_255.Q )
  );
  al_dffl _8604_ (
    .clk(CK),
    .d(\DFF_256.D ),
    .q(\DFF_256.Q )
  );
  al_dffl _8605_ (
    .clk(CK),
    .d(\DFF_257.D ),
    .q(\DFF_257.Q )
  );
  al_dffl _8606_ (
    .clk(CK),
    .d(\DFF_258.D ),
    .q(\DFF_258.Q )
  );
  al_dffl _8607_ (
    .clk(CK),
    .d(\DFF_259.D ),
    .q(\DFF_259.Q )
  );
  al_dffl _8608_ (
    .clk(CK),
    .d(\DFF_260.D ),
    .q(\DFF_260.Q )
  );
  al_dffl _8609_ (
    .clk(CK),
    .d(\DFF_261.D ),
    .q(\DFF_261.Q )
  );
  al_dffl _8610_ (
    .clk(CK),
    .d(\DFF_262.D ),
    .q(\DFF_262.Q )
  );
  al_dffl _8611_ (
    .clk(CK),
    .d(\DFF_263.D ),
    .q(\DFF_263.Q )
  );
  al_dffl _8612_ (
    .clk(CK),
    .d(\DFF_264.D ),
    .q(\DFF_264.Q )
  );
  al_dffl _8613_ (
    .clk(CK),
    .d(\DFF_265.D ),
    .q(\DFF_265.Q )
  );
  al_dffl _8614_ (
    .clk(CK),
    .d(\DFF_266.D ),
    .q(\DFF_266.Q )
  );
  al_dffl _8615_ (
    .clk(CK),
    .d(\DFF_267.D ),
    .q(\DFF_267.Q )
  );
  al_dffl _8616_ (
    .clk(CK),
    .d(\DFF_268.D ),
    .q(\DFF_268.Q )
  );
  al_dffl _8617_ (
    .clk(CK),
    .d(\DFF_269.D ),
    .q(\DFF_269.Q )
  );
  al_dffl _8618_ (
    .clk(CK),
    .d(\DFF_270.D ),
    .q(\DFF_270.Q )
  );
  al_dffl _8619_ (
    .clk(CK),
    .d(\DFF_271.D ),
    .q(\DFF_271.Q )
  );
  al_dffl _8620_ (
    .clk(CK),
    .d(\DFF_272.D ),
    .q(\DFF_272.Q )
  );
  al_dffl _8621_ (
    .clk(CK),
    .d(\DFF_273.D ),
    .q(\DFF_273.Q )
  );
  al_dffl _8622_ (
    .clk(CK),
    .d(\DFF_274.D ),
    .q(\DFF_274.Q )
  );
  al_dffl _8623_ (
    .clk(CK),
    .d(\DFF_275.D ),
    .q(\DFF_275.Q )
  );
  al_dffl _8624_ (
    .clk(CK),
    .d(\DFF_276.D ),
    .q(\DFF_276.Q )
  );
  al_dffl _8625_ (
    .clk(CK),
    .d(\DFF_277.D ),
    .q(\DFF_277.Q )
  );
  al_dffl _8626_ (
    .clk(CK),
    .d(\DFF_278.D ),
    .q(\DFF_278.Q )
  );
  al_dffl _8627_ (
    .clk(CK),
    .d(\DFF_279.D ),
    .q(\DFF_279.Q )
  );
  al_dffl _8628_ (
    .clk(CK),
    .d(\DFF_280.D ),
    .q(\DFF_280.Q )
  );
  al_dffl _8629_ (
    .clk(CK),
    .d(\DFF_281.D ),
    .q(\DFF_281.Q )
  );
  al_dffl _8630_ (
    .clk(CK),
    .d(\DFF_282.D ),
    .q(\DFF_282.Q )
  );
  al_dffl _8631_ (
    .clk(CK),
    .d(\DFF_283.D ),
    .q(\DFF_283.Q )
  );
  al_dffl _8632_ (
    .clk(CK),
    .d(\DFF_284.D ),
    .q(\DFF_284.Q )
  );
  al_dffl _8633_ (
    .clk(CK),
    .d(\DFF_285.D ),
    .q(\DFF_285.Q )
  );
  al_dffl _8634_ (
    .clk(CK),
    .d(\DFF_286.D ),
    .q(\DFF_286.Q )
  );
  al_dffl _8635_ (
    .clk(CK),
    .d(\DFF_287.D ),
    .q(\DFF_287.Q )
  );
  al_dffl _8636_ (
    .clk(CK),
    .d(\DFF_288.D ),
    .q(\DFF_288.Q )
  );
  al_dffl _8637_ (
    .clk(CK),
    .d(\DFF_289.D ),
    .q(\DFF_289.Q )
  );
  al_dffl _8638_ (
    .clk(CK),
    .d(\DFF_290.D ),
    .q(\DFF_290.Q )
  );
  al_dffl _8639_ (
    .clk(CK),
    .d(\DFF_291.D ),
    .q(\DFF_291.Q )
  );
  al_dffl _8640_ (
    .clk(CK),
    .d(\DFF_292.D ),
    .q(\DFF_292.Q )
  );
  al_dffl _8641_ (
    .clk(CK),
    .d(\DFF_293.D ),
    .q(\DFF_293.Q )
  );
  al_dffl _8642_ (
    .clk(CK),
    .d(\DFF_294.D ),
    .q(\DFF_294.Q )
  );
  al_dffl _8643_ (
    .clk(CK),
    .d(\DFF_295.D ),
    .q(\DFF_295.Q )
  );
  al_dffl _8644_ (
    .clk(CK),
    .d(\DFF_296.D ),
    .q(\DFF_296.Q )
  );
  al_dffl _8645_ (
    .clk(CK),
    .d(\DFF_297.D ),
    .q(\DFF_297.Q )
  );
  al_dffl _8646_ (
    .clk(CK),
    .d(\DFF_298.D ),
    .q(\DFF_298.Q )
  );
  al_dffl _8647_ (
    .clk(CK),
    .d(\DFF_298.Q ),
    .q(\DFF_299.Q )
  );
  al_dffl _8648_ (
    .clk(CK),
    .d(\DFF_300.D ),
    .q(\DFF_300.Q )
  );
  al_dffl _8649_ (
    .clk(CK),
    .d(\DFF_300.Q ),
    .q(\DFF_301.Q )
  );
  al_dffl _8650_ (
    .clk(CK),
    .d(\DFF_302.D ),
    .q(\DFF_302.Q )
  );
  al_dffl _8651_ (
    .clk(CK),
    .d(\DFF_302.Q ),
    .q(\DFF_303.Q )
  );
  al_dffl _8652_ (
    .clk(CK),
    .d(\DFF_304.D ),
    .q(\DFF_304.Q )
  );
  al_dffl _8653_ (
    .clk(CK),
    .d(\DFF_304.Q ),
    .q(\DFF_305.Q )
  );
  al_dffl _8654_ (
    .clk(CK),
    .d(\DFF_306.D ),
    .q(\DFF_306.Q )
  );
  al_dffl _8655_ (
    .clk(CK),
    .d(\DFF_306.Q ),
    .q(\DFF_307.Q )
  );
  al_dffl _8656_ (
    .clk(CK),
    .d(\DFF_308.D ),
    .q(\DFF_308.Q )
  );
  al_dffl _8657_ (
    .clk(CK),
    .d(\DFF_308.Q ),
    .q(\DFF_309.Q )
  );
  al_dffl _8658_ (
    .clk(CK),
    .d(\DFF_310.D ),
    .q(\DFF_310.Q )
  );
  al_dffl _8659_ (
    .clk(CK),
    .d(\DFF_310.Q ),
    .q(\DFF_311.Q )
  );
  al_dffl _8660_ (
    .clk(CK),
    .d(\DFF_312.D ),
    .q(\DFF_312.Q )
  );
  al_dffl _8661_ (
    .clk(CK),
    .d(\DFF_312.Q ),
    .q(\DFF_313.Q )
  );
  al_dffl _8662_ (
    .clk(CK),
    .d(\DFF_82.Q ),
    .q(\DFF_314.Q )
  );
  al_dffl _8663_ (
    .clk(CK),
    .d(\DFF_314.Q ),
    .q(\DFF_315.Q )
  );
  al_dffl _8664_ (
    .clk(CK),
    .d(\DFF_316.D ),
    .q(\DFF_316.Q )
  );
  al_dffl _8665_ (
    .clk(CK),
    .d(\DFF_317.D ),
    .q(\DFF_317.Q )
  );
  al_dffl _8666_ (
    .clk(CK),
    .d(\DFF_328.D ),
    .q(\DFF_328.Q )
  );
  al_dffl _8667_ (
    .clk(CK),
    .d(\DFF_253.Q ),
    .q(\DFF_329.Q )
  );
  al_dffl _8668_ (
    .clk(CK),
    .d(\DFF_329.Q ),
    .q(\DFF_330.Q )
  );
  al_dffl _8669_ (
    .clk(CK),
    .d(\DFF_254.Q ),
    .q(\DFF_331.Q )
  );
  al_dffl _8670_ (
    .clk(CK),
    .d(\DFF_331.Q ),
    .q(\DFF_332.Q )
  );
  al_dffl _8671_ (
    .clk(CK),
    .d(\DFF_255.Q ),
    .q(\DFF_333.Q )
  );
  al_dffl _8672_ (
    .clk(CK),
    .d(\DFF_333.Q ),
    .q(\DFF_334.Q )
  );
  al_dffl _8673_ (
    .clk(CK),
    .d(\DFF_256.Q ),
    .q(\DFF_335.Q )
  );
  al_dffl _8674_ (
    .clk(CK),
    .d(\DFF_335.Q ),
    .q(\DFF_336.Q )
  );
  al_dffl _8675_ (
    .clk(CK),
    .d(\DFF_257.Q ),
    .q(\DFF_337.Q )
  );
  al_dffl _8676_ (
    .clk(CK),
    .d(\DFF_337.Q ),
    .q(\DFF_338.Q )
  );
  al_dffl _8677_ (
    .clk(CK),
    .d(\DFF_258.Q ),
    .q(\DFF_339.Q )
  );
  al_dffl _8678_ (
    .clk(CK),
    .d(\DFF_339.Q ),
    .q(\DFF_340.Q )
  );
  al_dffl _8679_ (
    .clk(CK),
    .d(\DFF_259.Q ),
    .q(\DFF_341.Q )
  );
  al_dffl _8680_ (
    .clk(CK),
    .d(\DFF_341.Q ),
    .q(\DFF_342.Q )
  );
  al_dffl _8681_ (
    .clk(CK),
    .d(\DFF_260.Q ),
    .q(\DFF_343.Q )
  );
  al_dffl _8682_ (
    .clk(CK),
    .d(\DFF_343.Q ),
    .q(\DFF_344.Q )
  );
  al_dffl _8683_ (
    .clk(CK),
    .d(\DFF_261.Q ),
    .q(\DFF_345.Q )
  );
  al_dffl _8684_ (
    .clk(CK),
    .d(\DFF_345.Q ),
    .q(\DFF_346.Q )
  );
  al_dffl _8685_ (
    .clk(CK),
    .d(\DFF_262.Q ),
    .q(\DFF_347.Q )
  );
  al_dffl _8686_ (
    .clk(CK),
    .d(\DFF_347.Q ),
    .q(\DFF_348.Q )
  );
  al_dffl _8687_ (
    .clk(CK),
    .d(\DFF_263.Q ),
    .q(\DFF_349.Q )
  );
  al_dffl _8688_ (
    .clk(CK),
    .d(\DFF_349.Q ),
    .q(\DFF_350.Q )
  );
  al_dffl _8689_ (
    .clk(CK),
    .d(\DFF_264.Q ),
    .q(\DFF_351.Q )
  );
  al_dffl _8690_ (
    .clk(CK),
    .d(\DFF_351.Q ),
    .q(\DFF_352.Q )
  );
  al_dffl _8691_ (
    .clk(CK),
    .d(\DFF_359.D ),
    .q(\DFF_359.Q )
  );
  al_dffl _8692_ (
    .clk(CK),
    .d(\DFF_360.D ),
    .q(\DFF_360.Q )
  );
  al_dffl _8693_ (
    .clk(CK),
    .d(\DFF_361.D ),
    .q(\DFF_361.Q )
  );
  al_dffl _8694_ (
    .clk(CK),
    .d(\DFF_362.D ),
    .q(\DFF_362.Q )
  );
  al_dffl _8695_ (
    .clk(CK),
    .d(\DFF_362.Q ),
    .q(\DFF_363.Q )
  );
  al_dffl _8696_ (
    .clk(CK),
    .d(\DFF_363.Q ),
    .q(\DFF_364.Q )
  );
  al_dffl _8697_ (
    .clk(CK),
    .d(\DFF_383.Q ),
    .q(\DFF_365.Q )
  );
  al_dffl _8698_ (
    .clk(CK),
    .d(\DFF_365.Q ),
    .q(\DFF_366.Q )
  );
  al_dffl _8699_ (
    .clk(CK),
    .d(\DFF_384.Q ),
    .q(\DFF_367.Q )
  );
  al_dffl _8700_ (
    .clk(CK),
    .d(\DFF_367.Q ),
    .q(\DFF_368.Q )
  );
  al_dffl _8701_ (
    .clk(CK),
    .d(\DFF_385.Q ),
    .q(\DFF_369.Q )
  );
  al_dffl _8702_ (
    .clk(CK),
    .d(\DFF_369.Q ),
    .q(\DFF_370.Q )
  );
  al_dffl _8703_ (
    .clk(CK),
    .d(\DFF_392.Q ),
    .q(\DFF_371.Q )
  );
  al_dffl _8704_ (
    .clk(CK),
    .d(\DFF_371.Q ),
    .q(\DFF_372.Q )
  );
  al_dffl _8705_ (
    .clk(CK),
    .d(\DFF_393.Q ),
    .q(\DFF_373.Q )
  );
  al_dffl _8706_ (
    .clk(CK),
    .d(\DFF_373.Q ),
    .q(\DFF_374.Q )
  );
  al_dffl _8707_ (
    .clk(CK),
    .d(\DFF_394.Q ),
    .q(\DFF_375.Q )
  );
  al_dffl _8708_ (
    .clk(CK),
    .d(\DFF_375.Q ),
    .q(\DFF_376.Q )
  );
  al_dffl _8709_ (
    .clk(CK),
    .d(\DFF_380.D ),
    .q(\DFF_380.Q )
  );
  al_dffl _8710_ (
    .clk(CK),
    .d(\DFF_381.D ),
    .q(\DFF_381.Q )
  );
  al_dffl _8711_ (
    .clk(CK),
    .d(\DFF_382.D ),
    .q(\DFF_382.Q )
  );
  al_dffl _8712_ (
    .clk(CK),
    .d(\DFF_383.D ),
    .q(\DFF_383.Q )
  );
  al_dffl _8713_ (
    .clk(CK),
    .d(\DFF_384.D ),
    .q(\DFF_384.Q )
  );
  al_dffl _8714_ (
    .clk(CK),
    .d(\DFF_385.D ),
    .q(\DFF_385.Q )
  );
  al_dffl _8715_ (
    .clk(CK),
    .d(\DFF_386.D ),
    .q(\DFF_386.Q )
  );
  al_dffl _8716_ (
    .clk(CK),
    .d(\DFF_387.D ),
    .q(\DFF_387.Q )
  );
  al_dffl _8717_ (
    .clk(CK),
    .d(\DFF_388.D ),
    .q(\DFF_388.Q )
  );
  al_dffl _8718_ (
    .clk(CK),
    .d(\DFF_389.D ),
    .q(\DFF_389.Q )
  );
  al_dffl _8719_ (
    .clk(CK),
    .d(\DFF_390.D ),
    .q(\DFF_390.Q )
  );
  al_dffl _8720_ (
    .clk(CK),
    .d(\DFF_391.D ),
    .q(\DFF_391.Q )
  );
  al_dffl _8721_ (
    .clk(CK),
    .d(\DFF_392.D ),
    .q(\DFF_392.Q )
  );
  al_dffl _8722_ (
    .clk(CK),
    .d(\DFF_393.D ),
    .q(\DFF_393.Q )
  );
  al_dffl _8723_ (
    .clk(CK),
    .d(\DFF_394.D ),
    .q(\DFF_394.Q )
  );
  al_dffl _8724_ (
    .clk(CK),
    .d(\DFF_395.D ),
    .q(\DFF_395.Q )
  );
  al_dffl _8725_ (
    .clk(CK),
    .d(\DFF_395.Q ),
    .q(\DFF_396.Q )
  );
  al_dffl _8726_ (
    .clk(CK),
    .d(\DFF_396.Q ),
    .q(\DFF_397.Q )
  );
  al_dffl _8727_ (
    .clk(CK),
    .d(\DFF_398.D ),
    .q(\DFF_398.Q )
  );
  al_dffl _8728_ (
    .clk(CK),
    .d(\DFF_398.Q ),
    .q(\DFF_399.Q )
  );
  al_dffl _8729_ (
    .clk(CK),
    .d(\DFF_400.D ),
    .q(\DFF_400.Q )
  );
  al_dffl _8730_ (
    .clk(CK),
    .d(\DFF_401.D ),
    .q(\DFF_401.Q )
  );
  al_dffl _8731_ (
    .clk(CK),
    .d(\DFF_401.Q ),
    .q(\DFF_402.Q )
  );
  al_dffl _8732_ (
    .clk(CK),
    .d(\DFF_403.D ),
    .q(\DFF_403.Q )
  );
  al_dffl _8733_ (
    .clk(CK),
    .d(\DFF_403.Q ),
    .q(\DFF_404.Q )
  );
  al_dffl _8734_ (
    .clk(CK),
    .d(\DFF_405.D ),
    .q(\DFF_405.Q )
  );
  al_dffl _8735_ (
    .clk(CK),
    .d(\DFF_406.D ),
    .q(\DFF_406.Q )
  );
  al_dffl _8736_ (
    .clk(CK),
    .d(\DFF_407.D ),
    .q(\DFF_407.Q )
  );
  al_dffl _8737_ (
    .clk(CK),
    .d(\DFF_408.D ),
    .q(\DFF_408.Q )
  );
  al_dffl _8738_ (
    .clk(CK),
    .d(\DFF_409.D ),
    .q(\DFF_409.Q )
  );
  al_dffl _8739_ (
    .clk(CK),
    .d(\DFF_410.D ),
    .q(\DFF_410.Q )
  );
  al_dffl _8740_ (
    .clk(CK),
    .d(\DFF_411.D ),
    .q(\DFF_411.Q )
  );
  al_dffl _8741_ (
    .clk(CK),
    .d(\DFF_412.D ),
    .q(\DFF_412.Q )
  );
  al_dffl _8742_ (
    .clk(CK),
    .d(\DFF_413.D ),
    .q(\DFF_413.Q )
  );
  al_dffl _8743_ (
    .clk(CK),
    .d(\DFF_414.D ),
    .q(\DFF_414.Q )
  );
  al_dffl _8744_ (
    .clk(CK),
    .d(\DFF_415.D ),
    .q(\DFF_415.Q )
  );
  al_dffl _8745_ (
    .clk(CK),
    .d(\DFF_416.D ),
    .q(\DFF_416.Q )
  );
  al_dffl _8746_ (
    .clk(CK),
    .d(\DFF_417.D ),
    .q(\DFF_417.Q )
  );
  al_dffl _8747_ (
    .clk(CK),
    .d(\DFF_418.D ),
    .q(\DFF_418.Q )
  );
  al_dffl _8748_ (
    .clk(CK),
    .d(\DFF_419.D ),
    .q(\DFF_419.Q )
  );
  al_dffl _8749_ (
    .clk(CK),
    .d(\DFF_420.D ),
    .q(\DFF_420.Q )
  );
  al_dffl _8750_ (
    .clk(CK),
    .d(\DFF_421.D ),
    .q(\DFF_421.Q )
  );
  al_dffl _8751_ (
    .clk(CK),
    .d(\DFF_422.D ),
    .q(\DFF_422.Q )
  );
  al_dffl _8752_ (
    .clk(CK),
    .d(\DFF_423.D ),
    .q(\DFF_423.Q )
  );
  al_dffl _8753_ (
    .clk(CK),
    .d(\DFF_424.D ),
    .q(\DFF_424.Q )
  );
  al_dffl _8754_ (
    .clk(CK),
    .d(\DFF_425.D ),
    .q(\DFF_425.Q )
  );
  al_dffl _8755_ (
    .clk(CK),
    .d(\DFF_426.D ),
    .q(\DFF_426.Q )
  );
  al_dffl _8756_ (
    .clk(CK),
    .d(\DFF_427.D ),
    .q(\DFF_427.Q )
  );
  al_dffl _8757_ (
    .clk(CK),
    .d(\DFF_428.D ),
    .q(\DFF_428.Q )
  );
  al_dffl _8758_ (
    .clk(CK),
    .d(\DFF_429.D ),
    .q(\DFF_429.Q )
  );
  al_dffl _8759_ (
    .clk(CK),
    .d(\DFF_430.D ),
    .q(\DFF_430.Q )
  );
  al_dffl _8760_ (
    .clk(CK),
    .d(\DFF_431.D ),
    .q(\DFF_431.Q )
  );
  al_dffl _8761_ (
    .clk(CK),
    .d(\DFF_402.Q ),
    .q(\DFF_432.Q )
  );
  al_dffl _8762_ (
    .clk(CK),
    .d(\DFF_433.D ),
    .q(\DFF_433.Q )
  );
  al_dffl _8763_ (
    .clk(CK),
    .d(\DFF_442.D ),
    .q(\DFF_442.Q )
  );
  al_dffl _8764_ (
    .clk(CK),
    .d(\DFF_442.Q ),
    .q(\DFF_443.Q )
  );
  al_dffl _8765_ (
    .clk(CK),
    .d(\DFF_444.D ),
    .q(\DFF_444.Q )
  );
  al_dffl _8766_ (
    .clk(CK),
    .d(\DFF_445.D ),
    .q(\DFF_445.Q )
  );
  al_dffl _8767_ (
    .clk(CK),
    .d(\DFF_446.D ),
    .q(\DFF_446.Q )
  );
  al_dffl _8768_ (
    .clk(CK),
    .d(\DFF_447.D ),
    .q(\DFF_447.Q )
  );
  al_dffl _8769_ (
    .clk(CK),
    .d(\DFF_448.D ),
    .q(\DFF_448.Q )
  );
  al_dffl _8770_ (
    .clk(CK),
    .d(\DFF_449.D ),
    .q(\DFF_449.Q )
  );
  al_dffl _8771_ (
    .clk(CK),
    .d(\DFF_450.D ),
    .q(\DFF_450.Q )
  );
  al_dffl _8772_ (
    .clk(CK),
    .d(\DFF_451.D ),
    .q(\DFF_451.Q )
  );
  al_dffl _8773_ (
    .clk(CK),
    .d(\DFF_452.D ),
    .q(\DFF_452.Q )
  );
  al_dffl _8774_ (
    .clk(CK),
    .d(\DFF_453.D ),
    .q(\DFF_453.Q )
  );
  al_dffl _8775_ (
    .clk(CK),
    .d(\DFF_457.D ),
    .q(\DFF_457.Q )
  );
  al_dffl _8776_ (
    .clk(CK),
    .d(\DFF_458.D ),
    .q(\DFF_458.Q )
  );
  al_dffl _8777_ (
    .clk(CK),
    .d(\DFF_459.D ),
    .q(\DFF_459.Q )
  );
  al_dffl _8778_ (
    .clk(CK),
    .d(\DFF_460.D ),
    .q(\DFF_460.Q )
  );
  al_dffl _8779_ (
    .clk(CK),
    .d(\DFF_461.D ),
    .q(\DFF_461.Q )
  );
  al_dffl _8780_ (
    .clk(CK),
    .d(\DFF_462.D ),
    .q(\DFF_462.Q )
  );
  al_dffl _8781_ (
    .clk(CK),
    .d(\DFF_463.D ),
    .q(\DFF_463.Q )
  );
  al_dffl _8782_ (
    .clk(CK),
    .d(\DFF_464.D ),
    .q(\DFF_464.Q )
  );
  al_dffl _8783_ (
    .clk(CK),
    .d(\DFF_465.D ),
    .q(\DFF_465.Q )
  );
  al_dffl _8784_ (
    .clk(CK),
    .d(\DFF_466.D ),
    .q(\DFF_466.Q )
  );
  al_dffl _8785_ (
    .clk(CK),
    .d(\DFF_467.D ),
    .q(\DFF_467.Q )
  );
  al_dffl _8786_ (
    .clk(CK),
    .d(\DFF_468.D ),
    .q(\DFF_468.Q )
  );
  al_dffl _8787_ (
    .clk(CK),
    .d(\DFF_469.D ),
    .q(\DFF_469.Q )
  );
  al_dffl _8788_ (
    .clk(CK),
    .d(\DFF_470.D ),
    .q(\DFF_470.Q )
  );
  al_dffl _8789_ (
    .clk(CK),
    .d(\DFF_471.D ),
    .q(\DFF_471.Q )
  );
  al_dffl _8790_ (
    .clk(CK),
    .d(\DFF_472.D ),
    .q(\DFF_472.Q )
  );
  al_dffl _8791_ (
    .clk(CK),
    .d(\DFF_473.D ),
    .q(\DFF_473.Q )
  );
  al_dffl _8792_ (
    .clk(CK),
    .d(\DFF_474.D ),
    .q(\DFF_474.Q )
  );
  al_dffl _8793_ (
    .clk(CK),
    .d(\DFF_475.D ),
    .q(\DFF_475.Q )
  );
  al_dffl _8794_ (
    .clk(CK),
    .d(\DFF_476.D ),
    .q(\DFF_476.Q )
  );
  al_dffl _8795_ (
    .clk(CK),
    .d(\DFF_477.D ),
    .q(\DFF_477.Q )
  );
  al_dffl _8796_ (
    .clk(CK),
    .d(\DFF_478.D ),
    .q(\DFF_478.Q )
  );
  al_dffl _8797_ (
    .clk(CK),
    .d(\DFF_479.D ),
    .q(\DFF_479.Q )
  );
  al_dffl _8798_ (
    .clk(CK),
    .d(\DFF_480.D ),
    .q(\DFF_480.Q )
  );
  al_dffl _8799_ (
    .clk(CK),
    .d(\DFF_481.D ),
    .q(\DFF_481.Q )
  );
  al_dffl _8800_ (
    .clk(CK),
    .d(\DFF_482.D ),
    .q(\DFF_482.Q )
  );
  al_dffl _8801_ (
    .clk(CK),
    .d(\DFF_483.D ),
    .q(\DFF_483.Q )
  );
  al_dffl _8802_ (
    .clk(CK),
    .d(\DFF_484.D ),
    .q(\DFF_484.Q )
  );
  al_dffl _8803_ (
    .clk(CK),
    .d(\DFF_485.D ),
    .q(\DFF_485.Q )
  );
  al_dffl _8804_ (
    .clk(CK),
    .d(\DFF_486.D ),
    .q(\DFF_486.Q )
  );
  al_dffl _8805_ (
    .clk(CK),
    .d(\DFF_487.D ),
    .q(\DFF_487.Q )
  );
  al_dffl _8806_ (
    .clk(CK),
    .d(\DFF_488.D ),
    .q(\DFF_488.Q )
  );
  al_dffl _8807_ (
    .clk(CK),
    .d(\DFF_489.D ),
    .q(\DFF_489.Q )
  );
  al_dffl _8808_ (
    .clk(CK),
    .d(\DFF_490.D ),
    .q(\DFF_490.Q )
  );
  al_dffl _8809_ (
    .clk(CK),
    .d(\DFF_491.D ),
    .q(\DFF_491.Q )
  );
  al_dffl _8810_ (
    .clk(CK),
    .d(\DFF_492.D ),
    .q(\DFF_492.Q )
  );
  al_dffl _8811_ (
    .clk(CK),
    .d(\DFF_493.D ),
    .q(\DFF_493.Q )
  );
  al_dffl _8812_ (
    .clk(CK),
    .d(\DFF_494.D ),
    .q(\DFF_494.Q )
  );
  al_dffl _8813_ (
    .clk(CK),
    .d(\DFF_495.D ),
    .q(\DFF_495.Q )
  );
  al_dffl _8814_ (
    .clk(CK),
    .d(\DFF_496.D ),
    .q(\DFF_496.Q )
  );
  al_dffl _8815_ (
    .clk(CK),
    .d(\DFF_497.D ),
    .q(\DFF_497.Q )
  );
  al_dffl _8816_ (
    .clk(CK),
    .d(\DFF_498.D ),
    .q(\DFF_498.Q )
  );
  al_dffl _8817_ (
    .clk(CK),
    .d(\DFF_499.D ),
    .q(\DFF_499.Q )
  );
  al_dffl _8818_ (
    .clk(CK),
    .d(\DFF_500.D ),
    .q(\DFF_500.Q )
  );
  al_dffl _8819_ (
    .clk(CK),
    .d(\DFF_501.D ),
    .q(\DFF_501.Q )
  );
  al_dffl _8820_ (
    .clk(CK),
    .d(\DFF_502.D ),
    .q(\DFF_502.Q )
  );
  al_dffl _8821_ (
    .clk(CK),
    .d(\DFF_503.D ),
    .q(\DFF_503.Q )
  );
  al_dffl _8822_ (
    .clk(CK),
    .d(\DFF_504.D ),
    .q(\DFF_504.Q )
  );
  al_dffl _8823_ (
    .clk(CK),
    .d(\DFF_505.D ),
    .q(\DFF_505.Q )
  );
  al_dffl _8824_ (
    .clk(CK),
    .d(\DFF_506.D ),
    .q(\DFF_506.Q )
  );
  al_dffl _8825_ (
    .clk(CK),
    .d(\DFF_507.D ),
    .q(\DFF_507.Q )
  );
  al_dffl _8826_ (
    .clk(CK),
    .d(\DFF_508.D ),
    .q(\DFF_508.Q )
  );
  al_dffl _8827_ (
    .clk(CK),
    .d(\DFF_509.D ),
    .q(\DFF_509.Q )
  );
  al_dffl _8828_ (
    .clk(CK),
    .d(\DFF_510.D ),
    .q(\DFF_510.Q )
  );
  al_dffl _8829_ (
    .clk(CK),
    .d(\DFF_514.D ),
    .q(\DFF_514.Q )
  );
  al_dffl _8830_ (
    .clk(CK),
    .d(\DFF_515.D ),
    .q(\DFF_515.Q )
  );
  al_dffl _8831_ (
    .clk(CK),
    .d(\DFF_516.D ),
    .q(\DFF_516.Q )
  );
  al_dffl _8832_ (
    .clk(CK),
    .d(\DFF_517.D ),
    .q(\DFF_517.Q )
  );
  al_dffl _8833_ (
    .clk(CK),
    .d(\DFF_518.D ),
    .q(\DFF_518.Q )
  );
  al_dffl _8834_ (
    .clk(CK),
    .d(\DFF_519.D ),
    .q(\DFF_519.Q )
  );
  al_dffl _8835_ (
    .clk(CK),
    .d(\DFF_520.D ),
    .q(\DFF_520.Q )
  );
  al_dffl _8836_ (
    .clk(CK),
    .d(\DFF_521.D ),
    .q(\DFF_521.Q )
  );
  al_dffl _8837_ (
    .clk(CK),
    .d(\DFF_522.D ),
    .q(\DFF_522.Q )
  );
  al_dffl _8838_ (
    .clk(CK),
    .d(\DFF_523.D ),
    .q(\DFF_523.Q )
  );
  al_dffl _8839_ (
    .clk(CK),
    .d(\DFF_524.D ),
    .q(\DFF_524.Q )
  );
  al_dffl _8840_ (
    .clk(CK),
    .d(\DFF_525.D ),
    .q(\DFF_525.Q )
  );
  al_dffl _8841_ (
    .clk(CK),
    .d(\DFF_526.D ),
    .q(\DFF_526.Q )
  );
  al_dffl _8842_ (
    .clk(CK),
    .d(\DFF_527.D ),
    .q(\DFF_527.Q )
  );
  al_dffl _8843_ (
    .clk(CK),
    .d(\DFF_528.D ),
    .q(\DFF_528.Q )
  );
  al_dffl _8844_ (
    .clk(CK),
    .d(\DFF_529.D ),
    .q(\DFF_529.Q )
  );
  al_dffl _8845_ (
    .clk(CK),
    .d(\DFF_530.D ),
    .q(\DFF_530.Q )
  );
  al_dffl _8846_ (
    .clk(CK),
    .d(\DFF_531.D ),
    .q(\DFF_531.Q )
  );
  al_dffl _8847_ (
    .clk(CK),
    .d(\DFF_532.D ),
    .q(\DFF_532.Q )
  );
  al_dffl _8848_ (
    .clk(CK),
    .d(\DFF_533.D ),
    .q(\DFF_533.Q )
  );
  al_dffl _8849_ (
    .clk(CK),
    .d(\DFF_534.D ),
    .q(\DFF_534.Q )
  );
  al_dffl _8850_ (
    .clk(CK),
    .d(\DFF_535.D ),
    .q(\DFF_535.Q )
  );
  al_dffl _8851_ (
    .clk(CK),
    .d(\DFF_536.D ),
    .q(\DFF_536.Q )
  );
  al_dffl _8852_ (
    .clk(CK),
    .d(\DFF_537.D ),
    .q(\DFF_537.Q )
  );
  al_dffl _8853_ (
    .clk(CK),
    .d(\DFF_538.D ),
    .q(\DFF_538.Q )
  );
  al_dffl _8854_ (
    .clk(CK),
    .d(\DFF_539.D ),
    .q(\DFF_539.Q )
  );
  al_dffl _8855_ (
    .clk(CK),
    .d(\DFF_540.D ),
    .q(\DFF_540.Q )
  );
  al_dffl _8856_ (
    .clk(CK),
    .d(\DFF_541.D ),
    .q(\DFF_541.Q )
  );
  al_dffl _8857_ (
    .clk(CK),
    .d(\DFF_542.D ),
    .q(\DFF_542.Q )
  );
  al_dffl _8858_ (
    .clk(CK),
    .d(\DFF_543.D ),
    .q(\DFF_543.Q )
  );
  al_dffl _8859_ (
    .clk(CK),
    .d(\DFF_544.D ),
    .q(\DFF_544.Q )
  );
  al_dffl _8860_ (
    .clk(CK),
    .d(\DFF_545.D ),
    .q(\DFF_545.Q )
  );
  al_dffl _8861_ (
    .clk(CK),
    .d(\DFF_546.D ),
    .q(\DFF_546.Q )
  );
  al_dffl _8862_ (
    .clk(CK),
    .d(\DFF_547.D ),
    .q(\DFF_547.Q )
  );
  al_dffl _8863_ (
    .clk(CK),
    .d(\DFF_548.D ),
    .q(\DFF_548.Q )
  );
  al_dffl _8864_ (
    .clk(CK),
    .d(\DFF_549.D ),
    .q(\DFF_549.Q )
  );
  al_dffl _8865_ (
    .clk(CK),
    .d(\DFF_550.D ),
    .q(\DFF_550.Q )
  );
  al_dffl _8866_ (
    .clk(CK),
    .d(\DFF_551.D ),
    .q(\DFF_551.Q )
  );
  al_dffl _8867_ (
    .clk(CK),
    .d(\DFF_552.D ),
    .q(\DFF_552.Q )
  );
  al_dffl _8868_ (
    .clk(CK),
    .d(\DFF_553.D ),
    .q(\DFF_553.Q )
  );
  al_dffl _8869_ (
    .clk(CK),
    .d(\DFF_554.D ),
    .q(\DFF_554.Q )
  );
  al_dffl _8870_ (
    .clk(CK),
    .d(\DFF_555.D ),
    .q(\DFF_555.Q )
  );
  al_dffl _8871_ (
    .clk(CK),
    .d(\DFF_556.D ),
    .q(\DFF_556.Q )
  );
  al_dffl _8872_ (
    .clk(CK),
    .d(\DFF_557.D ),
    .q(\DFF_557.Q )
  );
  al_dffl _8873_ (
    .clk(CK),
    .d(\DFF_558.D ),
    .q(\DFF_558.Q )
  );
  al_dffl _8874_ (
    .clk(CK),
    .d(\DFF_559.D ),
    .q(\DFF_559.Q )
  );
  al_dffl _8875_ (
    .clk(CK),
    .d(\DFF_560.D ),
    .q(\DFF_560.Q )
  );
  al_dffl _8876_ (
    .clk(CK),
    .d(\DFF_561.D ),
    .q(\DFF_561.Q )
  );
  al_dffl _8877_ (
    .clk(CK),
    .d(\DFF_562.D ),
    .q(\DFF_562.Q )
  );
  al_dffl _8878_ (
    .clk(CK),
    .d(\DFF_563.D ),
    .q(\DFF_563.Q )
  );
  al_dffl _8879_ (
    .clk(CK),
    .d(\DFF_564.D ),
    .q(\DFF_564.Q )
  );
  al_dffl _8880_ (
    .clk(CK),
    .d(\DFF_565.D ),
    .q(\DFF_565.Q )
  );
  al_dffl _8881_ (
    .clk(CK),
    .d(\DFF_566.D ),
    .q(\DFF_566.Q )
  );
  al_dffl _8882_ (
    .clk(CK),
    .d(\DFF_567.D ),
    .q(\DFF_567.Q )
  );
  al_dffl _8883_ (
    .clk(CK),
    .d(\DFF_568.D ),
    .q(\DFF_568.Q )
  );
  al_dffl _8884_ (
    .clk(CK),
    .d(\DFF_569.D ),
    .q(\DFF_569.Q )
  );
  al_dffl _8885_ (
    .clk(CK),
    .d(\DFF_570.D ),
    .q(\DFF_570.Q )
  );
  al_dffl _8886_ (
    .clk(CK),
    .d(\DFF_571.D ),
    .q(\DFF_571.Q )
  );
  al_dffl _8887_ (
    .clk(CK),
    .d(\DFF_572.D ),
    .q(\DFF_572.Q )
  );
  al_dffl _8888_ (
    .clk(CK),
    .d(\DFF_573.D ),
    .q(\DFF_573.Q )
  );
  al_dffl _8889_ (
    .clk(CK),
    .d(\DFF_574.D ),
    .q(\DFF_574.Q )
  );
  al_dffl _8890_ (
    .clk(CK),
    .d(\DFF_575.D ),
    .q(\DFF_575.Q )
  );
  al_dffl _8891_ (
    .clk(CK),
    .d(\DFF_576.D ),
    .q(\DFF_576.Q )
  );
  al_dffl _8892_ (
    .clk(CK),
    .d(\DFF_577.D ),
    .q(\DFF_577.Q )
  );
  al_dffl _8893_ (
    .clk(CK),
    .d(\DFF_578.D ),
    .q(\DFF_578.Q )
  );
  al_dffl _8894_ (
    .clk(CK),
    .d(\DFF_579.D ),
    .q(\DFF_579.Q )
  );
  al_dffl _8895_ (
    .clk(CK),
    .d(\DFF_580.D ),
    .q(\DFF_580.Q )
  );
  al_dffl _8896_ (
    .clk(CK),
    .d(\DFF_581.D ),
    .q(\DFF_581.Q )
  );
  al_dffl _8897_ (
    .clk(CK),
    .d(\DFF_582.D ),
    .q(\DFF_582.Q )
  );
  al_dffl _8898_ (
    .clk(CK),
    .d(\DFF_583.D ),
    .q(\DFF_583.Q )
  );
  al_dffl _8899_ (
    .clk(CK),
    .d(\DFF_584.D ),
    .q(\DFF_584.Q )
  );
  al_dffl _8900_ (
    .clk(CK),
    .d(\DFF_585.D ),
    .q(\DFF_585.Q )
  );
  al_dffl _8901_ (
    .clk(CK),
    .d(\DFF_586.D ),
    .q(\DFF_586.Q )
  );
  al_dffl _8902_ (
    .clk(CK),
    .d(\DFF_587.D ),
    .q(\DFF_587.Q )
  );
  al_dffl _8903_ (
    .clk(CK),
    .d(\DFF_588.D ),
    .q(\DFF_588.Q )
  );
  al_dffl _8904_ (
    .clk(CK),
    .d(\DFF_589.D ),
    .q(\DFF_589.Q )
  );
  al_dffl _8905_ (
    .clk(CK),
    .d(\DFF_590.D ),
    .q(\DFF_590.Q )
  );
  al_dffl _8906_ (
    .clk(CK),
    .d(\DFF_591.D ),
    .q(\DFF_591.Q )
  );
  al_dffl _8907_ (
    .clk(CK),
    .d(\DFF_592.D ),
    .q(\DFF_592.Q )
  );
  al_dffl _8908_ (
    .clk(CK),
    .d(\DFF_593.D ),
    .q(\DFF_593.Q )
  );
  al_dffl _8909_ (
    .clk(CK),
    .d(\DFF_594.D ),
    .q(\DFF_594.Q )
  );
  al_dffl _8910_ (
    .clk(CK),
    .d(\DFF_595.D ),
    .q(\DFF_595.Q )
  );
  al_dffl _8911_ (
    .clk(CK),
    .d(\DFF_603.D ),
    .q(\DFF_603.Q )
  );
  al_dffl _8912_ (
    .clk(CK),
    .d(\DFF_604.D ),
    .q(\DFF_604.Q )
  );
  al_dffl _8913_ (
    .clk(CK),
    .d(\DFF_605.D ),
    .q(\DFF_605.Q )
  );
  al_dffl _8914_ (
    .clk(CK),
    .d(\DFF_606.D ),
    .q(\DFF_606.Q )
  );
  al_dffl _8915_ (
    .clk(CK),
    .d(\DFF_607.D ),
    .q(\DFF_607.Q )
  );
  al_dffl _8916_ (
    .clk(CK),
    .d(\DFF_608.D ),
    .q(\DFF_608.Q )
  );
  al_dffl _8917_ (
    .clk(CK),
    .d(\DFF_609.D ),
    .q(\DFF_609.Q )
  );
  al_dffl _8918_ (
    .clk(CK),
    .d(\DFF_610.D ),
    .q(\DFF_610.Q )
  );
  al_dffl _8919_ (
    .clk(CK),
    .d(\DFF_611.D ),
    .q(\DFF_611.Q )
  );
  al_dffl _8920_ (
    .clk(CK),
    .d(\DFF_612.D ),
    .q(\DFF_612.Q )
  );
  al_dffl _8921_ (
    .clk(CK),
    .d(\DFF_613.D ),
    .q(\DFF_613.Q )
  );
  al_dffl _8922_ (
    .clk(CK),
    .d(\DFF_614.D ),
    .q(\DFF_614.Q )
  );
  al_dffl _8923_ (
    .clk(CK),
    .d(\DFF_615.D ),
    .q(\DFF_615.Q )
  );
  al_dffl _8924_ (
    .clk(CK),
    .d(\DFF_616.D ),
    .q(\DFF_616.Q )
  );
  al_dffl _8925_ (
    .clk(CK),
    .d(\DFF_617.D ),
    .q(\DFF_617.Q )
  );
  al_dffl _8926_ (
    .clk(CK),
    .d(\DFF_618.D ),
    .q(\DFF_618.Q )
  );
  al_dffl _8927_ (
    .clk(CK),
    .d(\DFF_619.D ),
    .q(\DFF_619.Q )
  );
  al_dffl _8928_ (
    .clk(CK),
    .d(\DFF_620.D ),
    .q(\DFF_620.Q )
  );
  al_dffl _8929_ (
    .clk(CK),
    .d(\DFF_621.D ),
    .q(\DFF_621.Q )
  );
  al_dffl _8930_ (
    .clk(CK),
    .d(\DFF_622.D ),
    .q(\DFF_622.Q )
  );
  al_dffl _8931_ (
    .clk(CK),
    .d(\DFF_623.D ),
    .q(\DFF_623.Q )
  );
  al_dffl _8932_ (
    .clk(CK),
    .d(\DFF_624.D ),
    .q(\DFF_624.Q )
  );
  al_dffl _8933_ (
    .clk(CK),
    .d(\DFF_625.D ),
    .q(\DFF_625.Q )
  );
  al_dffl _8934_ (
    .clk(CK),
    .d(\DFF_626.D ),
    .q(\DFF_626.Q )
  );
  al_dffl _8935_ (
    .clk(CK),
    .d(\DFF_627.D ),
    .q(\DFF_627.Q )
  );
  al_dffl _8936_ (
    .clk(CK),
    .d(\DFF_628.D ),
    .q(\DFF_628.Q )
  );
  al_dffl _8937_ (
    .clk(CK),
    .d(\DFF_629.D ),
    .q(\DFF_629.Q )
  );
  al_dffl _8938_ (
    .clk(CK),
    .d(\DFF_630.D ),
    .q(\DFF_630.Q )
  );
  al_dffl _8939_ (
    .clk(CK),
    .d(\DFF_631.D ),
    .q(\DFF_631.Q )
  );
  al_dffl _8940_ (
    .clk(CK),
    .d(\DFF_632.D ),
    .q(\DFF_632.Q )
  );
  al_dffl _8941_ (
    .clk(CK),
    .d(\DFF_633.D ),
    .q(\DFF_633.Q )
  );
  al_dffl _8942_ (
    .clk(CK),
    .d(\DFF_634.D ),
    .q(\DFF_634.Q )
  );
  al_dffl _8943_ (
    .clk(CK),
    .d(\DFF_635.D ),
    .q(\DFF_635.Q )
  );
  al_dffl _8944_ (
    .clk(CK),
    .d(\DFF_636.D ),
    .q(\DFF_636.Q )
  );
  al_dffl _8945_ (
    .clk(CK),
    .d(\DFF_637.D ),
    .q(\DFF_637.Q )
  );
  al_dffl _8946_ (
    .clk(CK),
    .d(\DFF_638.D ),
    .q(\DFF_638.Q )
  );
  al_dffl _8947_ (
    .clk(CK),
    .d(\DFF_639.D ),
    .q(\DFF_639.Q )
  );
  al_dffl _8948_ (
    .clk(CK),
    .d(\DFF_640.D ),
    .q(\DFF_640.Q )
  );
  al_dffl _8949_ (
    .clk(CK),
    .d(\DFF_641.D ),
    .q(\DFF_641.Q )
  );
  al_dffl _8950_ (
    .clk(CK),
    .d(\DFF_642.D ),
    .q(\DFF_642.Q )
  );
  al_dffl _8951_ (
    .clk(CK),
    .d(\DFF_643.D ),
    .q(\DFF_643.Q )
  );
  al_dffl _8952_ (
    .clk(CK),
    .d(\DFF_644.D ),
    .q(\DFF_644.Q )
  );
  al_dffl _8953_ (
    .clk(CK),
    .d(\DFF_645.D ),
    .q(\DFF_645.Q )
  );
  al_dffl _8954_ (
    .clk(CK),
    .d(\DFF_646.D ),
    .q(\DFF_646.Q )
  );
  al_dffl _8955_ (
    .clk(CK),
    .d(\DFF_647.D ),
    .q(\DFF_647.Q )
  );
  al_dffl _8956_ (
    .clk(CK),
    .d(\DFF_648.D ),
    .q(\DFF_648.Q )
  );
  al_dffl _8957_ (
    .clk(CK),
    .d(\DFF_648.Q ),
    .q(\DFF_649.Q )
  );
  al_dffl _8958_ (
    .clk(CK),
    .d(\DFF_650.D ),
    .q(\DFF_650.Q )
  );
  al_dffl _8959_ (
    .clk(CK),
    .d(\DFF_650.Q ),
    .q(\DFF_651.Q )
  );
  al_dffl _8960_ (
    .clk(CK),
    .d(\DFF_652.D ),
    .q(\DFF_652.Q )
  );
  al_dffl _8961_ (
    .clk(CK),
    .d(\DFF_652.Q ),
    .q(\DFF_653.Q )
  );
  al_dffl _8962_ (
    .clk(CK),
    .d(\DFF_654.D ),
    .q(\DFF_654.Q )
  );
  al_dffl _8963_ (
    .clk(CK),
    .d(\DFF_654.Q ),
    .q(\DFF_655.Q )
  );
  al_dffl _8964_ (
    .clk(CK),
    .d(\DFF_656.D ),
    .q(\DFF_656.Q )
  );
  al_dffl _8965_ (
    .clk(CK),
    .d(\DFF_656.Q ),
    .q(\DFF_657.Q )
  );
  al_dffl _8966_ (
    .clk(CK),
    .d(\DFF_658.D ),
    .q(\DFF_658.Q )
  );
  al_dffl _8967_ (
    .clk(CK),
    .d(\DFF_658.Q ),
    .q(\DFF_659.Q )
  );
  al_dffl _8968_ (
    .clk(CK),
    .d(\DFF_660.D ),
    .q(\DFF_660.Q )
  );
  al_dffl _8969_ (
    .clk(CK),
    .d(\DFF_660.Q ),
    .q(\DFF_661.Q )
  );
  al_dffl _8970_ (
    .clk(CK),
    .d(\DFF_662.D ),
    .q(\DFF_662.Q )
  );
  al_dffl _8971_ (
    .clk(CK),
    .d(\DFF_662.Q ),
    .q(\DFF_663.Q )
  );
  al_dffl _8972_ (
    .clk(CK),
    .d(\DFF_64.Q ),
    .q(\DFF_664.Q )
  );
  al_dffl _8973_ (
    .clk(CK),
    .d(\DFF_664.Q ),
    .q(\DFF_665.Q )
  );
  al_dffl _8974_ (
    .clk(CK),
    .d(\DFF_666.D ),
    .q(\DFF_666.Q )
  );
  al_dffl _8975_ (
    .clk(CK),
    .d(\DFF_667.D ),
    .q(\DFF_667.Q )
  );
  al_dffl _8976_ (
    .clk(CK),
    .d(\DFF_678.D ),
    .q(\DFF_678.Q )
  );
  al_dffl _8977_ (
    .clk(CK),
    .d(\DFF_603.Q ),
    .q(\DFF_679.Q )
  );
  al_dffl _8978_ (
    .clk(CK),
    .d(\DFF_679.Q ),
    .q(\DFF_680.Q )
  );
  al_dffl _8979_ (
    .clk(CK),
    .d(\DFF_604.Q ),
    .q(\DFF_681.Q )
  );
  al_dffl _8980_ (
    .clk(CK),
    .d(\DFF_681.Q ),
    .q(\DFF_682.Q )
  );
  al_dffl _8981_ (
    .clk(CK),
    .d(\DFF_605.Q ),
    .q(\DFF_683.Q )
  );
  al_dffl _8982_ (
    .clk(CK),
    .d(\DFF_683.Q ),
    .q(\DFF_684.Q )
  );
  al_dffl _8983_ (
    .clk(CK),
    .d(\DFF_606.Q ),
    .q(\DFF_685.Q )
  );
  al_dffl _8984_ (
    .clk(CK),
    .d(\DFF_685.Q ),
    .q(\DFF_686.Q )
  );
  al_dffl _8985_ (
    .clk(CK),
    .d(\DFF_607.Q ),
    .q(\DFF_687.Q )
  );
  al_dffl _8986_ (
    .clk(CK),
    .d(\DFF_687.Q ),
    .q(\DFF_688.Q )
  );
  al_dffl _8987_ (
    .clk(CK),
    .d(\DFF_608.Q ),
    .q(\DFF_689.Q )
  );
  al_dffl _8988_ (
    .clk(CK),
    .d(\DFF_689.Q ),
    .q(\DFF_690.Q )
  );
  al_dffl _8989_ (
    .clk(CK),
    .d(\DFF_609.Q ),
    .q(\DFF_691.Q )
  );
  al_dffl _8990_ (
    .clk(CK),
    .d(\DFF_691.Q ),
    .q(\DFF_692.Q )
  );
  al_dffl _8991_ (
    .clk(CK),
    .d(\DFF_610.Q ),
    .q(\DFF_693.Q )
  );
  al_dffl _8992_ (
    .clk(CK),
    .d(\DFF_693.Q ),
    .q(\DFF_694.Q )
  );
  al_dffl _8993_ (
    .clk(CK),
    .d(\DFF_611.Q ),
    .q(\DFF_695.Q )
  );
  al_dffl _8994_ (
    .clk(CK),
    .d(\DFF_695.Q ),
    .q(\DFF_696.Q )
  );
  al_dffl _8995_ (
    .clk(CK),
    .d(\DFF_612.Q ),
    .q(\DFF_697.Q )
  );
  al_dffl _8996_ (
    .clk(CK),
    .d(\DFF_697.Q ),
    .q(\DFF_698.Q )
  );
  al_dffl _8997_ (
    .clk(CK),
    .d(\DFF_613.Q ),
    .q(\DFF_699.Q )
  );
  al_dffl _8998_ (
    .clk(CK),
    .d(\DFF_699.Q ),
    .q(\DFF_700.Q )
  );
  al_dffl _8999_ (
    .clk(CK),
    .d(\DFF_614.Q ),
    .q(\DFF_701.Q )
  );
  al_dffl _9000_ (
    .clk(CK),
    .d(\DFF_701.Q ),
    .q(\DFF_702.Q )
  );
  al_dffl _9001_ (
    .clk(CK),
    .d(\DFF_709.D ),
    .q(\DFF_709.Q )
  );
  al_dffl _9002_ (
    .clk(CK),
    .d(\DFF_710.D ),
    .q(\DFF_710.Q )
  );
  al_dffl _9003_ (
    .clk(CK),
    .d(\DFF_711.D ),
    .q(\DFF_711.Q )
  );
  al_dffl _9004_ (
    .clk(CK),
    .d(\DFF_712.D ),
    .q(\DFF_712.Q )
  );
  al_dffl _9005_ (
    .clk(CK),
    .d(\DFF_712.Q ),
    .q(\DFF_713.Q )
  );
  al_dffl _9006_ (
    .clk(CK),
    .d(\DFF_713.Q ),
    .q(\DFF_714.Q )
  );
  al_dffl _9007_ (
    .clk(CK),
    .d(\DFF_733.Q ),
    .q(\DFF_715.Q )
  );
  al_dffl _9008_ (
    .clk(CK),
    .d(\DFF_715.Q ),
    .q(\DFF_716.Q )
  );
  al_dffl _9009_ (
    .clk(CK),
    .d(\DFF_734.Q ),
    .q(\DFF_717.Q )
  );
  al_dffl _9010_ (
    .clk(CK),
    .d(\DFF_717.Q ),
    .q(\DFF_718.Q )
  );
  al_dffl _9011_ (
    .clk(CK),
    .d(\DFF_735.Q ),
    .q(\DFF_719.Q )
  );
  al_dffl _9012_ (
    .clk(CK),
    .d(\DFF_719.Q ),
    .q(\DFF_720.Q )
  );
  al_dffl _9013_ (
    .clk(CK),
    .d(\DFF_742.Q ),
    .q(\DFF_721.Q )
  );
  al_dffl _9014_ (
    .clk(CK),
    .d(\DFF_721.Q ),
    .q(\DFF_722.Q )
  );
  al_dffl _9015_ (
    .clk(CK),
    .d(\DFF_743.Q ),
    .q(\DFF_723.Q )
  );
  al_dffl _9016_ (
    .clk(CK),
    .d(\DFF_723.Q ),
    .q(\DFF_724.Q )
  );
  al_dffl _9017_ (
    .clk(CK),
    .d(\DFF_744.Q ),
    .q(\DFF_725.Q )
  );
  al_dffl _9018_ (
    .clk(CK),
    .d(\DFF_725.Q ),
    .q(\DFF_726.Q )
  );
  al_dffl _9019_ (
    .clk(CK),
    .d(\DFF_730.D ),
    .q(\DFF_730.Q )
  );
  al_dffl _9020_ (
    .clk(CK),
    .d(\DFF_731.D ),
    .q(\DFF_731.Q )
  );
  al_dffl _9021_ (
    .clk(CK),
    .d(\DFF_732.D ),
    .q(\DFF_732.Q )
  );
  al_dffl _9022_ (
    .clk(CK),
    .d(\DFF_733.D ),
    .q(\DFF_733.Q )
  );
  al_dffl _9023_ (
    .clk(CK),
    .d(\DFF_734.D ),
    .q(\DFF_734.Q )
  );
  al_dffl _9024_ (
    .clk(CK),
    .d(\DFF_735.D ),
    .q(\DFF_735.Q )
  );
  al_dffl _9025_ (
    .clk(CK),
    .d(\DFF_736.D ),
    .q(\DFF_736.Q )
  );
  al_dffl _9026_ (
    .clk(CK),
    .d(\DFF_737.D ),
    .q(\DFF_737.Q )
  );
  al_dffl _9027_ (
    .clk(CK),
    .d(\DFF_738.D ),
    .q(\DFF_738.Q )
  );
  al_dffl _9028_ (
    .clk(CK),
    .d(\DFF_739.D ),
    .q(\DFF_739.Q )
  );
  al_dffl _9029_ (
    .clk(CK),
    .d(\DFF_740.D ),
    .q(\DFF_740.Q )
  );
  al_dffl _9030_ (
    .clk(CK),
    .d(\DFF_741.D ),
    .q(\DFF_741.Q )
  );
  al_dffl _9031_ (
    .clk(CK),
    .d(\DFF_742.D ),
    .q(\DFF_742.Q )
  );
  al_dffl _9032_ (
    .clk(CK),
    .d(\DFF_743.D ),
    .q(\DFF_743.Q )
  );
  al_dffl _9033_ (
    .clk(CK),
    .d(\DFF_744.D ),
    .q(\DFF_744.Q )
  );
  al_dffl _9034_ (
    .clk(CK),
    .d(\DFF_745.D ),
    .q(\DFF_745.Q )
  );
  al_dffl _9035_ (
    .clk(CK),
    .d(\DFF_745.Q ),
    .q(\DFF_746.Q )
  );
  al_dffl _9036_ (
    .clk(CK),
    .d(\DFF_746.Q ),
    .q(\DFF_747.Q )
  );
  al_dffl _9037_ (
    .clk(CK),
    .d(\DFF_748.D ),
    .q(\DFF_748.Q )
  );
  al_dffl _9038_ (
    .clk(CK),
    .d(\DFF_748.Q ),
    .q(\DFF_749.Q )
  );
  al_dffl _9039_ (
    .clk(CK),
    .d(\DFF_750.D ),
    .q(\DFF_750.Q )
  );
  al_dffl _9040_ (
    .clk(CK),
    .d(\DFF_751.D ),
    .q(\DFF_751.Q )
  );
  al_dffl _9041_ (
    .clk(CK),
    .d(\DFF_751.Q ),
    .q(\DFF_752.Q )
  );
  al_dffl _9042_ (
    .clk(CK),
    .d(\DFF_753.D ),
    .q(\DFF_753.Q )
  );
  al_dffl _9043_ (
    .clk(CK),
    .d(\DFF_753.Q ),
    .q(\DFF_754.Q )
  );
  al_dffl _9044_ (
    .clk(CK),
    .d(\DFF_755.D ),
    .q(\DFF_755.Q )
  );
  al_dffl _9045_ (
    .clk(CK),
    .d(\DFF_756.D ),
    .q(\DFF_756.Q )
  );
  al_dffl _9046_ (
    .clk(CK),
    .d(\DFF_757.D ),
    .q(\DFF_757.Q )
  );
  al_dffl _9047_ (
    .clk(CK),
    .d(\DFF_758.D ),
    .q(\DFF_758.Q )
  );
  al_dffl _9048_ (
    .clk(CK),
    .d(\DFF_759.D ),
    .q(\DFF_759.Q )
  );
  al_dffl _9049_ (
    .clk(CK),
    .d(\DFF_760.D ),
    .q(\DFF_760.Q )
  );
  al_dffl _9050_ (
    .clk(CK),
    .d(\DFF_761.D ),
    .q(\DFF_761.Q )
  );
  al_dffl _9051_ (
    .clk(CK),
    .d(\DFF_762.D ),
    .q(\DFF_762.Q )
  );
  al_dffl _9052_ (
    .clk(CK),
    .d(\DFF_763.D ),
    .q(\DFF_763.Q )
  );
  al_dffl _9053_ (
    .clk(CK),
    .d(\DFF_764.D ),
    .q(\DFF_764.Q )
  );
  al_dffl _9054_ (
    .clk(CK),
    .d(\DFF_765.D ),
    .q(\DFF_765.Q )
  );
  al_dffl _9055_ (
    .clk(CK),
    .d(\DFF_766.D ),
    .q(\DFF_766.Q )
  );
  al_dffl _9056_ (
    .clk(CK),
    .d(\DFF_767.D ),
    .q(\DFF_767.Q )
  );
  al_dffl _9057_ (
    .clk(CK),
    .d(\DFF_768.D ),
    .q(\DFF_768.Q )
  );
  al_dffl _9058_ (
    .clk(CK),
    .d(\DFF_769.D ),
    .q(\DFF_769.Q )
  );
  al_dffl _9059_ (
    .clk(CK),
    .d(\DFF_770.D ),
    .q(\DFF_770.Q )
  );
  al_dffl _9060_ (
    .clk(CK),
    .d(\DFF_771.D ),
    .q(\DFF_771.Q )
  );
  al_dffl _9061_ (
    .clk(CK),
    .d(\DFF_772.D ),
    .q(\DFF_772.Q )
  );
  al_dffl _9062_ (
    .clk(CK),
    .d(\DFF_773.D ),
    .q(\DFF_773.Q )
  );
  al_dffl _9063_ (
    .clk(CK),
    .d(\DFF_774.D ),
    .q(\DFF_774.Q )
  );
  al_dffl _9064_ (
    .clk(CK),
    .d(\DFF_775.D ),
    .q(\DFF_775.Q )
  );
  al_dffl _9065_ (
    .clk(CK),
    .d(\DFF_776.D ),
    .q(\DFF_776.Q )
  );
  al_dffl _9066_ (
    .clk(CK),
    .d(\DFF_777.D ),
    .q(\DFF_777.Q )
  );
  al_dffl _9067_ (
    .clk(CK),
    .d(\DFF_778.D ),
    .q(\DFF_778.Q )
  );
  al_dffl _9068_ (
    .clk(CK),
    .d(\DFF_779.D ),
    .q(\DFF_779.Q )
  );
  al_dffl _9069_ (
    .clk(CK),
    .d(\DFF_780.D ),
    .q(\DFF_780.Q )
  );
  al_dffl _9070_ (
    .clk(CK),
    .d(\DFF_781.D ),
    .q(\DFF_781.Q )
  );
  al_dffl _9071_ (
    .clk(CK),
    .d(\DFF_752.Q ),
    .q(\DFF_782.Q )
  );
  al_dffl _9072_ (
    .clk(CK),
    .d(\DFF_783.D ),
    .q(\DFF_783.Q )
  );
  al_dffl _9073_ (
    .clk(CK),
    .d(\DFF_792.D ),
    .q(\DFF_792.Q )
  );
  al_dffl _9074_ (
    .clk(CK),
    .d(\DFF_792.Q ),
    .q(\DFF_793.Q )
  );
  al_dffl _9075_ (
    .clk(CK),
    .d(\DFF_794.D ),
    .q(\DFF_794.Q )
  );
  al_dffl _9076_ (
    .clk(CK),
    .d(\DFF_795.D ),
    .q(\DFF_795.Q )
  );
  al_dffl _9077_ (
    .clk(CK),
    .d(\DFF_796.D ),
    .q(\DFF_796.Q )
  );
  al_dffl _9078_ (
    .clk(CK),
    .d(\DFF_797.D ),
    .q(\DFF_797.Q )
  );
  al_dffl _9079_ (
    .clk(CK),
    .d(\DFF_798.D ),
    .q(\DFF_798.Q )
  );
  al_dffl _9080_ (
    .clk(CK),
    .d(\DFF_799.D ),
    .q(\DFF_799.Q )
  );
  al_dffl _9081_ (
    .clk(CK),
    .d(\DFF_800.D ),
    .q(\DFF_800.Q )
  );
  al_dffl _9082_ (
    .clk(CK),
    .d(\DFF_801.D ),
    .q(\DFF_801.Q )
  );
  al_dffl _9083_ (
    .clk(CK),
    .d(\DFF_802.D ),
    .q(\DFF_802.Q )
  );
  al_dffl _9084_ (
    .clk(CK),
    .d(\DFF_803.D ),
    .q(\DFF_803.Q )
  );
  al_dffl _9085_ (
    .clk(CK),
    .d(\DFF_807.D ),
    .q(\DFF_807.Q )
  );
  al_dffl _9086_ (
    .clk(CK),
    .d(\DFF_808.D ),
    .q(\DFF_808.Q )
  );
  al_dffl _9087_ (
    .clk(CK),
    .d(\DFF_809.D ),
    .q(\DFF_809.Q )
  );
  al_dffl _9088_ (
    .clk(CK),
    .d(\DFF_810.D ),
    .q(\DFF_810.Q )
  );
  al_dffl _9089_ (
    .clk(CK),
    .d(\DFF_811.D ),
    .q(\DFF_811.Q )
  );
  al_dffl _9090_ (
    .clk(CK),
    .d(\DFF_812.D ),
    .q(\DFF_812.Q )
  );
  al_dffl _9091_ (
    .clk(CK),
    .d(\DFF_813.D ),
    .q(\DFF_813.Q )
  );
  al_dffl _9092_ (
    .clk(CK),
    .d(\DFF_814.D ),
    .q(\DFF_814.Q )
  );
  al_dffl _9093_ (
    .clk(CK),
    .d(\DFF_815.D ),
    .q(\DFF_815.Q )
  );
  al_dffl _9094_ (
    .clk(CK),
    .d(\DFF_816.D ),
    .q(\DFF_816.Q )
  );
  al_dffl _9095_ (
    .clk(CK),
    .d(\DFF_817.D ),
    .q(\DFF_817.Q )
  );
  al_dffl _9096_ (
    .clk(CK),
    .d(\DFF_818.D ),
    .q(\DFF_818.Q )
  );
  al_dffl _9097_ (
    .clk(CK),
    .d(\DFF_819.D ),
    .q(\DFF_819.Q )
  );
  al_dffl _9098_ (
    .clk(CK),
    .d(\DFF_820.D ),
    .q(\DFF_820.Q )
  );
  al_dffl _9099_ (
    .clk(CK),
    .d(\DFF_821.D ),
    .q(\DFF_821.Q )
  );
  al_dffl _9100_ (
    .clk(CK),
    .d(\DFF_822.D ),
    .q(\DFF_822.Q )
  );
  al_dffl _9101_ (
    .clk(CK),
    .d(\DFF_823.D ),
    .q(\DFF_823.Q )
  );
  al_dffl _9102_ (
    .clk(CK),
    .d(\DFF_824.D ),
    .q(\DFF_824.Q )
  );
  al_dffl _9103_ (
    .clk(CK),
    .d(\DFF_825.D ),
    .q(\DFF_825.Q )
  );
  al_dffl _9104_ (
    .clk(CK),
    .d(\DFF_826.D ),
    .q(\DFF_826.Q )
  );
  al_dffl _9105_ (
    .clk(CK),
    .d(\DFF_827.D ),
    .q(\DFF_827.Q )
  );
  al_dffl _9106_ (
    .clk(CK),
    .d(\DFF_828.D ),
    .q(\DFF_828.Q )
  );
  al_dffl _9107_ (
    .clk(CK),
    .d(\DFF_829.D ),
    .q(\DFF_829.Q )
  );
  al_dffl _9108_ (
    .clk(CK),
    .d(\DFF_830.D ),
    .q(\DFF_830.Q )
  );
  al_dffl _9109_ (
    .clk(CK),
    .d(\DFF_831.D ),
    .q(\DFF_831.Q )
  );
  al_dffl _9110_ (
    .clk(CK),
    .d(\DFF_832.D ),
    .q(\DFF_832.Q )
  );
  al_dffl _9111_ (
    .clk(CK),
    .d(\DFF_833.D ),
    .q(\DFF_833.Q )
  );
  al_dffl _9112_ (
    .clk(CK),
    .d(\DFF_834.D ),
    .q(\DFF_834.Q )
  );
  al_dffl _9113_ (
    .clk(CK),
    .d(\DFF_835.D ),
    .q(\DFF_835.Q )
  );
  al_dffl _9114_ (
    .clk(CK),
    .d(\DFF_836.D ),
    .q(\DFF_836.Q )
  );
  al_dffl _9115_ (
    .clk(CK),
    .d(\DFF_837.D ),
    .q(\DFF_837.Q )
  );
  al_dffl _9116_ (
    .clk(CK),
    .d(\DFF_838.D ),
    .q(\DFF_838.Q )
  );
  al_dffl _9117_ (
    .clk(CK),
    .d(\DFF_839.D ),
    .q(\DFF_839.Q )
  );
  al_dffl _9118_ (
    .clk(CK),
    .d(\DFF_840.D ),
    .q(\DFF_840.Q )
  );
  al_dffl _9119_ (
    .clk(CK),
    .d(\DFF_841.D ),
    .q(\DFF_841.Q )
  );
  al_dffl _9120_ (
    .clk(CK),
    .d(\DFF_842.D ),
    .q(\DFF_842.Q )
  );
  al_dffl _9121_ (
    .clk(CK),
    .d(\DFF_843.D ),
    .q(\DFF_843.Q )
  );
  al_dffl _9122_ (
    .clk(CK),
    .d(\DFF_844.D ),
    .q(\DFF_844.Q )
  );
  al_dffl _9123_ (
    .clk(CK),
    .d(\DFF_845.D ),
    .q(\DFF_845.Q )
  );
  al_dffl _9124_ (
    .clk(CK),
    .d(\DFF_846.D ),
    .q(\DFF_846.Q )
  );
  al_dffl _9125_ (
    .clk(CK),
    .d(\DFF_847.D ),
    .q(\DFF_847.Q )
  );
  al_dffl _9126_ (
    .clk(CK),
    .d(\DFF_848.D ),
    .q(\DFF_848.Q )
  );
  al_dffl _9127_ (
    .clk(CK),
    .d(\DFF_849.D ),
    .q(\DFF_849.Q )
  );
  al_dffl _9128_ (
    .clk(CK),
    .d(\DFF_850.D ),
    .q(\DFF_850.Q )
  );
  al_dffl _9129_ (
    .clk(CK),
    .d(\DFF_851.D ),
    .q(\DFF_851.Q )
  );
  al_dffl _9130_ (
    .clk(CK),
    .d(\DFF_852.D ),
    .q(\DFF_852.Q )
  );
  al_dffl _9131_ (
    .clk(CK),
    .d(\DFF_853.D ),
    .q(\DFF_853.Q )
  );
  al_dffl _9132_ (
    .clk(CK),
    .d(\DFF_854.D ),
    .q(\DFF_854.Q )
  );
  al_dffl _9133_ (
    .clk(CK),
    .d(\DFF_855.D ),
    .q(\DFF_855.Q )
  );
  al_dffl _9134_ (
    .clk(CK),
    .d(\DFF_856.D ),
    .q(\DFF_856.Q )
  );
  al_dffl _9135_ (
    .clk(CK),
    .d(\DFF_857.D ),
    .q(\DFF_857.Q )
  );
  al_dffl _9136_ (
    .clk(CK),
    .d(\DFF_858.D ),
    .q(\DFF_858.Q )
  );
  al_dffl _9137_ (
    .clk(CK),
    .d(\DFF_859.D ),
    .q(\DFF_859.Q )
  );
  al_dffl _9138_ (
    .clk(CK),
    .d(\DFF_860.D ),
    .q(\DFF_860.Q )
  );
  al_dffl _9139_ (
    .clk(CK),
    .d(\DFF_864.D ),
    .q(\DFF_864.Q )
  );
  al_dffl _9140_ (
    .clk(CK),
    .d(\DFF_865.D ),
    .q(\DFF_865.Q )
  );
  al_dffl _9141_ (
    .clk(CK),
    .d(\DFF_866.D ),
    .q(\DFF_866.Q )
  );
  al_dffl _9142_ (
    .clk(CK),
    .d(\DFF_867.D ),
    .q(\DFF_867.Q )
  );
  al_dffl _9143_ (
    .clk(CK),
    .d(\DFF_868.D ),
    .q(\DFF_868.Q )
  );
  al_dffl _9144_ (
    .clk(CK),
    .d(\DFF_869.D ),
    .q(\DFF_869.Q )
  );
  al_dffl _9145_ (
    .clk(CK),
    .d(\DFF_870.D ),
    .q(\DFF_870.Q )
  );
  al_dffl _9146_ (
    .clk(CK),
    .d(\DFF_871.D ),
    .q(\DFF_871.Q )
  );
  al_dffl _9147_ (
    .clk(CK),
    .d(\DFF_872.D ),
    .q(\DFF_872.Q )
  );
  al_dffl _9148_ (
    .clk(CK),
    .d(\DFF_873.D ),
    .q(\DFF_873.Q )
  );
  al_dffl _9149_ (
    .clk(CK),
    .d(\DFF_874.D ),
    .q(\DFF_874.Q )
  );
  al_dffl _9150_ (
    .clk(CK),
    .d(\DFF_875.D ),
    .q(\DFF_875.Q )
  );
  al_dffl _9151_ (
    .clk(CK),
    .d(\DFF_876.D ),
    .q(\DFF_876.Q )
  );
  al_dffl _9152_ (
    .clk(CK),
    .d(\DFF_877.D ),
    .q(\DFF_877.Q )
  );
  al_dffl _9153_ (
    .clk(CK),
    .d(\DFF_878.D ),
    .q(\DFF_878.Q )
  );
  al_dffl _9154_ (
    .clk(CK),
    .d(\DFF_879.D ),
    .q(\DFF_879.Q )
  );
  al_dffl _9155_ (
    .clk(CK),
    .d(\DFF_880.D ),
    .q(\DFF_880.Q )
  );
  al_dffl _9156_ (
    .clk(CK),
    .d(\DFF_881.D ),
    .q(\DFF_881.Q )
  );
  al_dffl _9157_ (
    .clk(CK),
    .d(\DFF_882.D ),
    .q(\DFF_882.Q )
  );
  al_dffl _9158_ (
    .clk(CK),
    .d(\DFF_883.D ),
    .q(\DFF_883.Q )
  );
  al_dffl _9159_ (
    .clk(CK),
    .d(\DFF_884.D ),
    .q(\DFF_884.Q )
  );
  al_dffl _9160_ (
    .clk(CK),
    .d(\DFF_885.D ),
    .q(\DFF_885.Q )
  );
  al_dffl _9161_ (
    .clk(CK),
    .d(\DFF_886.D ),
    .q(\DFF_886.Q )
  );
  al_dffl _9162_ (
    .clk(CK),
    .d(\DFF_887.D ),
    .q(\DFF_887.Q )
  );
  al_dffl _9163_ (
    .clk(CK),
    .d(\DFF_888.D ),
    .q(\DFF_888.Q )
  );
  al_dffl _9164_ (
    .clk(CK),
    .d(\DFF_889.D ),
    .q(\DFF_889.Q )
  );
  al_dffl _9165_ (
    .clk(CK),
    .d(\DFF_890.D ),
    .q(\DFF_890.Q )
  );
  al_dffl _9166_ (
    .clk(CK),
    .d(\DFF_891.D ),
    .q(\DFF_891.Q )
  );
  al_dffl _9167_ (
    .clk(CK),
    .d(\DFF_892.D ),
    .q(\DFF_892.Q )
  );
  al_dffl _9168_ (
    .clk(CK),
    .d(\DFF_893.D ),
    .q(\DFF_893.Q )
  );
  al_dffl _9169_ (
    .clk(CK),
    .d(\DFF_894.D ),
    .q(\DFF_894.Q )
  );
  al_dffl _9170_ (
    .clk(CK),
    .d(\DFF_895.D ),
    .q(\DFF_895.Q )
  );
  al_dffl _9171_ (
    .clk(CK),
    .d(\DFF_896.D ),
    .q(\DFF_896.Q )
  );
  al_dffl _9172_ (
    .clk(CK),
    .d(\DFF_897.D ),
    .q(\DFF_897.Q )
  );
  al_dffl _9173_ (
    .clk(CK),
    .d(\DFF_898.D ),
    .q(\DFF_898.Q )
  );
  al_dffl _9174_ (
    .clk(CK),
    .d(\DFF_899.D ),
    .q(\DFF_899.Q )
  );
  al_dffl _9175_ (
    .clk(CK),
    .d(\DFF_900.D ),
    .q(\DFF_900.Q )
  );
  al_dffl _9176_ (
    .clk(CK),
    .d(\DFF_901.D ),
    .q(\DFF_901.Q )
  );
  al_dffl _9177_ (
    .clk(CK),
    .d(\DFF_902.D ),
    .q(\DFF_902.Q )
  );
  al_dffl _9178_ (
    .clk(CK),
    .d(\DFF_903.D ),
    .q(\DFF_903.Q )
  );
  al_dffl _9179_ (
    .clk(CK),
    .d(\DFF_904.D ),
    .q(\DFF_904.Q )
  );
  al_dffl _9180_ (
    .clk(CK),
    .d(\DFF_905.D ),
    .q(\DFF_905.Q )
  );
  al_dffl _9181_ (
    .clk(CK),
    .d(\DFF_906.D ),
    .q(\DFF_906.Q )
  );
  al_dffl _9182_ (
    .clk(CK),
    .d(\DFF_907.D ),
    .q(\DFF_907.Q )
  );
  al_dffl _9183_ (
    .clk(CK),
    .d(\DFF_908.D ),
    .q(\DFF_908.Q )
  );
  al_dffl _9184_ (
    .clk(CK),
    .d(\DFF_909.D ),
    .q(\DFF_909.Q )
  );
  al_dffl _9185_ (
    .clk(CK),
    .d(\DFF_910.D ),
    .q(\DFF_910.Q )
  );
  al_dffl _9186_ (
    .clk(CK),
    .d(\DFF_911.D ),
    .q(\DFF_911.Q )
  );
  al_dffl _9187_ (
    .clk(CK),
    .d(\DFF_912.D ),
    .q(\DFF_912.Q )
  );
  al_dffl _9188_ (
    .clk(CK),
    .d(\DFF_913.D ),
    .q(\DFF_913.Q )
  );
  al_dffl _9189_ (
    .clk(CK),
    .d(\DFF_914.D ),
    .q(\DFF_914.Q )
  );
  al_dffl _9190_ (
    .clk(CK),
    .d(\DFF_915.D ),
    .q(\DFF_915.Q )
  );
  al_dffl _9191_ (
    .clk(CK),
    .d(\DFF_916.D ),
    .q(\DFF_916.Q )
  );
  al_dffl _9192_ (
    .clk(CK),
    .d(\DFF_917.D ),
    .q(\DFF_917.Q )
  );
  al_dffl _9193_ (
    .clk(CK),
    .d(\DFF_918.D ),
    .q(\DFF_918.Q )
  );
  al_dffl _9194_ (
    .clk(CK),
    .d(\DFF_919.D ),
    .q(\DFF_919.Q )
  );
  al_dffl _9195_ (
    .clk(CK),
    .d(\DFF_920.D ),
    .q(\DFF_920.Q )
  );
  al_dffl _9196_ (
    .clk(CK),
    .d(\DFF_921.D ),
    .q(\DFF_921.Q )
  );
  al_dffl _9197_ (
    .clk(CK),
    .d(\DFF_922.D ),
    .q(\DFF_922.Q )
  );
  al_dffl _9198_ (
    .clk(CK),
    .d(\DFF_923.D ),
    .q(\DFF_923.Q )
  );
  al_dffl _9199_ (
    .clk(CK),
    .d(\DFF_924.D ),
    .q(\DFF_924.Q )
  );
  al_dffl _9200_ (
    .clk(CK),
    .d(\DFF_925.D ),
    .q(\DFF_925.Q )
  );
  al_dffl _9201_ (
    .clk(CK),
    .d(\DFF_926.D ),
    .q(\DFF_926.Q )
  );
  al_dffl _9202_ (
    .clk(CK),
    .d(\DFF_927.D ),
    .q(\DFF_927.Q )
  );
  al_dffl _9203_ (
    .clk(CK),
    .d(\DFF_928.D ),
    .q(\DFF_928.Q )
  );
  al_dffl _9204_ (
    .clk(CK),
    .d(\DFF_929.D ),
    .q(\DFF_929.Q )
  );
  al_dffl _9205_ (
    .clk(CK),
    .d(\DFF_930.D ),
    .q(\DFF_930.Q )
  );
  al_dffl _9206_ (
    .clk(CK),
    .d(\DFF_931.D ),
    .q(\DFF_931.Q )
  );
  al_dffl _9207_ (
    .clk(CK),
    .d(\DFF_932.D ),
    .q(\DFF_932.Q )
  );
  al_dffl _9208_ (
    .clk(CK),
    .d(\DFF_933.D ),
    .q(\DFF_933.Q )
  );
  al_dffl _9209_ (
    .clk(CK),
    .d(\DFF_934.D ),
    .q(\DFF_934.Q )
  );
  al_dffl _9210_ (
    .clk(CK),
    .d(\DFF_935.D ),
    .q(\DFF_935.Q )
  );
  al_dffl _9211_ (
    .clk(CK),
    .d(\DFF_936.D ),
    .q(\DFF_936.Q )
  );
  al_dffl _9212_ (
    .clk(CK),
    .d(\DFF_937.D ),
    .q(\DFF_937.Q )
  );
  al_dffl _9213_ (
    .clk(CK),
    .d(\DFF_938.D ),
    .q(\DFF_938.Q )
  );
  al_dffl _9214_ (
    .clk(CK),
    .d(\DFF_939.D ),
    .q(\DFF_939.Q )
  );
  al_dffl _9215_ (
    .clk(CK),
    .d(\DFF_940.D ),
    .q(\DFF_940.Q )
  );
  al_dffl _9216_ (
    .clk(CK),
    .d(\DFF_941.D ),
    .q(\DFF_941.Q )
  );
  al_dffl _9217_ (
    .clk(CK),
    .d(\DFF_942.D ),
    .q(\DFF_942.Q )
  );
  al_dffl _9218_ (
    .clk(CK),
    .d(\DFF_943.D ),
    .q(\DFF_943.Q )
  );
  al_dffl _9219_ (
    .clk(CK),
    .d(\DFF_944.D ),
    .q(\DFF_944.Q )
  );
  al_dffl _9220_ (
    .clk(CK),
    .d(\DFF_945.D ),
    .q(\DFF_945.Q )
  );
  al_dffl _9221_ (
    .clk(CK),
    .d(\DFF_953.D ),
    .q(\DFF_953.Q )
  );
  al_dffl _9222_ (
    .clk(CK),
    .d(\DFF_954.D ),
    .q(\DFF_954.Q )
  );
  al_dffl _9223_ (
    .clk(CK),
    .d(\DFF_955.D ),
    .q(\DFF_955.Q )
  );
  al_dffl _9224_ (
    .clk(CK),
    .d(\DFF_956.D ),
    .q(\DFF_956.Q )
  );
  al_dffl _9225_ (
    .clk(CK),
    .d(\DFF_957.D ),
    .q(\DFF_957.Q )
  );
  al_dffl _9226_ (
    .clk(CK),
    .d(\DFF_958.D ),
    .q(\DFF_958.Q )
  );
  al_dffl _9227_ (
    .clk(CK),
    .d(\DFF_959.D ),
    .q(\DFF_959.Q )
  );
  al_dffl _9228_ (
    .clk(CK),
    .d(\DFF_960.D ),
    .q(\DFF_960.Q )
  );
  al_dffl _9229_ (
    .clk(CK),
    .d(\DFF_961.D ),
    .q(\DFF_961.Q )
  );
  al_dffl _9230_ (
    .clk(CK),
    .d(\DFF_962.D ),
    .q(\DFF_962.Q )
  );
  al_dffl _9231_ (
    .clk(CK),
    .d(\DFF_963.D ),
    .q(\DFF_963.Q )
  );
  al_dffl _9232_ (
    .clk(CK),
    .d(\DFF_964.D ),
    .q(\DFF_964.Q )
  );
  al_dffl _9233_ (
    .clk(CK),
    .d(\DFF_965.D ),
    .q(\DFF_965.Q )
  );
  al_dffl _9234_ (
    .clk(CK),
    .d(\DFF_966.D ),
    .q(\DFF_966.Q )
  );
  al_dffl _9235_ (
    .clk(CK),
    .d(\DFF_967.D ),
    .q(\DFF_967.Q )
  );
  al_dffl _9236_ (
    .clk(CK),
    .d(\DFF_968.D ),
    .q(\DFF_968.Q )
  );
  al_dffl _9237_ (
    .clk(CK),
    .d(\DFF_969.D ),
    .q(\DFF_969.Q )
  );
  al_dffl _9238_ (
    .clk(CK),
    .d(\DFF_970.D ),
    .q(\DFF_970.Q )
  );
  al_dffl _9239_ (
    .clk(CK),
    .d(\DFF_971.D ),
    .q(\DFF_971.Q )
  );
  al_dffl _9240_ (
    .clk(CK),
    .d(\DFF_972.D ),
    .q(\DFF_972.Q )
  );
  al_dffl _9241_ (
    .clk(CK),
    .d(\DFF_973.D ),
    .q(\DFF_973.Q )
  );
  al_dffl _9242_ (
    .clk(CK),
    .d(\DFF_974.D ),
    .q(\DFF_974.Q )
  );
  al_dffl _9243_ (
    .clk(CK),
    .d(\DFF_975.D ),
    .q(\DFF_975.Q )
  );
  al_dffl _9244_ (
    .clk(CK),
    .d(\DFF_976.D ),
    .q(\DFF_976.Q )
  );
  al_dffl _9245_ (
    .clk(CK),
    .d(\DFF_977.D ),
    .q(\DFF_977.Q )
  );
  al_dffl _9246_ (
    .clk(CK),
    .d(\DFF_978.D ),
    .q(\DFF_978.Q )
  );
  al_dffl _9247_ (
    .clk(CK),
    .d(\DFF_979.D ),
    .q(\DFF_979.Q )
  );
  al_dffl _9248_ (
    .clk(CK),
    .d(\DFF_980.D ),
    .q(\DFF_980.Q )
  );
  al_dffl _9249_ (
    .clk(CK),
    .d(\DFF_981.D ),
    .q(\DFF_981.Q )
  );
  al_dffl _9250_ (
    .clk(CK),
    .d(\DFF_982.D ),
    .q(\DFF_982.Q )
  );
  al_dffl _9251_ (
    .clk(CK),
    .d(\DFF_983.D ),
    .q(\DFF_983.Q )
  );
  al_dffl _9252_ (
    .clk(CK),
    .d(\DFF_984.D ),
    .q(\DFF_984.Q )
  );
  al_dffl _9253_ (
    .clk(CK),
    .d(\DFF_985.D ),
    .q(\DFF_985.Q )
  );
  al_dffl _9254_ (
    .clk(CK),
    .d(\DFF_986.D ),
    .q(\DFF_986.Q )
  );
  al_dffl _9255_ (
    .clk(CK),
    .d(\DFF_987.D ),
    .q(\DFF_987.Q )
  );
  al_dffl _9256_ (
    .clk(CK),
    .d(\DFF_988.D ),
    .q(\DFF_988.Q )
  );
  al_dffl _9257_ (
    .clk(CK),
    .d(\DFF_989.D ),
    .q(\DFF_989.Q )
  );
  al_dffl _9258_ (
    .clk(CK),
    .d(\DFF_990.D ),
    .q(\DFF_990.Q )
  );
  al_dffl _9259_ (
    .clk(CK),
    .d(\DFF_991.D ),
    .q(\DFF_991.Q )
  );
  al_dffl _9260_ (
    .clk(CK),
    .d(\DFF_992.D ),
    .q(\DFF_992.Q )
  );
  al_dffl _9261_ (
    .clk(CK),
    .d(\DFF_993.D ),
    .q(\DFF_993.Q )
  );
  al_dffl _9262_ (
    .clk(CK),
    .d(\DFF_994.D ),
    .q(\DFF_994.Q )
  );
  al_dffl _9263_ (
    .clk(CK),
    .d(\DFF_995.D ),
    .q(\DFF_995.Q )
  );
  al_dffl _9264_ (
    .clk(CK),
    .d(\DFF_996.D ),
    .q(\DFF_996.Q )
  );
  al_dffl _9265_ (
    .clk(CK),
    .d(\DFF_997.D ),
    .q(\DFF_997.Q )
  );
  al_dffl _9266_ (
    .clk(CK),
    .d(\DFF_998.D ),
    .q(\DFF_998.Q )
  );
  al_dffl _9267_ (
    .clk(CK),
    .d(\DFF_998.Q ),
    .q(\DFF_999.Q )
  );
  al_dffl _9268_ (
    .clk(CK),
    .d(\DFF_1000.D ),
    .q(\DFF_1000.Q )
  );
  al_dffl _9269_ (
    .clk(CK),
    .d(\DFF_1000.Q ),
    .q(\DFF_1001.Q )
  );
  al_dffl _9270_ (
    .clk(CK),
    .d(\DFF_1002.D ),
    .q(\DFF_1002.Q )
  );
  al_dffl _9271_ (
    .clk(CK),
    .d(\DFF_1002.Q ),
    .q(\DFF_1003.Q )
  );
  al_dffl _9272_ (
    .clk(CK),
    .d(\DFF_1004.D ),
    .q(\DFF_1004.Q )
  );
  al_dffl _9273_ (
    .clk(CK),
    .d(\DFF_1004.Q ),
    .q(\DFF_1005.Q )
  );
  al_dffl _9274_ (
    .clk(CK),
    .d(\DFF_1006.D ),
    .q(\DFF_1006.Q )
  );
  al_dffl _9275_ (
    .clk(CK),
    .d(\DFF_1006.Q ),
    .q(\DFF_1007.Q )
  );
  al_dffl _9276_ (
    .clk(CK),
    .d(\DFF_1008.D ),
    .q(\DFF_1008.Q )
  );
  al_dffl _9277_ (
    .clk(CK),
    .d(\DFF_1008.Q ),
    .q(\DFF_1009.Q )
  );
  al_dffl _9278_ (
    .clk(CK),
    .d(\DFF_1010.D ),
    .q(\DFF_1010.Q )
  );
  al_dffl _9279_ (
    .clk(CK),
    .d(\DFF_1010.Q ),
    .q(\DFF_1011.Q )
  );
  al_dffl _9280_ (
    .clk(CK),
    .d(\DFF_1012.D ),
    .q(\DFF_1012.Q )
  );
  al_dffl _9281_ (
    .clk(CK),
    .d(\DFF_1012.Q ),
    .q(\DFF_1013.Q )
  );
  al_dffl _9282_ (
    .clk(CK),
    .d(\DFF_46.Q ),
    .q(\DFF_1014.Q )
  );
  al_dffl _9283_ (
    .clk(CK),
    .d(\DFF_1014.Q ),
    .q(\DFF_1015.Q )
  );
  al_dffl _9284_ (
    .clk(CK),
    .d(\DFF_1016.D ),
    .q(\DFF_1016.Q )
  );
  al_dffl _9285_ (
    .clk(CK),
    .d(\DFF_1017.D ),
    .q(\DFF_1017.Q )
  );
  al_dffl _9286_ (
    .clk(CK),
    .d(\DFF_1028.D ),
    .q(\DFF_1028.Q )
  );
  al_dffl _9287_ (
    .clk(CK),
    .d(\DFF_953.Q ),
    .q(\DFF_1029.Q )
  );
  al_dffl _9288_ (
    .clk(CK),
    .d(\DFF_1029.Q ),
    .q(\DFF_1030.Q )
  );
  al_dffl _9289_ (
    .clk(CK),
    .d(\DFF_954.Q ),
    .q(\DFF_1031.Q )
  );
  al_dffl _9290_ (
    .clk(CK),
    .d(\DFF_1031.Q ),
    .q(\DFF_1032.Q )
  );
  al_dffl _9291_ (
    .clk(CK),
    .d(\DFF_955.Q ),
    .q(\DFF_1033.Q )
  );
  al_dffl _9292_ (
    .clk(CK),
    .d(\DFF_1033.Q ),
    .q(\DFF_1034.Q )
  );
  al_dffl _9293_ (
    .clk(CK),
    .d(\DFF_956.Q ),
    .q(\DFF_1035.Q )
  );
  al_dffl _9294_ (
    .clk(CK),
    .d(\DFF_1035.Q ),
    .q(\DFF_1036.Q )
  );
  al_dffl _9295_ (
    .clk(CK),
    .d(\DFF_957.Q ),
    .q(\DFF_1037.Q )
  );
  al_dffl _9296_ (
    .clk(CK),
    .d(\DFF_1037.Q ),
    .q(\DFF_1038.Q )
  );
  al_dffl _9297_ (
    .clk(CK),
    .d(\DFF_958.Q ),
    .q(\DFF_1039.Q )
  );
  al_dffl _9298_ (
    .clk(CK),
    .d(\DFF_1039.Q ),
    .q(\DFF_1040.Q )
  );
  al_dffl _9299_ (
    .clk(CK),
    .d(\DFF_959.Q ),
    .q(\DFF_1041.Q )
  );
  al_dffl _9300_ (
    .clk(CK),
    .d(\DFF_1041.Q ),
    .q(\DFF_1042.Q )
  );
  al_dffl _9301_ (
    .clk(CK),
    .d(\DFF_960.Q ),
    .q(\DFF_1043.Q )
  );
  al_dffl _9302_ (
    .clk(CK),
    .d(\DFF_1043.Q ),
    .q(\DFF_1044.Q )
  );
  al_dffl _9303_ (
    .clk(CK),
    .d(\DFF_961.Q ),
    .q(\DFF_1045.Q )
  );
  al_dffl _9304_ (
    .clk(CK),
    .d(\DFF_1045.Q ),
    .q(\DFF_1046.Q )
  );
  al_dffl _9305_ (
    .clk(CK),
    .d(\DFF_962.Q ),
    .q(\DFF_1047.Q )
  );
  al_dffl _9306_ (
    .clk(CK),
    .d(\DFF_1047.Q ),
    .q(\DFF_1048.Q )
  );
  al_dffl _9307_ (
    .clk(CK),
    .d(\DFF_963.Q ),
    .q(\DFF_1049.Q )
  );
  al_dffl _9308_ (
    .clk(CK),
    .d(\DFF_1049.Q ),
    .q(\DFF_1050.Q )
  );
  al_dffl _9309_ (
    .clk(CK),
    .d(\DFF_964.Q ),
    .q(\DFF_1051.Q )
  );
  al_dffl _9310_ (
    .clk(CK),
    .d(\DFF_1051.Q ),
    .q(\DFF_1052.Q )
  );
  al_dffl _9311_ (
    .clk(CK),
    .d(\DFF_1059.D ),
    .q(\DFF_1059.Q )
  );
  al_dffl _9312_ (
    .clk(CK),
    .d(\DFF_1060.D ),
    .q(\DFF_1060.Q )
  );
  al_dffl _9313_ (
    .clk(CK),
    .d(\DFF_1061.D ),
    .q(\DFF_1061.Q )
  );
  al_dffl _9314_ (
    .clk(CK),
    .d(\DFF_1062.D ),
    .q(\DFF_1062.Q )
  );
  al_dffl _9315_ (
    .clk(CK),
    .d(\DFF_1062.Q ),
    .q(\DFF_1063.Q )
  );
  al_dffl _9316_ (
    .clk(CK),
    .d(\DFF_1063.Q ),
    .q(\DFF_1064.Q )
  );
  al_dffl _9317_ (
    .clk(CK),
    .d(\DFF_1083.Q ),
    .q(\DFF_1065.Q )
  );
  al_dffl _9318_ (
    .clk(CK),
    .d(\DFF_1065.Q ),
    .q(\DFF_1066.Q )
  );
  al_dffl _9319_ (
    .clk(CK),
    .d(\DFF_1084.Q ),
    .q(\DFF_1067.Q )
  );
  al_dffl _9320_ (
    .clk(CK),
    .d(\DFF_1067.Q ),
    .q(\DFF_1068.Q )
  );
  al_dffl _9321_ (
    .clk(CK),
    .d(\DFF_1085.Q ),
    .q(\DFF_1069.Q )
  );
  al_dffl _9322_ (
    .clk(CK),
    .d(\DFF_1069.Q ),
    .q(\DFF_1070.Q )
  );
  al_dffl _9323_ (
    .clk(CK),
    .d(\DFF_1092.Q ),
    .q(\DFF_1071.Q )
  );
  al_dffl _9324_ (
    .clk(CK),
    .d(\DFF_1071.Q ),
    .q(\DFF_1072.Q )
  );
  al_dffl _9325_ (
    .clk(CK),
    .d(\DFF_1093.Q ),
    .q(\DFF_1073.Q )
  );
  al_dffl _9326_ (
    .clk(CK),
    .d(\DFF_1073.Q ),
    .q(\DFF_1074.Q )
  );
  al_dffl _9327_ (
    .clk(CK),
    .d(\DFF_1094.Q ),
    .q(\DFF_1075.Q )
  );
  al_dffl _9328_ (
    .clk(CK),
    .d(\DFF_1075.Q ),
    .q(\DFF_1076.Q )
  );
  al_dffl _9329_ (
    .clk(CK),
    .d(\DFF_1080.D ),
    .q(\DFF_1080.Q )
  );
  al_dffl _9330_ (
    .clk(CK),
    .d(\DFF_1081.D ),
    .q(\DFF_1081.Q )
  );
  al_dffl _9331_ (
    .clk(CK),
    .d(\DFF_1082.D ),
    .q(\DFF_1082.Q )
  );
  al_dffl _9332_ (
    .clk(CK),
    .d(\DFF_1083.D ),
    .q(\DFF_1083.Q )
  );
  al_dffl _9333_ (
    .clk(CK),
    .d(\DFF_1084.D ),
    .q(\DFF_1084.Q )
  );
  al_dffl _9334_ (
    .clk(CK),
    .d(\DFF_1085.D ),
    .q(\DFF_1085.Q )
  );
  al_dffl _9335_ (
    .clk(CK),
    .d(\DFF_1086.D ),
    .q(\DFF_1086.Q )
  );
  al_dffl _9336_ (
    .clk(CK),
    .d(\DFF_1087.D ),
    .q(\DFF_1087.Q )
  );
  al_dffl _9337_ (
    .clk(CK),
    .d(\DFF_1088.D ),
    .q(\DFF_1088.Q )
  );
  al_dffl _9338_ (
    .clk(CK),
    .d(\DFF_1089.D ),
    .q(\DFF_1089.Q )
  );
  al_dffl _9339_ (
    .clk(CK),
    .d(\DFF_1090.D ),
    .q(\DFF_1090.Q )
  );
  al_dffl _9340_ (
    .clk(CK),
    .d(\DFF_1091.D ),
    .q(\DFF_1091.Q )
  );
  al_dffl _9341_ (
    .clk(CK),
    .d(\DFF_1092.D ),
    .q(\DFF_1092.Q )
  );
  al_dffl _9342_ (
    .clk(CK),
    .d(\DFF_1093.D ),
    .q(\DFF_1093.Q )
  );
  al_dffl _9343_ (
    .clk(CK),
    .d(\DFF_1094.D ),
    .q(\DFF_1094.Q )
  );
  al_dffl _9344_ (
    .clk(CK),
    .d(\DFF_1095.D ),
    .q(\DFF_1095.Q )
  );
  al_dffl _9345_ (
    .clk(CK),
    .d(\DFF_1095.Q ),
    .q(\DFF_1096.Q )
  );
  al_dffl _9346_ (
    .clk(CK),
    .d(\DFF_1096.Q ),
    .q(\DFF_1097.Q )
  );
  al_dffl _9347_ (
    .clk(CK),
    .d(\DFF_1098.D ),
    .q(\DFF_1098.Q )
  );
  al_dffl _9348_ (
    .clk(CK),
    .d(\DFF_1098.Q ),
    .q(\DFF_1099.Q )
  );
  al_dffl _9349_ (
    .clk(CK),
    .d(\DFF_1100.D ),
    .q(\DFF_1100.Q )
  );
  al_dffl _9350_ (
    .clk(CK),
    .d(\DFF_1101.D ),
    .q(\DFF_1101.Q )
  );
  al_dffl _9351_ (
    .clk(CK),
    .d(\DFF_1101.Q ),
    .q(\DFF_1102.Q )
  );
  al_dffl _9352_ (
    .clk(CK),
    .d(\DFF_1103.D ),
    .q(\DFF_1103.Q )
  );
  al_dffl _9353_ (
    .clk(CK),
    .d(\DFF_1103.Q ),
    .q(\DFF_1104.Q )
  );
  al_dffl _9354_ (
    .clk(CK),
    .d(\DFF_1105.D ),
    .q(\DFF_1105.Q )
  );
  al_dffl _9355_ (
    .clk(CK),
    .d(\DFF_1106.D ),
    .q(\DFF_1106.Q )
  );
  al_dffl _9356_ (
    .clk(CK),
    .d(\DFF_1107.D ),
    .q(\DFF_1107.Q )
  );
  al_dffl _9357_ (
    .clk(CK),
    .d(\DFF_1108.D ),
    .q(\DFF_1108.Q )
  );
  al_dffl _9358_ (
    .clk(CK),
    .d(\DFF_1109.D ),
    .q(\DFF_1109.Q )
  );
  al_dffl _9359_ (
    .clk(CK),
    .d(\DFF_1110.D ),
    .q(\DFF_1110.Q )
  );
  al_dffl _9360_ (
    .clk(CK),
    .d(\DFF_1111.D ),
    .q(\DFF_1111.Q )
  );
  al_dffl _9361_ (
    .clk(CK),
    .d(\DFF_1112.D ),
    .q(\DFF_1112.Q )
  );
  al_dffl _9362_ (
    .clk(CK),
    .d(\DFF_1113.D ),
    .q(\DFF_1113.Q )
  );
  al_dffl _9363_ (
    .clk(CK),
    .d(\DFF_1114.D ),
    .q(\DFF_1114.Q )
  );
  al_dffl _9364_ (
    .clk(CK),
    .d(\DFF_1115.D ),
    .q(\DFF_1115.Q )
  );
  al_dffl _9365_ (
    .clk(CK),
    .d(\DFF_1116.D ),
    .q(\DFF_1116.Q )
  );
  al_dffl _9366_ (
    .clk(CK),
    .d(\DFF_1117.D ),
    .q(\DFF_1117.Q )
  );
  al_dffl _9367_ (
    .clk(CK),
    .d(\DFF_1118.D ),
    .q(\DFF_1118.Q )
  );
  al_dffl _9368_ (
    .clk(CK),
    .d(\DFF_1119.D ),
    .q(\DFF_1119.Q )
  );
  al_dffl _9369_ (
    .clk(CK),
    .d(\DFF_1120.D ),
    .q(\DFF_1120.Q )
  );
  al_dffl _9370_ (
    .clk(CK),
    .d(\DFF_1121.D ),
    .q(\DFF_1121.Q )
  );
  al_dffl _9371_ (
    .clk(CK),
    .d(\DFF_1122.D ),
    .q(\DFF_1122.Q )
  );
  al_dffl _9372_ (
    .clk(CK),
    .d(\DFF_1123.D ),
    .q(\DFF_1123.Q )
  );
  al_dffl _9373_ (
    .clk(CK),
    .d(\DFF_1124.D ),
    .q(\DFF_1124.Q )
  );
  al_dffl _9374_ (
    .clk(CK),
    .d(\DFF_1125.D ),
    .q(\DFF_1125.Q )
  );
  al_dffl _9375_ (
    .clk(CK),
    .d(\DFF_1126.D ),
    .q(\DFF_1126.Q )
  );
  al_dffl _9376_ (
    .clk(CK),
    .d(\DFF_1127.D ),
    .q(\DFF_1127.Q )
  );
  al_dffl _9377_ (
    .clk(CK),
    .d(\DFF_1128.D ),
    .q(\DFF_1128.Q )
  );
  al_dffl _9378_ (
    .clk(CK),
    .d(\DFF_1129.D ),
    .q(\DFF_1129.Q )
  );
  al_dffl _9379_ (
    .clk(CK),
    .d(\DFF_1130.D ),
    .q(\DFF_1130.Q )
  );
  al_dffl _9380_ (
    .clk(CK),
    .d(\DFF_1131.D ),
    .q(\DFF_1131.Q )
  );
  al_dffl _9381_ (
    .clk(CK),
    .d(\DFF_1102.Q ),
    .q(\DFF_1132.Q )
  );
  al_dffl _9382_ (
    .clk(CK),
    .d(\DFF_1133.D ),
    .q(\DFF_1133.Q )
  );
  al_dffl _9383_ (
    .clk(CK),
    .d(\DFF_1142.D ),
    .q(\DFF_1142.Q )
  );
  al_dffl _9384_ (
    .clk(CK),
    .d(\DFF_1142.Q ),
    .q(\DFF_1143.Q )
  );
  al_dffl _9385_ (
    .clk(CK),
    .d(\DFF_1144.D ),
    .q(\DFF_1144.Q )
  );
  al_dffl _9386_ (
    .clk(CK),
    .d(\DFF_1145.D ),
    .q(\DFF_1145.Q )
  );
  al_dffl _9387_ (
    .clk(CK),
    .d(\DFF_1146.D ),
    .q(\DFF_1146.Q )
  );
  al_dffl _9388_ (
    .clk(CK),
    .d(\DFF_1147.D ),
    .q(\DFF_1147.Q )
  );
  al_dffl _9389_ (
    .clk(CK),
    .d(\DFF_1148.D ),
    .q(\DFF_1148.Q )
  );
  al_dffl _9390_ (
    .clk(CK),
    .d(\DFF_1149.D ),
    .q(\DFF_1149.Q )
  );
  al_dffl _9391_ (
    .clk(CK),
    .d(\DFF_1150.D ),
    .q(\DFF_1150.Q )
  );
  al_dffl _9392_ (
    .clk(CK),
    .d(\DFF_1151.D ),
    .q(\DFF_1151.Q )
  );
  al_dffl _9393_ (
    .clk(CK),
    .d(\DFF_1152.D ),
    .q(\DFF_1152.Q )
  );
  al_dffl _9394_ (
    .clk(CK),
    .d(\DFF_1153.D ),
    .q(\DFF_1153.Q )
  );
  al_dffl _9395_ (
    .clk(CK),
    .d(\DFF_1157.D ),
    .q(\DFF_1157.Q )
  );
  al_dffl _9396_ (
    .clk(CK),
    .d(\DFF_1158.D ),
    .q(\DFF_1158.Q )
  );
  al_dffl _9397_ (
    .clk(CK),
    .d(\DFF_1159.D ),
    .q(\DFF_1159.Q )
  );
  al_dffl _9398_ (
    .clk(CK),
    .d(\DFF_1160.D ),
    .q(\DFF_1160.Q )
  );
  al_dffl _9399_ (
    .clk(CK),
    .d(\DFF_1161.D ),
    .q(\DFF_1161.Q )
  );
  al_dffl _9400_ (
    .clk(CK),
    .d(\DFF_1162.D ),
    .q(\DFF_1162.Q )
  );
  al_dffl _9401_ (
    .clk(CK),
    .d(\DFF_1163.D ),
    .q(\DFF_1163.Q )
  );
  al_dffl _9402_ (
    .clk(CK),
    .d(\DFF_1164.D ),
    .q(\DFF_1164.Q )
  );
  al_dffl _9403_ (
    .clk(CK),
    .d(\DFF_1165.D ),
    .q(\DFF_1165.Q )
  );
  al_dffl _9404_ (
    .clk(CK),
    .d(\DFF_1166.D ),
    .q(\DFF_1166.Q )
  );
  al_dffl _9405_ (
    .clk(CK),
    .d(\DFF_1167.D ),
    .q(\DFF_1167.Q )
  );
  al_dffl _9406_ (
    .clk(CK),
    .d(\DFF_1168.D ),
    .q(\DFF_1168.Q )
  );
  al_dffl _9407_ (
    .clk(CK),
    .d(\DFF_1169.D ),
    .q(\DFF_1169.Q )
  );
  al_dffl _9408_ (
    .clk(CK),
    .d(\DFF_1170.D ),
    .q(\DFF_1170.Q )
  );
  al_dffl _9409_ (
    .clk(CK),
    .d(\DFF_1171.D ),
    .q(\DFF_1171.Q )
  );
  al_dffl _9410_ (
    .clk(CK),
    .d(\DFF_1172.D ),
    .q(\DFF_1172.Q )
  );
  al_dffl _9411_ (
    .clk(CK),
    .d(\DFF_1173.D ),
    .q(\DFF_1173.Q )
  );
  al_dffl _9412_ (
    .clk(CK),
    .d(\DFF_1174.D ),
    .q(\DFF_1174.Q )
  );
  al_dffl _9413_ (
    .clk(CK),
    .d(\DFF_1175.D ),
    .q(\DFF_1175.Q )
  );
  al_dffl _9414_ (
    .clk(CK),
    .d(\DFF_1176.D ),
    .q(\DFF_1176.Q )
  );
  al_dffl _9415_ (
    .clk(CK),
    .d(\DFF_1177.D ),
    .q(\DFF_1177.Q )
  );
  al_dffl _9416_ (
    .clk(CK),
    .d(\DFF_1178.D ),
    .q(\DFF_1178.Q )
  );
  al_dffl _9417_ (
    .clk(CK),
    .d(\DFF_1179.D ),
    .q(\DFF_1179.Q )
  );
  al_dffl _9418_ (
    .clk(CK),
    .d(\DFF_1180.D ),
    .q(\DFF_1180.Q )
  );
  al_dffl _9419_ (
    .clk(CK),
    .d(\DFF_1181.D ),
    .q(\DFF_1181.Q )
  );
  al_dffl _9420_ (
    .clk(CK),
    .d(\DFF_1182.D ),
    .q(\DFF_1182.Q )
  );
  al_dffl _9421_ (
    .clk(CK),
    .d(\DFF_1183.D ),
    .q(\DFF_1183.Q )
  );
  al_dffl _9422_ (
    .clk(CK),
    .d(\DFF_1184.D ),
    .q(\DFF_1184.Q )
  );
  al_dffl _9423_ (
    .clk(CK),
    .d(\DFF_1185.D ),
    .q(\DFF_1185.Q )
  );
  al_dffl _9424_ (
    .clk(CK),
    .d(\DFF_1186.D ),
    .q(\DFF_1186.Q )
  );
  al_dffl _9425_ (
    .clk(CK),
    .d(\DFF_1187.D ),
    .q(\DFF_1187.Q )
  );
  al_dffl _9426_ (
    .clk(CK),
    .d(\DFF_1188.D ),
    .q(\DFF_1188.Q )
  );
  al_dffl _9427_ (
    .clk(CK),
    .d(\DFF_1189.D ),
    .q(\DFF_1189.Q )
  );
  al_dffl _9428_ (
    .clk(CK),
    .d(\DFF_1190.D ),
    .q(\DFF_1190.Q )
  );
  al_dffl _9429_ (
    .clk(CK),
    .d(\DFF_1191.D ),
    .q(\DFF_1191.Q )
  );
  al_dffl _9430_ (
    .clk(CK),
    .d(\DFF_1192.D ),
    .q(\DFF_1192.Q )
  );
  al_dffl _9431_ (
    .clk(CK),
    .d(\DFF_1193.D ),
    .q(\DFF_1193.Q )
  );
  al_dffl _9432_ (
    .clk(CK),
    .d(\DFF_1194.D ),
    .q(\DFF_1194.Q )
  );
  al_dffl _9433_ (
    .clk(CK),
    .d(\DFF_1195.D ),
    .q(\DFF_1195.Q )
  );
  al_dffl _9434_ (
    .clk(CK),
    .d(\DFF_1196.D ),
    .q(\DFF_1196.Q )
  );
  al_dffl _9435_ (
    .clk(CK),
    .d(\DFF_1197.D ),
    .q(\DFF_1197.Q )
  );
  al_dffl _9436_ (
    .clk(CK),
    .d(\DFF_1198.D ),
    .q(\DFF_1198.Q )
  );
  al_dffl _9437_ (
    .clk(CK),
    .d(\DFF_1199.D ),
    .q(\DFF_1199.Q )
  );
  al_dffl _9438_ (
    .clk(CK),
    .d(\DFF_1200.D ),
    .q(\DFF_1200.Q )
  );
  al_dffl _9439_ (
    .clk(CK),
    .d(\DFF_1201.D ),
    .q(\DFF_1201.Q )
  );
  al_dffl _9440_ (
    .clk(CK),
    .d(\DFF_1202.D ),
    .q(\DFF_1202.Q )
  );
  al_dffl _9441_ (
    .clk(CK),
    .d(\DFF_1203.D ),
    .q(\DFF_1203.Q )
  );
  al_dffl _9442_ (
    .clk(CK),
    .d(\DFF_1204.D ),
    .q(\DFF_1204.Q )
  );
  al_dffl _9443_ (
    .clk(CK),
    .d(\DFF_1205.D ),
    .q(\DFF_1205.Q )
  );
  al_dffl _9444_ (
    .clk(CK),
    .d(\DFF_1206.D ),
    .q(\DFF_1206.Q )
  );
  al_dffl _9445_ (
    .clk(CK),
    .d(\DFF_1207.D ),
    .q(\DFF_1207.Q )
  );
  al_dffl _9446_ (
    .clk(CK),
    .d(\DFF_1208.D ),
    .q(\DFF_1208.Q )
  );
  al_dffl _9447_ (
    .clk(CK),
    .d(\DFF_1209.D ),
    .q(\DFF_1209.Q )
  );
  al_dffl _9448_ (
    .clk(CK),
    .d(\DFF_1210.D ),
    .q(\DFF_1210.Q )
  );
  al_dffl _9449_ (
    .clk(CK),
    .d(\DFF_1214.D ),
    .q(\DFF_1214.Q )
  );
  al_dffl _9450_ (
    .clk(CK),
    .d(\DFF_1215.D ),
    .q(\DFF_1215.Q )
  );
  al_dffl _9451_ (
    .clk(CK),
    .d(\DFF_1216.D ),
    .q(\DFF_1216.Q )
  );
  al_dffl _9452_ (
    .clk(CK),
    .d(\DFF_1217.D ),
    .q(\DFF_1217.Q )
  );
  al_dffl _9453_ (
    .clk(CK),
    .d(\DFF_1218.D ),
    .q(\DFF_1218.Q )
  );
  al_dffl _9454_ (
    .clk(CK),
    .d(\DFF_1219.D ),
    .q(\DFF_1219.Q )
  );
  al_dffl _9455_ (
    .clk(CK),
    .d(\DFF_1220.D ),
    .q(\DFF_1220.Q )
  );
  al_dffl _9456_ (
    .clk(CK),
    .d(\DFF_1221.D ),
    .q(\DFF_1221.Q )
  );
  al_dffl _9457_ (
    .clk(CK),
    .d(\DFF_1222.D ),
    .q(\DFF_1222.Q )
  );
  al_dffl _9458_ (
    .clk(CK),
    .d(\DFF_1223.D ),
    .q(\DFF_1223.Q )
  );
  al_dffl _9459_ (
    .clk(CK),
    .d(\DFF_1224.D ),
    .q(\DFF_1224.Q )
  );
  al_dffl _9460_ (
    .clk(CK),
    .d(\DFF_1225.D ),
    .q(\DFF_1225.Q )
  );
  al_dffl _9461_ (
    .clk(CK),
    .d(\DFF_1226.D ),
    .q(\DFF_1226.Q )
  );
  al_dffl _9462_ (
    .clk(CK),
    .d(\DFF_1227.D ),
    .q(\DFF_1227.Q )
  );
  al_dffl _9463_ (
    .clk(CK),
    .d(\DFF_1228.D ),
    .q(\DFF_1228.Q )
  );
  al_dffl _9464_ (
    .clk(CK),
    .d(\DFF_1229.D ),
    .q(\DFF_1229.Q )
  );
  al_dffl _9465_ (
    .clk(CK),
    .d(\DFF_1230.D ),
    .q(\DFF_1230.Q )
  );
  al_dffl _9466_ (
    .clk(CK),
    .d(\DFF_1231.D ),
    .q(\DFF_1231.Q )
  );
  al_dffl _9467_ (
    .clk(CK),
    .d(\DFF_1232.D ),
    .q(\DFF_1232.Q )
  );
  al_dffl _9468_ (
    .clk(CK),
    .d(\DFF_1233.D ),
    .q(\DFF_1233.Q )
  );
  al_dffl _9469_ (
    .clk(CK),
    .d(\DFF_1234.D ),
    .q(\DFF_1234.Q )
  );
  al_dffl _9470_ (
    .clk(CK),
    .d(\DFF_1235.D ),
    .q(\DFF_1235.Q )
  );
  al_dffl _9471_ (
    .clk(CK),
    .d(\DFF_1236.D ),
    .q(\DFF_1236.Q )
  );
  al_dffl _9472_ (
    .clk(CK),
    .d(\DFF_1237.D ),
    .q(\DFF_1237.Q )
  );
  al_dffl _9473_ (
    .clk(CK),
    .d(\DFF_1238.D ),
    .q(\DFF_1238.Q )
  );
  al_dffl _9474_ (
    .clk(CK),
    .d(\DFF_1239.D ),
    .q(\DFF_1239.Q )
  );
  al_dffl _9475_ (
    .clk(CK),
    .d(\DFF_1240.D ),
    .q(\DFF_1240.Q )
  );
  al_dffl _9476_ (
    .clk(CK),
    .d(\DFF_1241.D ),
    .q(\DFF_1241.Q )
  );
  al_dffl _9477_ (
    .clk(CK),
    .d(\DFF_1242.D ),
    .q(\DFF_1242.Q )
  );
  al_dffl _9478_ (
    .clk(CK),
    .d(\DFF_1243.D ),
    .q(\DFF_1243.Q )
  );
  al_dffl _9479_ (
    .clk(CK),
    .d(\DFF_1244.D ),
    .q(\DFF_1244.Q )
  );
  al_dffl _9480_ (
    .clk(CK),
    .d(\DFF_1245.D ),
    .q(\DFF_1245.Q )
  );
  al_dffl _9481_ (
    .clk(CK),
    .d(\DFF_1246.D ),
    .q(\DFF_1246.Q )
  );
  al_dffl _9482_ (
    .clk(CK),
    .d(\DFF_1247.D ),
    .q(\DFF_1247.Q )
  );
  al_dffl _9483_ (
    .clk(CK),
    .d(\DFF_1248.D ),
    .q(\DFF_1248.Q )
  );
  al_dffl _9484_ (
    .clk(CK),
    .d(\DFF_1249.D ),
    .q(\DFF_1249.Q )
  );
  al_dffl _9485_ (
    .clk(CK),
    .d(\DFF_1250.D ),
    .q(\DFF_1250.Q )
  );
  al_dffl _9486_ (
    .clk(CK),
    .d(\DFF_1251.D ),
    .q(\DFF_1251.Q )
  );
  al_dffl _9487_ (
    .clk(CK),
    .d(\DFF_1252.D ),
    .q(\DFF_1252.Q )
  );
  al_dffl _9488_ (
    .clk(CK),
    .d(\DFF_1253.D ),
    .q(\DFF_1253.Q )
  );
  al_dffl _9489_ (
    .clk(CK),
    .d(\DFF_1254.D ),
    .q(\DFF_1254.Q )
  );
  al_dffl _9490_ (
    .clk(CK),
    .d(\DFF_1255.D ),
    .q(\DFF_1255.Q )
  );
  al_dffl _9491_ (
    .clk(CK),
    .d(\DFF_1256.D ),
    .q(\DFF_1256.Q )
  );
  al_dffl _9492_ (
    .clk(CK),
    .d(\DFF_1257.D ),
    .q(\DFF_1257.Q )
  );
  al_dffl _9493_ (
    .clk(CK),
    .d(\DFF_1258.D ),
    .q(\DFF_1258.Q )
  );
  al_dffl _9494_ (
    .clk(CK),
    .d(\DFF_1259.D ),
    .q(\DFF_1259.Q )
  );
  al_dffl _9495_ (
    .clk(CK),
    .d(\DFF_1260.D ),
    .q(\DFF_1260.Q )
  );
  al_dffl _9496_ (
    .clk(CK),
    .d(\DFF_1261.D ),
    .q(\DFF_1261.Q )
  );
  al_dffl _9497_ (
    .clk(CK),
    .d(\DFF_1262.D ),
    .q(\DFF_1262.Q )
  );
  al_dffl _9498_ (
    .clk(CK),
    .d(\DFF_1263.D ),
    .q(\DFF_1263.Q )
  );
  al_dffl _9499_ (
    .clk(CK),
    .d(\DFF_1264.D ),
    .q(\DFF_1264.Q )
  );
  al_dffl _9500_ (
    .clk(CK),
    .d(\DFF_1265.D ),
    .q(\DFF_1265.Q )
  );
  al_dffl _9501_ (
    .clk(CK),
    .d(\DFF_1266.D ),
    .q(\DFF_1266.Q )
  );
  al_dffl _9502_ (
    .clk(CK),
    .d(\DFF_1267.D ),
    .q(\DFF_1267.Q )
  );
  al_dffl _9503_ (
    .clk(CK),
    .d(\DFF_1268.D ),
    .q(\DFF_1268.Q )
  );
  al_dffl _9504_ (
    .clk(CK),
    .d(\DFF_1269.D ),
    .q(\DFF_1269.Q )
  );
  al_dffl _9505_ (
    .clk(CK),
    .d(\DFF_1270.D ),
    .q(\DFF_1270.Q )
  );
  al_dffl _9506_ (
    .clk(CK),
    .d(\DFF_1271.D ),
    .q(\DFF_1271.Q )
  );
  al_dffl _9507_ (
    .clk(CK),
    .d(\DFF_1272.D ),
    .q(\DFF_1272.Q )
  );
  al_dffl _9508_ (
    .clk(CK),
    .d(\DFF_1273.D ),
    .q(\DFF_1273.Q )
  );
  al_dffl _9509_ (
    .clk(CK),
    .d(\DFF_1274.D ),
    .q(\DFF_1274.Q )
  );
  al_dffl _9510_ (
    .clk(CK),
    .d(\DFF_1275.D ),
    .q(\DFF_1275.Q )
  );
  al_dffl _9511_ (
    .clk(CK),
    .d(\DFF_1276.D ),
    .q(\DFF_1276.Q )
  );
  al_dffl _9512_ (
    .clk(CK),
    .d(\DFF_1277.D ),
    .q(\DFF_1277.Q )
  );
  al_dffl _9513_ (
    .clk(CK),
    .d(\DFF_1278.D ),
    .q(\DFF_1278.Q )
  );
  al_dffl _9514_ (
    .clk(CK),
    .d(\DFF_1279.D ),
    .q(\DFF_1279.Q )
  );
  al_dffl _9515_ (
    .clk(CK),
    .d(\DFF_1280.D ),
    .q(\DFF_1280.Q )
  );
  al_dffl _9516_ (
    .clk(CK),
    .d(\DFF_1281.D ),
    .q(\DFF_1281.Q )
  );
  al_dffl _9517_ (
    .clk(CK),
    .d(\DFF_1282.D ),
    .q(\DFF_1282.Q )
  );
  al_dffl _9518_ (
    .clk(CK),
    .d(\DFF_1283.D ),
    .q(\DFF_1283.Q )
  );
  al_dffl _9519_ (
    .clk(CK),
    .d(\DFF_1284.D ),
    .q(\DFF_1284.Q )
  );
  al_dffl _9520_ (
    .clk(CK),
    .d(\DFF_1285.D ),
    .q(\DFF_1285.Q )
  );
  al_dffl _9521_ (
    .clk(CK),
    .d(\DFF_1286.D ),
    .q(\DFF_1286.Q )
  );
  al_dffl _9522_ (
    .clk(CK),
    .d(\DFF_1287.D ),
    .q(\DFF_1287.Q )
  );
  al_dffl _9523_ (
    .clk(CK),
    .d(\DFF_1288.D ),
    .q(\DFF_1288.Q )
  );
  al_dffl _9524_ (
    .clk(CK),
    .d(\DFF_1289.D ),
    .q(\DFF_1289.Q )
  );
  al_dffl _9525_ (
    .clk(CK),
    .d(\DFF_1290.D ),
    .q(\DFF_1290.Q )
  );
  al_dffl _9526_ (
    .clk(CK),
    .d(\DFF_1291.D ),
    .q(\DFF_1291.Q )
  );
  al_dffl _9527_ (
    .clk(CK),
    .d(\DFF_1292.D ),
    .q(\DFF_1292.Q )
  );
  al_dffl _9528_ (
    .clk(CK),
    .d(\DFF_1293.D ),
    .q(\DFF_1293.Q )
  );
  al_dffl _9529_ (
    .clk(CK),
    .d(\DFF_1294.D ),
    .q(\DFF_1294.Q )
  );
  al_dffl _9530_ (
    .clk(CK),
    .d(\DFF_1295.D ),
    .q(\DFF_1295.Q )
  );
  al_dffl _9531_ (
    .clk(CK),
    .d(\DFF_1296.D ),
    .q(\DFF_1296.Q )
  );
  al_dffl _9532_ (
    .clk(CK),
    .d(\DFF_1296.Q ),
    .q(\DFF_1297.Q )
  );
  al_dffl _9533_ (
    .clk(CK),
    .d(\DFF_1297.Q ),
    .q(\DFF_1302.Q )
  );
  al_dffl _9534_ (
    .clk(CK),
    .d(\DFF_1303.D ),
    .q(\DFF_1303.Q )
  );
  al_dffl _9535_ (
    .clk(CK),
    .d(\DFF_1304.D ),
    .q(\DFF_1304.Q )
  );
  al_dffl _9536_ (
    .clk(CK),
    .d(\DFF_1305.D ),
    .q(\DFF_1305.Q )
  );
  al_dffl _9537_ (
    .clk(CK),
    .d(\DFF_1306.D ),
    .q(\DFF_1306.Q )
  );
  al_dffl _9538_ (
    .clk(CK),
    .d(\DFF_1307.D ),
    .q(\DFF_1307.Q )
  );
  al_dffl _9539_ (
    .clk(CK),
    .d(\DFF_1308.D ),
    .q(\DFF_1308.Q )
  );
  al_dffl _9540_ (
    .clk(CK),
    .d(\DFF_1309.D ),
    .q(\DFF_1309.Q )
  );
  al_dffl _9541_ (
    .clk(CK),
    .d(\DFF_1310.D ),
    .q(\DFF_1310.Q )
  );
  al_dffl _9542_ (
    .clk(CK),
    .d(\DFF_1311.D ),
    .q(\DFF_1311.Q )
  );
  al_dffl _9543_ (
    .clk(CK),
    .d(\DFF_1312.D ),
    .q(\DFF_1312.Q )
  );
  al_dffl _9544_ (
    .clk(CK),
    .d(\DFF_1313.D ),
    .q(\DFF_1313.Q )
  );
  al_dffl _9545_ (
    .clk(CK),
    .d(\DFF_1314.D ),
    .q(\DFF_1314.Q )
  );
  al_dffl _9546_ (
    .clk(CK),
    .d(\DFF_1315.D ),
    .q(\DFF_1315.Q )
  );
  al_dffl _9547_ (
    .clk(CK),
    .d(\DFF_1316.D ),
    .q(\DFF_1316.Q )
  );
  al_dffl _9548_ (
    .clk(CK),
    .d(\DFF_1317.D ),
    .q(\DFF_1317.Q )
  );
  al_dffl _9549_ (
    .clk(CK),
    .d(\DFF_1318.D ),
    .q(\DFF_1318.Q )
  );
  al_dffl _9550_ (
    .clk(CK),
    .d(\DFF_1319.D ),
    .q(\DFF_1319.Q )
  );
  al_dffl _9551_ (
    .clk(CK),
    .d(\DFF_1320.D ),
    .q(\DFF_1320.Q )
  );
  al_dffl _9552_ (
    .clk(CK),
    .d(\DFF_1321.D ),
    .q(\DFF_1321.Q )
  );
  al_dffl _9553_ (
    .clk(CK),
    .d(\DFF_1322.D ),
    .q(\DFF_1322.Q )
  );
  al_dffl _9554_ (
    .clk(CK),
    .d(\DFF_1323.D ),
    .q(\DFF_1323.Q )
  );
  al_dffl _9555_ (
    .clk(CK),
    .d(\DFF_1324.D ),
    .q(\DFF_1324.Q )
  );
  al_dffl _9556_ (
    .clk(CK),
    .d(\DFF_1325.D ),
    .q(\DFF_1325.Q )
  );
  al_dffl _9557_ (
    .clk(CK),
    .d(\DFF_1326.D ),
    .q(\DFF_1326.Q )
  );
  al_dffl _9558_ (
    .clk(CK),
    .d(\DFF_1327.D ),
    .q(\DFF_1327.Q )
  );
  al_dffl _9559_ (
    .clk(CK),
    .d(\DFF_1328.D ),
    .q(\DFF_1328.Q )
  );
  al_dffl _9560_ (
    .clk(CK),
    .d(\DFF_1329.D ),
    .q(\DFF_1329.Q )
  );
  al_dffl _9561_ (
    .clk(CK),
    .d(\DFF_1330.D ),
    .q(\DFF_1330.Q )
  );
  al_dffl _9562_ (
    .clk(CK),
    .d(\DFF_1331.D ),
    .q(\DFF_1331.Q )
  );
  al_dffl _9563_ (
    .clk(CK),
    .d(\DFF_1332.D ),
    .q(\DFF_1332.Q )
  );
  al_dffl _9564_ (
    .clk(CK),
    .d(\DFF_1333.D ),
    .q(\DFF_1333.Q )
  );
  al_dffl _9565_ (
    .clk(CK),
    .d(\DFF_1334.D ),
    .q(\DFF_1334.Q )
  );
  al_dffl _9566_ (
    .clk(CK),
    .d(\DFF_1335.D ),
    .q(\DFF_1335.Q )
  );
  al_dffl _9567_ (
    .clk(CK),
    .d(\DFF_1336.D ),
    .q(\DFF_1336.Q )
  );
  al_dffl _9568_ (
    .clk(CK),
    .d(\DFF_1337.D ),
    .q(\DFF_1337.Q )
  );
  al_dffl _9569_ (
    .clk(CK),
    .d(\DFF_1338.D ),
    .q(\DFF_1338.Q )
  );
  al_dffl _9570_ (
    .clk(CK),
    .d(\DFF_1339.D ),
    .q(\DFF_1339.Q )
  );
  al_dffl _9571_ (
    .clk(CK),
    .d(\DFF_1340.D ),
    .q(\DFF_1340.Q )
  );
  al_dffl _9572_ (
    .clk(CK),
    .d(\DFF_1341.D ),
    .q(\DFF_1341.Q )
  );
  al_dffl _9573_ (
    .clk(CK),
    .d(\DFF_1342.D ),
    .q(\DFF_1342.Q )
  );
  al_dffl _9574_ (
    .clk(CK),
    .d(\DFF_1343.D ),
    .q(\DFF_1343.Q )
  );
  al_dffl _9575_ (
    .clk(CK),
    .d(\DFF_1344.D ),
    .q(\DFF_1344.Q )
  );
  al_dffl _9576_ (
    .clk(CK),
    .d(\DFF_1345.D ),
    .q(\DFF_1345.Q )
  );
  al_dffl _9577_ (
    .clk(CK),
    .d(\DFF_1346.D ),
    .q(\DFF_1346.Q )
  );
  al_dffl _9578_ (
    .clk(CK),
    .d(\DFF_1347.D ),
    .q(\DFF_1347.Q )
  );
  al_dffl _9579_ (
    .clk(CK),
    .d(\DFF_1348.D ),
    .q(\DFF_1348.Q )
  );
  al_dffl _9580_ (
    .clk(CK),
    .d(\DFF_1348.Q ),
    .q(\DFF_1349.Q )
  );
  al_dffl _9581_ (
    .clk(CK),
    .d(\DFF_1350.D ),
    .q(\DFF_1350.Q )
  );
  al_dffl _9582_ (
    .clk(CK),
    .d(\DFF_1350.Q ),
    .q(\DFF_1351.Q )
  );
  al_dffl _9583_ (
    .clk(CK),
    .d(\DFF_1352.D ),
    .q(\DFF_1352.Q )
  );
  al_dffl _9584_ (
    .clk(CK),
    .d(\DFF_1352.Q ),
    .q(\DFF_1353.Q )
  );
  al_dffl _9585_ (
    .clk(CK),
    .d(\DFF_1354.D ),
    .q(\DFF_1354.Q )
  );
  al_dffl _9586_ (
    .clk(CK),
    .d(\DFF_1354.Q ),
    .q(\DFF_1355.Q )
  );
  al_dffl _9587_ (
    .clk(CK),
    .d(\DFF_1356.D ),
    .q(\DFF_1356.Q )
  );
  al_dffl _9588_ (
    .clk(CK),
    .d(\DFF_1356.Q ),
    .q(\DFF_1357.Q )
  );
  al_dffl _9589_ (
    .clk(CK),
    .d(\DFF_1358.D ),
    .q(\DFF_1358.Q )
  );
  al_dffl _9590_ (
    .clk(CK),
    .d(\DFF_1358.Q ),
    .q(\DFF_1359.Q )
  );
  al_dffl _9591_ (
    .clk(CK),
    .d(\DFF_1360.D ),
    .q(\DFF_1360.Q )
  );
  al_dffl _9592_ (
    .clk(CK),
    .d(\DFF_1360.Q ),
    .q(\DFF_1361.Q )
  );
  al_dffl _9593_ (
    .clk(CK),
    .d(\DFF_1362.D ),
    .q(\DFF_1362.Q )
  );
  al_dffl _9594_ (
    .clk(CK),
    .d(\DFF_1362.Q ),
    .q(\DFF_1363.Q )
  );
  al_dffl _9595_ (
    .clk(CK),
    .d(\DFF_91.Q ),
    .q(\DFF_1364.Q )
  );
  al_dffl _9596_ (
    .clk(CK),
    .d(\DFF_1364.Q ),
    .q(\DFF_1365.Q )
  );
  al_dffl _9597_ (
    .clk(CK),
    .d(\DFF_1366.D ),
    .q(\DFF_1366.Q )
  );
  al_dffl _9598_ (
    .clk(CK),
    .d(\DFF_1367.D ),
    .q(\DFF_1367.Q )
  );
  al_dffl _9599_ (
    .clk(CK),
    .d(\DFF_1378.D ),
    .q(\DFF_1378.Q )
  );
  al_dffl _9600_ (
    .clk(CK),
    .d(\DFF_1303.Q ),
    .q(\DFF_1379.Q )
  );
  al_dffl _9601_ (
    .clk(CK),
    .d(\DFF_1379.Q ),
    .q(\DFF_1380.Q )
  );
  al_dffl _9602_ (
    .clk(CK),
    .d(\DFF_1304.Q ),
    .q(\DFF_1381.Q )
  );
  al_dffl _9603_ (
    .clk(CK),
    .d(\DFF_1381.Q ),
    .q(\DFF_1382.Q )
  );
  al_dffl _9604_ (
    .clk(CK),
    .d(\DFF_1305.Q ),
    .q(\DFF_1383.Q )
  );
  al_dffl _9605_ (
    .clk(CK),
    .d(\DFF_1383.Q ),
    .q(\DFF_1384.Q )
  );
  al_dffl _9606_ (
    .clk(CK),
    .d(\DFF_1306.Q ),
    .q(\DFF_1385.Q )
  );
  al_dffl _9607_ (
    .clk(CK),
    .d(\DFF_1385.Q ),
    .q(\DFF_1386.Q )
  );
  al_dffl _9608_ (
    .clk(CK),
    .d(\DFF_1307.Q ),
    .q(\DFF_1387.Q )
  );
  al_dffl _9609_ (
    .clk(CK),
    .d(\DFF_1387.Q ),
    .q(\DFF_1388.Q )
  );
  al_dffl _9610_ (
    .clk(CK),
    .d(\DFF_1308.Q ),
    .q(\DFF_1389.Q )
  );
  al_dffl _9611_ (
    .clk(CK),
    .d(\DFF_1389.Q ),
    .q(\DFF_1390.Q )
  );
  al_dffl _9612_ (
    .clk(CK),
    .d(\DFF_1309.Q ),
    .q(\DFF_1391.Q )
  );
  al_dffl _9613_ (
    .clk(CK),
    .d(\DFF_1391.Q ),
    .q(\DFF_1392.Q )
  );
  al_dffl _9614_ (
    .clk(CK),
    .d(\DFF_1310.Q ),
    .q(\DFF_1393.Q )
  );
  al_dffl _9615_ (
    .clk(CK),
    .d(\DFF_1393.Q ),
    .q(\DFF_1394.Q )
  );
  al_dffl _9616_ (
    .clk(CK),
    .d(\DFF_1311.Q ),
    .q(\DFF_1395.Q )
  );
  al_dffl _9617_ (
    .clk(CK),
    .d(\DFF_1395.Q ),
    .q(\DFF_1396.Q )
  );
  al_dffl _9618_ (
    .clk(CK),
    .d(\DFF_1312.Q ),
    .q(\DFF_1397.Q )
  );
  al_dffl _9619_ (
    .clk(CK),
    .d(\DFF_1397.Q ),
    .q(\DFF_1398.Q )
  );
  al_dffl _9620_ (
    .clk(CK),
    .d(\DFF_1313.Q ),
    .q(\DFF_1399.Q )
  );
  al_dffl _9621_ (
    .clk(CK),
    .d(\DFF_1399.Q ),
    .q(\DFF_1400.Q )
  );
  al_dffl _9622_ (
    .clk(CK),
    .d(\DFF_1314.Q ),
    .q(\DFF_1401.Q )
  );
  al_dffl _9623_ (
    .clk(CK),
    .d(\DFF_1401.Q ),
    .q(\DFF_1402.Q )
  );
  al_dffl _9624_ (
    .clk(CK),
    .d(\DFF_1409.D ),
    .q(\DFF_1409.Q )
  );
  al_dffl _9625_ (
    .clk(CK),
    .d(\DFF_1410.D ),
    .q(\DFF_1410.Q )
  );
  al_dffl _9626_ (
    .clk(CK),
    .d(\DFF_1411.D ),
    .q(\DFF_1411.Q )
  );
  al_dffl _9627_ (
    .clk(CK),
    .d(\DFF_1412.D ),
    .q(\DFF_1412.Q )
  );
  al_dffl _9628_ (
    .clk(CK),
    .d(\DFF_1412.Q ),
    .q(\DFF_1413.Q )
  );
  al_dffl _9629_ (
    .clk(CK),
    .d(\DFF_1413.Q ),
    .q(\DFF_1414.Q )
  );
  al_dffl _9630_ (
    .clk(CK),
    .d(\DFF_1433.Q ),
    .q(\DFF_1415.Q )
  );
  al_dffl _9631_ (
    .clk(CK),
    .d(\DFF_1415.Q ),
    .q(\DFF_1416.Q )
  );
  al_dffl _9632_ (
    .clk(CK),
    .d(\DFF_1434.Q ),
    .q(\DFF_1417.Q )
  );
  al_dffl _9633_ (
    .clk(CK),
    .d(\DFF_1417.Q ),
    .q(\DFF_1418.Q )
  );
  al_dffl _9634_ (
    .clk(CK),
    .d(\DFF_1435.Q ),
    .q(\DFF_1419.Q )
  );
  al_dffl _9635_ (
    .clk(CK),
    .d(\DFF_1419.Q ),
    .q(\DFF_1420.Q )
  );
  al_dffl _9636_ (
    .clk(CK),
    .d(\DFF_1442.Q ),
    .q(\DFF_1421.Q )
  );
  al_dffl _9637_ (
    .clk(CK),
    .d(\DFF_1421.Q ),
    .q(\DFF_1422.Q )
  );
  al_dffl _9638_ (
    .clk(CK),
    .d(\DFF_1443.Q ),
    .q(\DFF_1423.Q )
  );
  al_dffl _9639_ (
    .clk(CK),
    .d(\DFF_1423.Q ),
    .q(\DFF_1424.Q )
  );
  al_dffl _9640_ (
    .clk(CK),
    .d(\DFF_1444.Q ),
    .q(\DFF_1425.Q )
  );
  al_dffl _9641_ (
    .clk(CK),
    .d(\DFF_1425.Q ),
    .q(\DFF_1426.Q )
  );
  al_dffl _9642_ (
    .clk(CK),
    .d(\DFF_3.Q ),
    .q(\DFF_1427.Q )
  );
  al_dffl _9643_ (
    .clk(CK),
    .d(\DFF_1427.Q ),
    .q(\DFF_1428.Q )
  );
  al_dffl _9644_ (
    .clk(CK),
    .d(\DFF_1428.Q ),
    .q(\DFF_1429.Q )
  );
  al_dffl _9645_ (
    .clk(CK),
    .d(\DFF_1430.D ),
    .q(\DFF_1430.Q )
  );
  al_dffl _9646_ (
    .clk(CK),
    .d(\DFF_1431.D ),
    .q(\DFF_1431.Q )
  );
  al_dffl _9647_ (
    .clk(CK),
    .d(\DFF_1432.D ),
    .q(\DFF_1432.Q )
  );
  al_dffl _9648_ (
    .clk(CK),
    .d(\DFF_1433.D ),
    .q(\DFF_1433.Q )
  );
  al_dffl _9649_ (
    .clk(CK),
    .d(\DFF_1434.D ),
    .q(\DFF_1434.Q )
  );
  al_dffl _9650_ (
    .clk(CK),
    .d(\DFF_1435.D ),
    .q(\DFF_1435.Q )
  );
  al_dffl _9651_ (
    .clk(CK),
    .d(\DFF_1436.D ),
    .q(\DFF_1436.Q )
  );
  al_dffl _9652_ (
    .clk(CK),
    .d(\DFF_1437.D ),
    .q(\DFF_1437.Q )
  );
  al_dffl _9653_ (
    .clk(CK),
    .d(\DFF_1438.D ),
    .q(\DFF_1438.Q )
  );
  al_dffl _9654_ (
    .clk(CK),
    .d(\DFF_1439.D ),
    .q(\DFF_1439.Q )
  );
  al_dffl _9655_ (
    .clk(CK),
    .d(\DFF_1440.D ),
    .q(\DFF_1440.Q )
  );
  al_dffl _9656_ (
    .clk(CK),
    .d(\DFF_1441.D ),
    .q(\DFF_1441.Q )
  );
  al_dffl _9657_ (
    .clk(CK),
    .d(\DFF_1442.D ),
    .q(\DFF_1442.Q )
  );
  al_dffl _9658_ (
    .clk(CK),
    .d(\DFF_1443.D ),
    .q(\DFF_1443.Q )
  );
  al_dffl _9659_ (
    .clk(CK),
    .d(\DFF_1444.D ),
    .q(\DFF_1444.Q )
  );
  al_dffl _9660_ (
    .clk(CK),
    .d(\DFF_1445.D ),
    .q(\DFF_1445.Q )
  );
  al_dffl _9661_ (
    .clk(CK),
    .d(\DFF_1445.Q ),
    .q(\DFF_1446.Q )
  );
  al_dffl _9662_ (
    .clk(CK),
    .d(\DFF_1446.Q ),
    .q(\DFF_1447.Q )
  );
  al_dffl _9663_ (
    .clk(CK),
    .d(\DFF_1448.D ),
    .q(\DFF_1448.Q )
  );
  al_dffl _9664_ (
    .clk(CK),
    .d(\DFF_1448.Q ),
    .q(\DFF_1449.Q )
  );
  al_dffl _9665_ (
    .clk(CK),
    .d(\DFF_1450.D ),
    .q(\DFF_1450.Q )
  );
  al_dffl _9666_ (
    .clk(CK),
    .d(\DFF_1451.D ),
    .q(\DFF_1451.Q )
  );
  al_dffl _9667_ (
    .clk(CK),
    .d(\DFF_1451.Q ),
    .q(\DFF_1452.Q )
  );
  al_dffl _9668_ (
    .clk(CK),
    .d(\DFF_1453.D ),
    .q(\DFF_1453.Q )
  );
  al_dffl _9669_ (
    .clk(CK),
    .d(\DFF_1453.Q ),
    .q(\DFF_1454.Q )
  );
  al_dffl _9670_ (
    .clk(CK),
    .d(\DFF_1455.D ),
    .q(\DFF_1455.Q )
  );
  al_dffl _9671_ (
    .clk(CK),
    .d(\DFF_1456.D ),
    .q(\DFF_1456.Q )
  );
  al_dffl _9672_ (
    .clk(CK),
    .d(\DFF_1457.D ),
    .q(\DFF_1457.Q )
  );
  al_dffl _9673_ (
    .clk(CK),
    .d(\DFF_1458.D ),
    .q(\DFF_1458.Q )
  );
  al_dffl _9674_ (
    .clk(CK),
    .d(\DFF_1459.D ),
    .q(\DFF_1459.Q )
  );
  al_dffl _9675_ (
    .clk(CK),
    .d(\DFF_1460.D ),
    .q(\DFF_1460.Q )
  );
  al_dffl _9676_ (
    .clk(CK),
    .d(\DFF_1461.D ),
    .q(\DFF_1461.Q )
  );
  al_dffl _9677_ (
    .clk(CK),
    .d(\DFF_1462.D ),
    .q(\DFF_1462.Q )
  );
  al_dffl _9678_ (
    .clk(CK),
    .d(\DFF_1463.D ),
    .q(\DFF_1463.Q )
  );
  al_dffl _9679_ (
    .clk(CK),
    .d(\DFF_1464.D ),
    .q(\DFF_1464.Q )
  );
  al_dffl _9680_ (
    .clk(CK),
    .d(\DFF_1465.D ),
    .q(\DFF_1465.Q )
  );
  al_dffl _9681_ (
    .clk(CK),
    .d(\DFF_1466.D ),
    .q(\DFF_1466.Q )
  );
  al_dffl _9682_ (
    .clk(CK),
    .d(\DFF_1467.D ),
    .q(\DFF_1467.Q )
  );
  al_dffl _9683_ (
    .clk(CK),
    .d(\DFF_1468.D ),
    .q(\DFF_1468.Q )
  );
  al_dffl _9684_ (
    .clk(CK),
    .d(\DFF_1469.D ),
    .q(\DFF_1469.Q )
  );
  al_dffl _9685_ (
    .clk(CK),
    .d(\DFF_1470.D ),
    .q(\DFF_1470.Q )
  );
  al_dffl _9686_ (
    .clk(CK),
    .d(\DFF_1471.D ),
    .q(\DFF_1471.Q )
  );
  al_dffl _9687_ (
    .clk(CK),
    .d(\DFF_1472.D ),
    .q(\DFF_1472.Q )
  );
  al_dffl _9688_ (
    .clk(CK),
    .d(\DFF_1473.D ),
    .q(\DFF_1473.Q )
  );
  al_dffl _9689_ (
    .clk(CK),
    .d(\DFF_1474.D ),
    .q(\DFF_1474.Q )
  );
  al_dffl _9690_ (
    .clk(CK),
    .d(\DFF_1475.D ),
    .q(\DFF_1475.Q )
  );
  al_dffl _9691_ (
    .clk(CK),
    .d(\DFF_1476.D ),
    .q(\DFF_1476.Q )
  );
  al_dffl _9692_ (
    .clk(CK),
    .d(\DFF_1477.D ),
    .q(\DFF_1477.Q )
  );
  al_dffl _9693_ (
    .clk(CK),
    .d(\DFF_1478.D ),
    .q(\DFF_1478.Q )
  );
  al_dffl _9694_ (
    .clk(CK),
    .d(\DFF_1479.D ),
    .q(\DFF_1479.Q )
  );
  al_dffl _9695_ (
    .clk(CK),
    .d(\DFF_1480.D ),
    .q(\DFF_1480.Q )
  );
  al_dffl _9696_ (
    .clk(CK),
    .d(\DFF_1481.D ),
    .q(\DFF_1481.Q )
  );
  al_dffl _9697_ (
    .clk(CK),
    .d(\DFF_1452.Q ),
    .q(\DFF_1482.Q )
  );
  al_dffl _9698_ (
    .clk(CK),
    .d(\DFF_1483.D ),
    .q(\DFF_1483.Q )
  );
  al_dffl _9699_ (
    .clk(CK),
    .d(\DFF_1492.D ),
    .q(\DFF_1492.Q )
  );
  al_dffl _9700_ (
    .clk(CK),
    .d(\DFF_1492.Q ),
    .q(\DFF_1493.Q )
  );
  al_dffl _9701_ (
    .clk(CK),
    .d(\DFF_1494.D ),
    .q(\DFF_1494.Q )
  );
  al_dffl _9702_ (
    .clk(CK),
    .d(\DFF_1495.D ),
    .q(\DFF_1495.Q )
  );
  al_dffl _9703_ (
    .clk(CK),
    .d(\DFF_1496.D ),
    .q(\DFF_1496.Q )
  );
  al_dffl _9704_ (
    .clk(CK),
    .d(\DFF_1497.D ),
    .q(\DFF_1497.Q )
  );
  al_dffl _9705_ (
    .clk(CK),
    .d(\DFF_1498.D ),
    .q(\DFF_1498.Q )
  );
  al_dffl _9706_ (
    .clk(CK),
    .d(\DFF_1499.D ),
    .q(\DFF_1499.Q )
  );
  al_dffl _9707_ (
    .clk(CK),
    .d(\DFF_1500.D ),
    .q(\DFF_1500.Q )
  );
  al_dffl _9708_ (
    .clk(CK),
    .d(\DFF_1501.D ),
    .q(\DFF_1501.Q )
  );
  al_dffl _9709_ (
    .clk(CK),
    .d(\DFF_1502.D ),
    .q(\DFF_1502.Q )
  );
  al_dffl _9710_ (
    .clk(CK),
    .d(\DFF_1503.D ),
    .q(\DFF_1503.Q )
  );
  al_dffl _9711_ (
    .clk(CK),
    .d(\DFF_1563.Q ),
    .q(\DFF_1504.Q )
  );
  al_dffl _9712_ (
    .clk(CK),
    .d(\DFF_1504.Q ),
    .q(\DFF_1505.Q )
  );
  al_dffl _9713_ (
    .clk(CK),
    .d(\DFF_1505.Q ),
    .q(\DFF_1506.Q )
  );
  al_dffl _9714_ (
    .clk(CK),
    .d(\DFF_1507.D ),
    .q(\DFF_1507.Q )
  );
  al_dffl _9715_ (
    .clk(CK),
    .d(\DFF_1508.D ),
    .q(\DFF_1508.Q )
  );
  al_dffl _9716_ (
    .clk(CK),
    .d(\DFF_1509.D ),
    .q(\DFF_1509.Q )
  );
  al_dffl _9717_ (
    .clk(CK),
    .d(\DFF_1510.D ),
    .q(\DFF_1510.Q )
  );
  al_dffl _9718_ (
    .clk(CK),
    .d(\DFF_1511.D ),
    .q(\DFF_1511.Q )
  );
  al_dffl _9719_ (
    .clk(CK),
    .d(\DFF_1512.D ),
    .q(\DFF_1512.Q )
  );
  al_dffl _9720_ (
    .clk(CK),
    .d(\DFF_1513.D ),
    .q(\DFF_1513.Q )
  );
  al_dffl _9721_ (
    .clk(CK),
    .d(\DFF_1514.D ),
    .q(\DFF_1514.Q )
  );
  al_dffl _9722_ (
    .clk(CK),
    .d(\DFF_1515.D ),
    .q(\DFF_1515.Q )
  );
  al_dffl _9723_ (
    .clk(CK),
    .d(\DFF_1516.D ),
    .q(\DFF_1516.Q )
  );
  al_dffl _9724_ (
    .clk(CK),
    .d(\DFF_1517.D ),
    .q(\DFF_1517.Q )
  );
  al_dffl _9725_ (
    .clk(CK),
    .d(\DFF_1518.D ),
    .q(\DFF_1518.Q )
  );
  al_dffl _9726_ (
    .clk(CK),
    .d(\DFF_1519.D ),
    .q(\DFF_1519.Q )
  );
  al_dffl _9727_ (
    .clk(CK),
    .d(\DFF_1520.D ),
    .q(\DFF_1520.Q )
  );
  al_dffl _9728_ (
    .clk(CK),
    .d(\DFF_1521.D ),
    .q(\DFF_1521.Q )
  );
  al_dffl _9729_ (
    .clk(CK),
    .d(\DFF_1522.D ),
    .q(\DFF_1522.Q )
  );
  al_dffl _9730_ (
    .clk(CK),
    .d(\DFF_1523.D ),
    .q(\DFF_1523.Q )
  );
  al_dffl _9731_ (
    .clk(CK),
    .d(\DFF_1524.D ),
    .q(\DFF_1524.Q )
  );
  al_dffl _9732_ (
    .clk(CK),
    .d(\DFF_1525.D ),
    .q(\DFF_1525.Q )
  );
  al_dffl _9733_ (
    .clk(CK),
    .d(\DFF_1526.D ),
    .q(\DFF_1526.Q )
  );
  al_dffl _9734_ (
    .clk(CK),
    .d(\DFF_1527.D ),
    .q(\DFF_1527.Q )
  );
  al_dffl _9735_ (
    .clk(CK),
    .d(\DFF_1528.D ),
    .q(\DFF_1528.Q )
  );
  al_dffl _9736_ (
    .clk(CK),
    .d(\DFF_1529.D ),
    .q(\DFF_1529.Q )
  );
  al_dffl _9737_ (
    .clk(CK),
    .d(\DFF_1530.D ),
    .q(\DFF_1530.Q )
  );
  al_dffl _9738_ (
    .clk(CK),
    .d(\DFF_1531.D ),
    .q(\DFF_1531.Q )
  );
  al_dffl _9739_ (
    .clk(CK),
    .d(\DFF_1532.D ),
    .q(\DFF_1532.Q )
  );
  al_dffl _9740_ (
    .clk(CK),
    .d(\DFF_1533.D ),
    .q(\DFF_1533.Q )
  );
  al_dffl _9741_ (
    .clk(CK),
    .d(\DFF_1534.D ),
    .q(\DFF_1534.Q )
  );
  al_dffl _9742_ (
    .clk(CK),
    .d(\DFF_1535.D ),
    .q(\DFF_1535.Q )
  );
  al_dffl _9743_ (
    .clk(CK),
    .d(\DFF_1536.D ),
    .q(\DFF_1536.Q )
  );
  al_dffl _9744_ (
    .clk(CK),
    .d(\DFF_1537.D ),
    .q(\DFF_1537.Q )
  );
  al_dffl _9745_ (
    .clk(CK),
    .d(\DFF_1538.D ),
    .q(\DFF_1538.Q )
  );
  al_dffl _9746_ (
    .clk(CK),
    .d(\DFF_1539.D ),
    .q(\DFF_1539.Q )
  );
  al_dffl _9747_ (
    .clk(CK),
    .d(\DFF_1540.D ),
    .q(\DFF_1540.Q )
  );
  al_dffl _9748_ (
    .clk(CK),
    .d(\DFF_1541.D ),
    .q(\DFF_1541.Q )
  );
  al_dffl _9749_ (
    .clk(CK),
    .d(\DFF_1542.D ),
    .q(\DFF_1542.Q )
  );
  al_dffl _9750_ (
    .clk(CK),
    .d(\DFF_1543.D ),
    .q(\DFF_1543.Q )
  );
  al_dffl _9751_ (
    .clk(CK),
    .d(\DFF_1544.D ),
    .q(\DFF_1544.Q )
  );
  al_dffl _9752_ (
    .clk(CK),
    .d(\DFF_1545.D ),
    .q(\DFF_1545.Q )
  );
  al_dffl _9753_ (
    .clk(CK),
    .d(\DFF_1546.D ),
    .q(\DFF_1546.Q )
  );
  al_dffl _9754_ (
    .clk(CK),
    .d(\DFF_1547.D ),
    .q(\DFF_1547.Q )
  );
  al_dffl _9755_ (
    .clk(CK),
    .d(\DFF_1548.D ),
    .q(\DFF_1548.Q )
  );
  al_dffl _9756_ (
    .clk(CK),
    .d(\DFF_1549.D ),
    .q(\DFF_1549.Q )
  );
  al_dffl _9757_ (
    .clk(CK),
    .d(\DFF_1550.D ),
    .q(\DFF_1550.Q )
  );
  al_dffl _9758_ (
    .clk(CK),
    .d(\DFF_1551.D ),
    .q(\DFF_1551.Q )
  );
  al_dffl _9759_ (
    .clk(CK),
    .d(\DFF_1552.D ),
    .q(\DFF_1552.Q )
  );
  al_dffl _9760_ (
    .clk(CK),
    .d(\DFF_1553.D ),
    .q(\DFF_1553.Q )
  );
  al_dffl _9761_ (
    .clk(CK),
    .d(\DFF_1554.D ),
    .q(\DFF_1554.Q )
  );
  al_dffl _9762_ (
    .clk(CK),
    .d(\DFF_1555.D ),
    .q(\DFF_1555.Q )
  );
  al_dffl _9763_ (
    .clk(CK),
    .d(\DFF_1556.D ),
    .q(\DFF_1556.Q )
  );
  al_dffl _9764_ (
    .clk(CK),
    .d(\DFF_1557.D ),
    .q(\DFF_1557.Q )
  );
  al_dffl _9765_ (
    .clk(CK),
    .d(\DFF_1558.D ),
    .q(\DFF_1558.Q )
  );
  al_dffl _9766_ (
    .clk(CK),
    .d(\DFF_1559.D ),
    .q(\DFF_1559.Q )
  );
  al_dffl _9767_ (
    .clk(CK),
    .d(\DFF_1560.D ),
    .q(\DFF_1560.Q )
  );
  al_dffl _9768_ (
    .clk(CK),
    .d(\DFF_1561.D ),
    .q(\DFF_1561.Q )
  );
  al_dffl _9769_ (
    .clk(CK),
    .d(\DFF_1562.D ),
    .q(\DFF_1562.Q )
  );
  al_dffl _9770_ (
    .clk(CK),
    .d(\DFF_1563.D ),
    .q(\DFF_1563.Q )
  );
  al_dffl _9771_ (
    .clk(CK),
    .d(\DFF_1564.D ),
    .q(\DFF_1564.Q )
  );
  al_dffl _9772_ (
    .clk(CK),
    .d(\DFF_1565.D ),
    .q(\DFF_1565.Q )
  );
  al_dffl _9773_ (
    .clk(CK),
    .d(\DFF_1566.D ),
    .q(\DFF_1566.Q )
  );
  al_dffl _9774_ (
    .clk(CK),
    .d(\DFF_1567.D ),
    .q(\DFF_1567.Q )
  );
  al_dffl _9775_ (
    .clk(CK),
    .d(\DFF_1568.D ),
    .q(\DFF_1568.Q )
  );
  al_dffl _9776_ (
    .clk(CK),
    .d(\DFF_1569.D ),
    .q(\DFF_1569.Q )
  );
  al_dffl _9777_ (
    .clk(CK),
    .d(\DFF_1570.D ),
    .q(\DFF_1570.Q )
  );
  al_dffl _9778_ (
    .clk(CK),
    .d(\DFF_1571.D ),
    .q(\DFF_1571.Q )
  );
  al_dffl _9779_ (
    .clk(CK),
    .d(\DFF_1572.D ),
    .q(\DFF_1572.Q )
  );
  al_dffl _9780_ (
    .clk(CK),
    .d(\DFF_1573.D ),
    .q(\DFF_1573.Q )
  );
  al_dffl _9781_ (
    .clk(CK),
    .d(\DFF_1574.D ),
    .q(\DFF_1574.Q )
  );
  al_dffl _9782_ (
    .clk(CK),
    .d(\DFF_1575.D ),
    .q(\DFF_1575.Q )
  );
  al_dffl _9783_ (
    .clk(CK),
    .d(\DFF_1576.D ),
    .q(\DFF_1576.Q )
  );
  al_dffl _9784_ (
    .clk(CK),
    .d(\DFF_1577.D ),
    .q(\DFF_1577.Q )
  );
  al_dffl _9785_ (
    .clk(CK),
    .d(\DFF_1578.D ),
    .q(\DFF_1578.Q )
  );
  al_dffl _9786_ (
    .clk(CK),
    .d(\DFF_1579.D ),
    .q(\DFF_1579.Q )
  );
  al_dffl _9787_ (
    .clk(CK),
    .d(\DFF_1580.D ),
    .q(\DFF_1580.Q )
  );
  al_dffl _9788_ (
    .clk(CK),
    .d(\DFF_1581.D ),
    .q(\DFF_1581.Q )
  );
  al_dffl _9789_ (
    .clk(CK),
    .d(\DFF_1582.D ),
    .q(\DFF_1582.Q )
  );
  al_dffl _9790_ (
    .clk(CK),
    .d(\DFF_1583.D ),
    .q(\DFF_1583.Q )
  );
  al_dffl _9791_ (
    .clk(CK),
    .d(\DFF_1584.D ),
    .q(\DFF_1584.Q )
  );
  al_dffl _9792_ (
    .clk(CK),
    .d(\DFF_1585.D ),
    .q(\DFF_1585.Q )
  );
  al_dffl _9793_ (
    .clk(CK),
    .d(\DFF_1586.D ),
    .q(\DFF_1586.Q )
  );
  al_dffl _9794_ (
    .clk(CK),
    .d(\DFF_1587.D ),
    .q(\DFF_1587.Q )
  );
  al_dffl _9795_ (
    .clk(CK),
    .d(\DFF_1588.D ),
    .q(\DFF_1588.Q )
  );
  al_dffl _9796_ (
    .clk(CK),
    .d(\DFF_1589.D ),
    .q(\DFF_1589.Q )
  );
  al_dffl _9797_ (
    .clk(CK),
    .d(\DFF_1590.D ),
    .q(\DFF_1590.Q )
  );
  al_dffl _9798_ (
    .clk(CK),
    .d(\DFF_1591.D ),
    .q(\DFF_1591.Q )
  );
  al_dffl _9799_ (
    .clk(CK),
    .d(\DFF_1592.D ),
    .q(\DFF_1592.Q )
  );
  al_dffl _9800_ (
    .clk(CK),
    .d(\DFF_1593.D ),
    .q(\DFF_1593.Q )
  );
  al_dffl _9801_ (
    .clk(CK),
    .d(\DFF_1594.D ),
    .q(\DFF_1594.Q )
  );
  al_dffl _9802_ (
    .clk(CK),
    .d(\DFF_1595.D ),
    .q(\DFF_1595.Q )
  );
  al_dffl _9803_ (
    .clk(CK),
    .d(\DFF_1596.D ),
    .q(\DFF_1596.Q )
  );
  al_dffl _9804_ (
    .clk(CK),
    .d(\DFF_1597.D ),
    .q(\DFF_1597.Q )
  );
  al_dffl _9805_ (
    .clk(CK),
    .d(\DFF_1598.D ),
    .q(\DFF_1598.Q )
  );
  al_dffl _9806_ (
    .clk(CK),
    .d(\DFF_1599.D ),
    .q(\DFF_1599.Q )
  );
  al_dffl _9807_ (
    .clk(CK),
    .d(\DFF_1600.D ),
    .q(\DFF_1600.Q )
  );
  al_dffl _9808_ (
    .clk(CK),
    .d(\DFF_1601.D ),
    .q(\DFF_1601.Q )
  );
  al_dffl _9809_ (
    .clk(CK),
    .d(\DFF_1602.D ),
    .q(\DFF_1602.Q )
  );
  al_dffl _9810_ (
    .clk(CK),
    .d(\DFF_1603.D ),
    .q(\DFF_1603.Q )
  );
  al_dffl _9811_ (
    .clk(CK),
    .d(\DFF_1604.D ),
    .q(\DFF_1604.Q )
  );
  al_dffl _9812_ (
    .clk(CK),
    .d(\DFF_1605.D ),
    .q(\DFF_1605.Q )
  );
  al_dffl _9813_ (
    .clk(CK),
    .d(\DFF_1606.D ),
    .q(\DFF_1606.Q )
  );
  al_dffl _9814_ (
    .clk(CK),
    .d(\DFF_1607.D ),
    .q(\DFF_1607.Q )
  );
  al_dffl _9815_ (
    .clk(CK),
    .d(\DFF_1608.D ),
    .q(\DFF_1608.Q )
  );
  al_dffl _9816_ (
    .clk(CK),
    .d(\DFF_1609.D ),
    .q(\DFF_1609.Q )
  );
  al_dffl _9817_ (
    .clk(CK),
    .d(\DFF_1610.D ),
    .q(\DFF_1610.Q )
  );
  al_dffl _9818_ (
    .clk(CK),
    .d(g3234),
    .q(\DFF_1611.Q )
  );
  al_dffl _9819_ (
    .clk(CK),
    .d(\DFF_1611.Q ),
    .q(\DFF_1612.Q )
  );
  al_dffl _9820_ (
    .clk(CK),
    .d(\DFF_1613.D ),
    .q(\DFF_1613.Q )
  );
  al_dffl _9821_ (
    .clk(CK),
    .d(\DFF_1614.D ),
    .q(\DFF_1614.Q )
  );
  al_dffl _9822_ (
    .clk(CK),
    .d(\DFF_1615.D ),
    .q(\DFF_1615.Q )
  );
  al_dffl _9823_ (
    .clk(CK),
    .d(\DFF_1616.D ),
    .q(\DFF_1616.Q )
  );
  al_dffl _9824_ (
    .clk(CK),
    .d(\DFF_1617.D ),
    .q(\DFF_1617.Q )
  );
  al_dffl _9825_ (
    .clk(CK),
    .d(\DFF_1618.D ),
    .q(\DFF_1618.Q )
  );
  al_dffl _9826_ (
    .clk(CK),
    .d(\DFF_1619.D ),
    .q(\DFF_1619.Q )
  );
  al_dffl _9827_ (
    .clk(CK),
    .d(\DFF_1620.D ),
    .q(\DFF_1620.Q )
  );
  al_dffl _9828_ (
    .clk(CK),
    .d(\DFF_1621.D ),
    .q(\DFF_1621.Q )
  );
  al_dffl _9829_ (
    .clk(CK),
    .d(\DFF_1622.D ),
    .q(\DFF_1622.Q )
  );
  al_dffl _9830_ (
    .clk(CK),
    .d(\DFF_1623.D ),
    .q(\DFF_1623.Q )
  );
  al_dffl _9831_ (
    .clk(CK),
    .d(\DFF_1624.D ),
    .q(\DFF_1624.Q )
  );
  al_dffl _9832_ (
    .clk(CK),
    .d(\DFF_1625.D ),
    .q(\DFF_1625.Q )
  );
  al_dffl _9833_ (
    .clk(CK),
    .d(\DFF_1626.D ),
    .q(\DFF_1626.Q )
  );
  al_dffl _9834_ (
    .clk(CK),
    .d(\DFF_1627.D ),
    .q(\DFF_1627.Q )
  );
  al_dffl _9835_ (
    .clk(CK),
    .d(\DFF_1628.D ),
    .q(\DFF_1628.Q )
  );
  al_dffl _9836_ (
    .clk(CK),
    .d(\DFF_1629.D ),
    .q(\DFF_1629.Q )
  );
  al_dffl _9837_ (
    .clk(CK),
    .d(\DFF_1630.D ),
    .q(\DFF_1630.Q )
  );
  al_dffl _9838_ (
    .clk(CK),
    .d(\DFF_1631.D ),
    .q(\DFF_1631.Q )
  );
  al_dffl _9839_ (
    .clk(CK),
    .d(\DFF_1632.D ),
    .q(\DFF_1632.Q )
  );
  al_dffl _9840_ (
    .clk(CK),
    .d(\DFF_1633.D ),
    .q(\DFF_1633.Q )
  );
  al_dffl _9841_ (
    .clk(CK),
    .d(\DFF_1634.D ),
    .q(\DFF_1634.Q )
  );
  al_dffl _9842_ (
    .clk(CK),
    .d(\DFF_1635.D ),
    .q(\DFF_1635.Q )
  );
  assign \DFF_0.CK  = CK;
  assign \DFF_0.D  = g51;
  assign \DFF_0.Q  = \DFF_17.Q ;
  assign \DFF_1.CK  = CK;
  assign \DFF_10.CK  = CK;
  assign \DFF_100.CK  = CK;
  assign \DFF_1000.CK  = CK;
  assign \DFF_1001.CK  = CK;
  assign \DFF_1001.D  = \DFF_1000.Q ;
  assign \DFF_1002.CK  = CK;
  assign \DFF_1003.CK  = CK;
  assign \DFF_1003.D  = \DFF_1002.Q ;
  assign \DFF_1004.CK  = CK;
  assign \DFF_1005.CK  = CK;
  assign \DFF_1005.D  = \DFF_1004.Q ;
  assign \DFF_1006.CK  = CK;
  assign \DFF_1007.CK  = CK;
  assign \DFF_1007.D  = \DFF_1006.Q ;
  assign \DFF_1008.CK  = CK;
  assign \DFF_1009.CK  = CK;
  assign \DFF_1009.D  = \DFF_1008.Q ;
  assign \DFF_101.CK  = CK;
  assign \DFF_1010.CK  = CK;
  assign \DFF_1011.CK  = CK;
  assign \DFF_1011.D  = \DFF_1010.Q ;
  assign \DFF_1012.CK  = CK;
  assign \DFF_1013.CK  = CK;
  assign \DFF_1013.D  = \DFF_1012.Q ;
  assign \DFF_1014.CK  = CK;
  assign \DFF_1014.D  = \DFF_46.Q ;
  assign \DFF_1015.CK  = CK;
  assign \DFF_1015.D  = \DFF_1014.Q ;
  assign \DFF_1016.CK  = CK;
  assign \DFF_1017.CK  = CK;
  assign \DFF_1018.CK  = CK;
  assign \DFF_1019.CK  = CK;
  assign \DFF_102.CK  = CK;
  assign \DFF_1020.CK  = CK;
  assign \DFF_1021.CK  = CK;
  assign \DFF_1022.CK  = CK;
  assign \DFF_1023.CK  = CK;
  assign \DFF_1024.CK  = CK;
  assign \DFF_1025.CK  = CK;
  assign \DFF_1026.CK  = CK;
  assign \DFF_1027.CK  = CK;
  assign \DFF_1028.CK  = CK;
  assign \DFF_1029.CK  = CK;
  assign \DFF_1029.D  = \DFF_953.Q ;
  assign \DFF_103.CK  = CK;
  assign \DFF_1030.CK  = CK;
  assign \DFF_1030.D  = \DFF_1029.Q ;
  assign \DFF_1031.CK  = CK;
  assign \DFF_1031.D  = \DFF_954.Q ;
  assign \DFF_1032.CK  = CK;
  assign \DFF_1032.D  = \DFF_1031.Q ;
  assign \DFF_1033.CK  = CK;
  assign \DFF_1033.D  = \DFF_955.Q ;
  assign \DFF_1034.CK  = CK;
  assign \DFF_1034.D  = \DFF_1033.Q ;
  assign \DFF_1035.CK  = CK;
  assign \DFF_1035.D  = \DFF_956.Q ;
  assign \DFF_1036.CK  = CK;
  assign \DFF_1036.D  = \DFF_1035.Q ;
  assign \DFF_1037.CK  = CK;
  assign \DFF_1037.D  = \DFF_957.Q ;
  assign \DFF_1038.CK  = CK;
  assign \DFF_1038.D  = \DFF_1037.Q ;
  assign \DFF_1039.CK  = CK;
  assign \DFF_1039.D  = \DFF_958.Q ;
  assign \DFF_104.CK  = CK;
  assign \DFF_1040.CK  = CK;
  assign \DFF_1040.D  = \DFF_1039.Q ;
  assign \DFF_1041.CK  = CK;
  assign \DFF_1041.D  = \DFF_959.Q ;
  assign \DFF_1042.CK  = CK;
  assign \DFF_1042.D  = \DFF_1041.Q ;
  assign \DFF_1043.CK  = CK;
  assign \DFF_1043.D  = \DFF_960.Q ;
  assign \DFF_1044.CK  = CK;
  assign \DFF_1044.D  = \DFF_1043.Q ;
  assign \DFF_1045.CK  = CK;
  assign \DFF_1045.D  = \DFF_961.Q ;
  assign \DFF_1046.CK  = CK;
  assign \DFF_1046.D  = \DFF_1045.Q ;
  assign \DFF_1047.CK  = CK;
  assign \DFF_1047.D  = \DFF_962.Q ;
  assign \DFF_1048.CK  = CK;
  assign \DFF_1048.D  = \DFF_1047.Q ;
  assign \DFF_1049.CK  = CK;
  assign \DFF_1049.D  = \DFF_963.Q ;
  assign \DFF_105.CK  = CK;
  assign \DFF_1050.CK  = CK;
  assign \DFF_1050.D  = \DFF_1049.Q ;
  assign \DFF_1051.CK  = CK;
  assign \DFF_1051.D  = \DFF_964.Q ;
  assign \DFF_1052.CK  = CK;
  assign \DFF_1052.D  = \DFF_1051.Q ;
  assign \DFF_1053.CK  = CK;
  assign \DFF_1053.D  = \DFF_1563.Q ;
  assign \DFF_1053.Q  = \DFF_1504.Q ;
  assign \DFF_1054.CK  = CK;
  assign \DFF_1054.D  = \DFF_1504.Q ;
  assign \DFF_1054.Q  = \DFF_1505.Q ;
  assign \DFF_1055.CK  = CK;
  assign \DFF_1055.D  = \DFF_1505.Q ;
  assign \DFF_1055.Q  = \DFF_1506.Q ;
  assign \DFF_1056.CK  = CK;
  assign \DFF_1056.D  = \DFF_1563.Q ;
  assign \DFF_1056.Q  = \DFF_1504.Q ;
  assign \DFF_1057.CK  = CK;
  assign \DFF_1057.D  = \DFF_1504.Q ;
  assign \DFF_1057.Q  = \DFF_1505.Q ;
  assign \DFF_1058.CK  = CK;
  assign \DFF_1058.D  = \DFF_1505.Q ;
  assign \DFF_1058.Q  = \DFF_1506.Q ;
  assign \DFF_1059.CK  = CK;
  assign \DFF_106.CK  = CK;
  assign \DFF_1060.CK  = CK;
  assign \DFF_1061.CK  = CK;
  assign \DFF_1062.CK  = CK;
  assign \DFF_1063.CK  = CK;
  assign \DFF_1063.D  = \DFF_1062.Q ;
  assign \DFF_1064.CK  = CK;
  assign \DFF_1064.D  = \DFF_1063.Q ;
  assign \DFF_1065.CK  = CK;
  assign \DFF_1065.D  = \DFF_1083.Q ;
  assign \DFF_1066.CK  = CK;
  assign \DFF_1066.D  = \DFF_1065.Q ;
  assign \DFF_1067.CK  = CK;
  assign \DFF_1067.D  = \DFF_1084.Q ;
  assign \DFF_1068.CK  = CK;
  assign \DFF_1068.D  = \DFF_1067.Q ;
  assign \DFF_1069.CK  = CK;
  assign \DFF_1069.D  = \DFF_1085.Q ;
  assign \DFF_107.CK  = CK;
  assign \DFF_1070.CK  = CK;
  assign \DFF_1070.D  = \DFF_1069.Q ;
  assign \DFF_1071.CK  = CK;
  assign \DFF_1071.D  = \DFF_1092.Q ;
  assign \DFF_1072.CK  = CK;
  assign \DFF_1072.D  = \DFF_1071.Q ;
  assign \DFF_1073.CK  = CK;
  assign \DFF_1073.D  = \DFF_1093.Q ;
  assign \DFF_1074.CK  = CK;
  assign \DFF_1074.D  = \DFF_1073.Q ;
  assign \DFF_1075.CK  = CK;
  assign \DFF_1075.D  = \DFF_1094.Q ;
  assign \DFF_1076.CK  = CK;
  assign \DFF_1076.D  = \DFF_1075.Q ;
  assign \DFF_1077.CK  = CK;
  assign \DFF_1077.D  = \DFF_3.Q ;
  assign \DFF_1077.Q  = \DFF_1427.Q ;
  assign \DFF_1078.CK  = CK;
  assign \DFF_1078.D  = \DFF_1427.Q ;
  assign \DFF_1078.Q  = \DFF_1428.Q ;
  assign \DFF_1079.CK  = CK;
  assign \DFF_1079.D  = \DFF_1428.Q ;
  assign \DFF_1079.Q  = \DFF_1429.Q ;
  assign \DFF_108.CK  = CK;
  assign \DFF_1080.CK  = CK;
  assign \DFF_1081.CK  = CK;
  assign \DFF_1082.CK  = CK;
  assign \DFF_1083.CK  = CK;
  assign \DFF_1084.CK  = CK;
  assign \DFF_1085.CK  = CK;
  assign \DFF_1086.CK  = CK;
  assign \DFF_1087.CK  = CK;
  assign \DFF_1088.CK  = CK;
  assign \DFF_1089.CK  = CK;
  assign \DFF_109.CK  = CK;
  assign \DFF_1090.CK  = CK;
  assign \DFF_1091.CK  = CK;
  assign \DFF_1092.CK  = CK;
  assign \DFF_1093.CK  = CK;
  assign \DFF_1094.CK  = CK;
  assign \DFF_1095.CK  = CK;
  assign \DFF_1096.CK  = CK;
  assign \DFF_1096.D  = \DFF_1095.Q ;
  assign \DFF_1097.CK  = CK;
  assign \DFF_1097.D  = \DFF_1096.Q ;
  assign \DFF_1098.CK  = CK;
  assign \DFF_1099.CK  = CK;
  assign \DFF_1099.D  = \DFF_1098.Q ;
  assign \DFF_11.CK  = CK;
  assign \DFF_110.CK  = CK;
  assign \DFF_1100.CK  = CK;
  assign \DFF_1101.CK  = CK;
  assign \DFF_1102.CK  = CK;
  assign \DFF_1102.D  = \DFF_1101.Q ;
  assign \DFF_1103.CK  = CK;
  assign \DFF_1104.CK  = CK;
  assign \DFF_1104.D  = \DFF_1103.Q ;
  assign \DFF_1105.CK  = CK;
  assign \DFF_1106.CK  = CK;
  assign \DFF_1107.CK  = CK;
  assign \DFF_1108.CK  = CK;
  assign \DFF_1109.CK  = CK;
  assign \DFF_111.CK  = CK;
  assign \DFF_1110.CK  = CK;
  assign \DFF_1111.CK  = CK;
  assign \DFF_1112.CK  = CK;
  assign \DFF_1113.CK  = CK;
  assign \DFF_1114.CK  = CK;
  assign \DFF_1115.CK  = CK;
  assign \DFF_1116.CK  = CK;
  assign \DFF_1117.CK  = CK;
  assign \DFF_1118.CK  = CK;
  assign \DFF_1119.CK  = CK;
  assign \DFF_112.CK  = CK;
  assign \DFF_1120.CK  = CK;
  assign \DFF_1121.CK  = CK;
  assign \DFF_1122.CK  = CK;
  assign \DFF_1123.CK  = CK;
  assign \DFF_1124.CK  = CK;
  assign \DFF_1125.CK  = CK;
  assign \DFF_1126.CK  = CK;
  assign \DFF_1127.CK  = CK;
  assign \DFF_1128.CK  = CK;
  assign \DFF_1129.CK  = CK;
  assign \DFF_113.CK  = CK;
  assign \DFF_1130.CK  = CK;
  assign \DFF_1131.CK  = CK;
  assign \DFF_1132.CK  = CK;
  assign \DFF_1132.D  = \DFF_1102.Q ;
  assign \DFF_1133.CK  = CK;
  assign \DFF_1134.CK  = CK;
  assign \DFF_1135.CK  = CK;
  assign \DFF_1136.CK  = CK;
  assign \DFF_1137.CK  = CK;
  assign \DFF_1138.CK  = CK;
  assign \DFF_1139.CK  = CK;
  assign \DFF_114.CK  = CK;
  assign \DFF_1140.CK  = CK;
  assign \DFF_1141.CK  = CK;
  assign \DFF_1142.CK  = CK;
  assign \DFF_1143.CK  = CK;
  assign \DFF_1143.D  = \DFF_1142.Q ;
  assign \DFF_1144.CK  = CK;
  assign \DFF_1145.CK  = CK;
  assign \DFF_1146.CK  = CK;
  assign \DFF_1147.CK  = CK;
  assign \DFF_1148.CK  = CK;
  assign \DFF_1149.CK  = CK;
  assign \DFF_115.CK  = CK;
  assign \DFF_1150.CK  = CK;
  assign \DFF_1151.CK  = CK;
  assign \DFF_1152.CK  = CK;
  assign \DFF_1153.CK  = CK;
  assign \DFF_1154.CK  = CK;
  assign \DFF_1154.D  = \DFF_1563.Q ;
  assign \DFF_1154.Q  = \DFF_1504.Q ;
  assign \DFF_1155.CK  = CK;
  assign \DFF_1155.D  = \DFF_1504.Q ;
  assign \DFF_1155.Q  = \DFF_1505.Q ;
  assign \DFF_1156.CK  = CK;
  assign \DFF_1156.D  = \DFF_1505.Q ;
  assign \DFF_1156.Q  = \DFF_1506.Q ;
  assign \DFF_1157.CK  = CK;
  assign \DFF_1158.CK  = CK;
  assign \DFF_1159.CK  = CK;
  assign \DFF_116.CK  = CK;
  assign \DFF_1160.CK  = CK;
  assign \DFF_1161.CK  = CK;
  assign \DFF_1162.CK  = CK;
  assign \DFF_1163.CK  = CK;
  assign \DFF_1164.CK  = CK;
  assign \DFF_1165.CK  = CK;
  assign \DFF_1166.CK  = CK;
  assign \DFF_1167.CK  = CK;
  assign \DFF_1168.CK  = CK;
  assign \DFF_1169.CK  = CK;
  assign \DFF_117.CK  = CK;
  assign \DFF_1170.CK  = CK;
  assign \DFF_1171.CK  = CK;
  assign \DFF_1172.CK  = CK;
  assign \DFF_1173.CK  = CK;
  assign \DFF_1174.CK  = CK;
  assign \DFF_1175.CK  = CK;
  assign \DFF_1176.CK  = CK;
  assign \DFF_1177.CK  = CK;
  assign \DFF_1178.CK  = CK;
  assign \DFF_1179.CK  = CK;
  assign \DFF_118.CK  = CK;
  assign \DFF_1180.CK  = CK;
  assign \DFF_1181.CK  = CK;
  assign \DFF_1182.CK  = CK;
  assign \DFF_1183.CK  = CK;
  assign \DFF_1184.CK  = CK;
  assign \DFF_1185.CK  = CK;
  assign \DFF_1186.CK  = CK;
  assign \DFF_1187.CK  = CK;
  assign \DFF_1188.CK  = CK;
  assign \DFF_1189.CK  = CK;
  assign \DFF_119.CK  = CK;
  assign \DFF_1190.CK  = CK;
  assign \DFF_1191.CK  = CK;
  assign \DFF_1192.CK  = CK;
  assign \DFF_1193.CK  = CK;
  assign \DFF_1194.CK  = CK;
  assign \DFF_1195.CK  = CK;
  assign \DFF_1196.CK  = CK;
  assign \DFF_1197.CK  = CK;
  assign \DFF_1198.CK  = CK;
  assign \DFF_1199.CK  = CK;
  assign \DFF_12.CK  = CK;
  assign \DFF_120.CK  = CK;
  assign \DFF_1200.CK  = CK;
  assign \DFF_1201.CK  = CK;
  assign \DFF_1202.CK  = CK;
  assign \DFF_1203.CK  = CK;
  assign \DFF_1204.CK  = CK;
  assign \DFF_1205.CK  = CK;
  assign \DFF_1206.CK  = CK;
  assign \DFF_1207.CK  = CK;
  assign \DFF_1208.CK  = CK;
  assign \DFF_1209.CK  = CK;
  assign \DFF_121.CK  = CK;
  assign \DFF_1210.CK  = CK;
  assign \DFF_1211.CK  = CK;
  assign \DFF_1211.D  = \DFF_3.Q ;
  assign \DFF_1211.Q  = \DFF_1427.Q ;
  assign \DFF_1212.CK  = CK;
  assign \DFF_1212.D  = \DFF_1427.Q ;
  assign \DFF_1212.Q  = \DFF_1428.Q ;
  assign \DFF_1213.CK  = CK;
  assign \DFF_1213.D  = \DFF_1428.Q ;
  assign \DFF_1213.Q  = \DFF_1429.Q ;
  assign \DFF_1214.CK  = CK;
  assign \DFF_1215.CK  = CK;
  assign \DFF_1216.CK  = CK;
  assign \DFF_1217.CK  = CK;
  assign \DFF_1218.CK  = CK;
  assign \DFF_1219.CK  = CK;
  assign \DFF_122.CK  = CK;
  assign \DFF_1220.CK  = CK;
  assign \DFF_1221.CK  = CK;
  assign \DFF_1222.CK  = CK;
  assign \DFF_1223.CK  = CK;
  assign \DFF_1224.CK  = CK;
  assign \DFF_1225.CK  = CK;
  assign \DFF_1226.CK  = CK;
  assign \DFF_1227.CK  = CK;
  assign \DFF_1228.CK  = CK;
  assign \DFF_1229.CK  = CK;
  assign \DFF_123.CK  = CK;
  assign \DFF_1230.CK  = CK;
  assign \DFF_1231.CK  = CK;
  assign \DFF_1232.CK  = CK;
  assign \DFF_1233.CK  = CK;
  assign \DFF_1234.CK  = CK;
  assign \DFF_1235.CK  = CK;
  assign \DFF_1236.CK  = CK;
  assign \DFF_1237.CK  = CK;
  assign \DFF_1238.CK  = CK;
  assign \DFF_1239.CK  = CK;
  assign \DFF_124.CK  = CK;
  assign \DFF_1240.CK  = CK;
  assign \DFF_1241.CK  = CK;
  assign \DFF_1242.CK  = CK;
  assign \DFF_1243.CK  = CK;
  assign \DFF_1244.CK  = CK;
  assign \DFF_1245.CK  = CK;
  assign \DFF_1246.CK  = CK;
  assign \DFF_1247.CK  = CK;
  assign \DFF_1248.CK  = CK;
  assign \DFF_1249.CK  = CK;
  assign \DFF_125.CK  = CK;
  assign \DFF_1250.CK  = CK;
  assign \DFF_1251.CK  = CK;
  assign \DFF_1252.CK  = CK;
  assign \DFF_1253.CK  = CK;
  assign \DFF_1254.CK  = CK;
  assign \DFF_1255.CK  = CK;
  assign \DFF_1256.CK  = CK;
  assign \DFF_1257.CK  = CK;
  assign \DFF_1258.CK  = CK;
  assign \DFF_1259.CK  = CK;
  assign \DFF_126.CK  = CK;
  assign \DFF_1260.CK  = CK;
  assign \DFF_1261.CK  = CK;
  assign \DFF_1262.CK  = CK;
  assign \DFF_1263.CK  = CK;
  assign \DFF_1264.CK  = CK;
  assign \DFF_1265.CK  = CK;
  assign \DFF_1266.CK  = CK;
  assign \DFF_1267.CK  = CK;
  assign \DFF_1268.CK  = CK;
  assign \DFF_1269.CK  = CK;
  assign \DFF_127.CK  = CK;
  assign \DFF_1270.CK  = CK;
  assign \DFF_1271.CK  = CK;
  assign \DFF_1272.CK  = CK;
  assign \DFF_1273.CK  = CK;
  assign \DFF_1274.CK  = CK;
  assign \DFF_1275.CK  = CK;
  assign \DFF_1276.CK  = CK;
  assign \DFF_1277.CK  = CK;
  assign \DFF_1278.CK  = CK;
  assign \DFF_1279.CK  = CK;
  assign \DFF_128.CK  = CK;
  assign \DFF_1280.CK  = CK;
  assign \DFF_1281.CK  = CK;
  assign \DFF_1282.CK  = CK;
  assign \DFF_1283.CK  = CK;
  assign \DFF_1284.CK  = CK;
  assign \DFF_1285.CK  = CK;
  assign \DFF_1286.CK  = CK;
  assign \DFF_1287.CK  = CK;
  assign \DFF_1288.CK  = CK;
  assign \DFF_1289.CK  = CK;
  assign \DFF_129.CK  = CK;
  assign \DFF_1290.CK  = CK;
  assign \DFF_1291.CK  = CK;
  assign \DFF_1292.CK  = CK;
  assign \DFF_1293.CK  = CK;
  assign \DFF_1294.CK  = CK;
  assign \DFF_1295.CK  = CK;
  assign \DFF_1296.CK  = CK;
  assign \DFF_1297.CK  = CK;
  assign \DFF_1297.D  = \DFF_1296.Q ;
  assign \DFF_1298.CK  = CK;
  assign \DFF_1298.D  = \DFF_1297.Q ;
  assign \DFF_1298.Q  = \DFF_1302.Q ;
  assign \DFF_1299.CK  = CK;
  assign \DFF_1299.D  = \DFF_3.Q ;
  assign \DFF_1299.Q  = \DFF_1427.Q ;
  assign \DFF_13.CK  = CK;
  assign \DFF_130.CK  = CK;
  assign \DFF_1300.CK  = CK;
  assign \DFF_1300.D  = \DFF_1427.Q ;
  assign \DFF_1300.Q  = \DFF_1428.Q ;
  assign \DFF_1301.CK  = CK;
  assign \DFF_1301.D  = \DFF_1428.Q ;
  assign \DFF_1301.Q  = \DFF_1429.Q ;
  assign \DFF_1302.CK  = CK;
  assign \DFF_1302.D  = \DFF_1297.Q ;
  assign \DFF_1303.CK  = CK;
  assign \DFF_1304.CK  = CK;
  assign \DFF_1305.CK  = CK;
  assign \DFF_1306.CK  = CK;
  assign \DFF_1307.CK  = CK;
  assign \DFF_1308.CK  = CK;
  assign \DFF_1309.CK  = CK;
  assign \DFF_131.CK  = CK;
  assign \DFF_1310.CK  = CK;
  assign \DFF_1311.CK  = CK;
  assign \DFF_1312.CK  = CK;
  assign \DFF_1313.CK  = CK;
  assign \DFF_1314.CK  = CK;
  assign \DFF_1315.CK  = CK;
  assign \DFF_1316.CK  = CK;
  assign \DFF_1317.CK  = CK;
  assign \DFF_1318.CK  = CK;
  assign \DFF_1319.CK  = CK;
  assign \DFF_132.CK  = CK;
  assign \DFF_132.D  = \DFF_152.D ;
  assign \DFF_132.Q  = \DFF_152.Q ;
  assign \DFF_1320.CK  = CK;
  assign \DFF_1321.CK  = CK;
  assign \DFF_1322.CK  = CK;
  assign \DFF_1323.CK  = CK;
  assign \DFF_1324.CK  = CK;
  assign \DFF_1325.CK  = CK;
  assign \DFF_1326.CK  = CK;
  assign \DFF_1327.CK  = CK;
  assign \DFF_1328.CK  = CK;
  assign \DFF_1329.CK  = CK;
  assign \DFF_133.CK  = CK;
  assign \DFF_133.D  = \DFF_151.D ;
  assign \DFF_133.Q  = \DFF_151.Q ;
  assign \DFF_1330.CK  = CK;
  assign \DFF_1331.CK  = CK;
  assign \DFF_1332.CK  = CK;
  assign \DFF_1333.CK  = CK;
  assign \DFF_1334.CK  = CK;
  assign \DFF_1335.CK  = CK;
  assign \DFF_1336.CK  = CK;
  assign \DFF_1337.CK  = CK;
  assign \DFF_1338.CK  = CK;
  assign \DFF_1339.CK  = CK;
  assign \DFF_134.CK  = CK;
  assign \DFF_134.D  = \DFF_150.D ;
  assign \DFF_134.Q  = \DFF_150.Q ;
  assign \DFF_1340.CK  = CK;
  assign \DFF_1341.CK  = CK;
  assign \DFF_1342.CK  = CK;
  assign \DFF_1343.CK  = CK;
  assign \DFF_1344.CK  = CK;
  assign \DFF_1345.CK  = CK;
  assign \DFF_1346.CK  = CK;
  assign \DFF_1347.CK  = CK;
  assign \DFF_1348.CK  = CK;
  assign \DFF_1349.CK  = CK;
  assign \DFF_1349.D  = \DFF_1348.Q ;
  assign \DFF_135.CK  = CK;
  assign \DFF_135.D  = \DFF_156.D ;
  assign \DFF_135.Q  = \DFF_156.Q ;
  assign \DFF_1350.CK  = CK;
  assign \DFF_1351.CK  = CK;
  assign \DFF_1351.D  = \DFF_1350.Q ;
  assign \DFF_1352.CK  = CK;
  assign \DFF_1353.CK  = CK;
  assign \DFF_1353.D  = \DFF_1352.Q ;
  assign \DFF_1354.CK  = CK;
  assign \DFF_1355.CK  = CK;
  assign \DFF_1355.D  = \DFF_1354.Q ;
  assign \DFF_1356.CK  = CK;
  assign \DFF_1357.CK  = CK;
  assign \DFF_1357.D  = \DFF_1356.Q ;
  assign \DFF_1358.CK  = CK;
  assign \DFF_1359.CK  = CK;
  assign \DFF_1359.D  = \DFF_1358.Q ;
  assign \DFF_136.CK  = CK;
  assign \DFF_136.D  = \DFF_159.D ;
  assign \DFF_136.Q  = \DFF_159.Q ;
  assign \DFF_1360.CK  = CK;
  assign \DFF_1361.CK  = CK;
  assign \DFF_1361.D  = \DFF_1360.Q ;
  assign \DFF_1362.CK  = CK;
  assign \DFF_1363.CK  = CK;
  assign \DFF_1363.D  = \DFF_1362.Q ;
  assign \DFF_1364.CK  = CK;
  assign \DFF_1364.D  = \DFF_91.Q ;
  assign \DFF_1365.CK  = CK;
  assign \DFF_1365.D  = \DFF_1364.Q ;
  assign \DFF_1366.CK  = CK;
  assign \DFF_1367.CK  = CK;
  assign \DFF_1368.CK  = CK;
  assign \DFF_1369.CK  = CK;
  assign \DFF_137.CK  = CK;
  assign \DFF_137.D  = \DFF_158.D ;
  assign \DFF_137.Q  = \DFF_158.Q ;
  assign \DFF_1370.CK  = CK;
  assign \DFF_1371.CK  = CK;
  assign \DFF_1372.CK  = CK;
  assign \DFF_1373.CK  = CK;
  assign \DFF_1374.CK  = CK;
  assign \DFF_1375.CK  = CK;
  assign \DFF_1376.CK  = CK;
  assign \DFF_1377.CK  = CK;
  assign \DFF_1378.CK  = CK;
  assign \DFF_1379.CK  = CK;
  assign \DFF_1379.D  = \DFF_1303.Q ;
  assign \DFF_138.CK  = CK;
  assign \DFF_138.D  = \DFF_157.D ;
  assign \DFF_138.Q  = \DFF_157.Q ;
  assign \DFF_1380.CK  = CK;
  assign \DFF_1380.D  = \DFF_1379.Q ;
  assign \DFF_1381.CK  = CK;
  assign \DFF_1381.D  = \DFF_1304.Q ;
  assign \DFF_1382.CK  = CK;
  assign \DFF_1382.D  = \DFF_1381.Q ;
  assign \DFF_1383.CK  = CK;
  assign \DFF_1383.D  = \DFF_1305.Q ;
  assign \DFF_1384.CK  = CK;
  assign \DFF_1384.D  = \DFF_1383.Q ;
  assign \DFF_1385.CK  = CK;
  assign \DFF_1385.D  = \DFF_1306.Q ;
  assign \DFF_1386.CK  = CK;
  assign \DFF_1386.D  = \DFF_1385.Q ;
  assign \DFF_1387.CK  = CK;
  assign \DFF_1387.D  = \DFF_1307.Q ;
  assign \DFF_1388.CK  = CK;
  assign \DFF_1388.D  = \DFF_1387.Q ;
  assign \DFF_1389.CK  = CK;
  assign \DFF_1389.D  = \DFF_1308.Q ;
  assign \DFF_139.CK  = CK;
  assign \DFF_139.D  = \DFF_160.D ;
  assign \DFF_139.Q  = \DFF_160.Q ;
  assign \DFF_1390.CK  = CK;
  assign \DFF_1390.D  = \DFF_1389.Q ;
  assign \DFF_1391.CK  = CK;
  assign \DFF_1391.D  = \DFF_1309.Q ;
  assign \DFF_1392.CK  = CK;
  assign \DFF_1392.D  = \DFF_1391.Q ;
  assign \DFF_1393.CK  = CK;
  assign \DFF_1393.D  = \DFF_1310.Q ;
  assign \DFF_1394.CK  = CK;
  assign \DFF_1394.D  = \DFF_1393.Q ;
  assign \DFF_1395.CK  = CK;
  assign \DFF_1395.D  = \DFF_1311.Q ;
  assign \DFF_1396.CK  = CK;
  assign \DFF_1396.D  = \DFF_1395.Q ;
  assign \DFF_1397.CK  = CK;
  assign \DFF_1397.D  = \DFF_1312.Q ;
  assign \DFF_1398.CK  = CK;
  assign \DFF_1398.D  = \DFF_1397.Q ;
  assign \DFF_1399.CK  = CK;
  assign \DFF_1399.D  = \DFF_1313.Q ;
  assign \DFF_14.CK  = CK;
  assign \DFF_140.CK  = CK;
  assign \DFF_140.D  = \DFF_158.D ;
  assign \DFF_140.Q  = \DFF_158.Q ;
  assign \DFF_1400.CK  = CK;
  assign \DFF_1400.D  = \DFF_1399.Q ;
  assign \DFF_1401.CK  = CK;
  assign \DFF_1401.D  = \DFF_1314.Q ;
  assign \DFF_1402.CK  = CK;
  assign \DFF_1402.D  = \DFF_1401.Q ;
  assign \DFF_1403.CK  = CK;
  assign \DFF_1403.D  = \DFF_1563.Q ;
  assign \DFF_1403.Q  = \DFF_1504.Q ;
  assign \DFF_1404.CK  = CK;
  assign \DFF_1404.D  = \DFF_1504.Q ;
  assign \DFF_1404.Q  = \DFF_1505.Q ;
  assign \DFF_1405.CK  = CK;
  assign \DFF_1405.D  = \DFF_1505.Q ;
  assign \DFF_1405.Q  = \DFF_1506.Q ;
  assign \DFF_1406.CK  = CK;
  assign \DFF_1406.D  = \DFF_1563.Q ;
  assign \DFF_1406.Q  = \DFF_1504.Q ;
  assign \DFF_1407.CK  = CK;
  assign \DFF_1407.D  = \DFF_1504.Q ;
  assign \DFF_1407.Q  = \DFF_1505.Q ;
  assign \DFF_1408.CK  = CK;
  assign \DFF_1408.D  = \DFF_1505.Q ;
  assign \DFF_1408.Q  = \DFF_1506.Q ;
  assign \DFF_1409.CK  = CK;
  assign \DFF_141.CK  = CK;
  assign \DFF_1410.CK  = CK;
  assign \DFF_1411.CK  = CK;
  assign \DFF_1412.CK  = CK;
  assign \DFF_1413.CK  = CK;
  assign \DFF_1413.D  = \DFF_1412.Q ;
  assign \DFF_1414.CK  = CK;
  assign \DFF_1414.D  = \DFF_1413.Q ;
  assign \DFF_1415.CK  = CK;
  assign \DFF_1415.D  = \DFF_1433.Q ;
  assign \DFF_1416.CK  = CK;
  assign \DFF_1416.D  = \DFF_1415.Q ;
  assign \DFF_1417.CK  = CK;
  assign \DFF_1417.D  = \DFF_1434.Q ;
  assign \DFF_1418.CK  = CK;
  assign \DFF_1418.D  = \DFF_1417.Q ;
  assign \DFF_1419.CK  = CK;
  assign \DFF_1419.D  = \DFF_1435.Q ;
  assign \DFF_142.CK  = CK;
  assign \DFF_142.D  = \DFF_156.D ;
  assign \DFF_142.Q  = \DFF_156.Q ;
  assign \DFF_1420.CK  = CK;
  assign \DFF_1420.D  = \DFF_1419.Q ;
  assign \DFF_1421.CK  = CK;
  assign \DFF_1421.D  = \DFF_1442.Q ;
  assign \DFF_1422.CK  = CK;
  assign \DFF_1422.D  = \DFF_1421.Q ;
  assign \DFF_1423.CK  = CK;
  assign \DFF_1423.D  = \DFF_1443.Q ;
  assign \DFF_1424.CK  = CK;
  assign \DFF_1424.D  = \DFF_1423.Q ;
  assign \DFF_1425.CK  = CK;
  assign \DFF_1425.D  = \DFF_1444.Q ;
  assign \DFF_1426.CK  = CK;
  assign \DFF_1426.D  = \DFF_1425.Q ;
  assign \DFF_1427.CK  = CK;
  assign \DFF_1427.D  = \DFF_3.Q ;
  assign \DFF_1428.CK  = CK;
  assign \DFF_1428.D  = \DFF_1427.Q ;
  assign \DFF_1429.CK  = CK;
  assign \DFF_1429.D  = \DFF_1428.Q ;
  assign \DFF_143.CK  = CK;
  assign \DFF_143.D  = \DFF_150.D ;
  assign \DFF_143.Q  = \DFF_150.Q ;
  assign \DFF_1430.CK  = CK;
  assign \DFF_1431.CK  = CK;
  assign \DFF_1432.CK  = CK;
  assign \DFF_1433.CK  = CK;
  assign \DFF_1434.CK  = CK;
  assign \DFF_1435.CK  = CK;
  assign \DFF_1436.CK  = CK;
  assign \DFF_1437.CK  = CK;
  assign \DFF_1438.CK  = CK;
  assign \DFF_1439.CK  = CK;
  assign \DFF_144.CK  = CK;
  assign \DFF_1440.CK  = CK;
  assign \DFF_1441.CK  = CK;
  assign \DFF_1442.CK  = CK;
  assign \DFF_1443.CK  = CK;
  assign \DFF_1444.CK  = CK;
  assign \DFF_1445.CK  = CK;
  assign \DFF_1446.CK  = CK;
  assign \DFF_1446.D  = \DFF_1445.Q ;
  assign \DFF_1447.CK  = CK;
  assign \DFF_1447.D  = \DFF_1446.Q ;
  assign \DFF_1448.CK  = CK;
  assign \DFF_1449.CK  = CK;
  assign \DFF_1449.D  = \DFF_1448.Q ;
  assign \DFF_145.CK  = CK;
  assign \DFF_145.D  = \DFF_152.D ;
  assign \DFF_145.Q  = \DFF_152.Q ;
  assign \DFF_1450.CK  = CK;
  assign \DFF_1451.CK  = CK;
  assign \DFF_1452.CK  = CK;
  assign \DFF_1452.D  = \DFF_1451.Q ;
  assign \DFF_1453.CK  = CK;
  assign \DFF_1454.CK  = CK;
  assign \DFF_1454.D  = \DFF_1453.Q ;
  assign \DFF_1455.CK  = CK;
  assign \DFF_1456.CK  = CK;
  assign \DFF_1457.CK  = CK;
  assign \DFF_1458.CK  = CK;
  assign \DFF_1459.CK  = CK;
  assign \DFF_146.CK  = CK;
  assign \DFF_1460.CK  = CK;
  assign \DFF_1461.CK  = CK;
  assign \DFF_1462.CK  = CK;
  assign \DFF_1463.CK  = CK;
  assign \DFF_1464.CK  = CK;
  assign \DFF_1465.CK  = CK;
  assign \DFF_1466.CK  = CK;
  assign \DFF_1467.CK  = CK;
  assign \DFF_1468.CK  = CK;
  assign \DFF_1469.CK  = CK;
  assign \DFF_147.CK  = CK;
  assign \DFF_147.D  = \DFF_158.D ;
  assign \DFF_147.Q  = \DFF_158.Q ;
  assign \DFF_1470.CK  = CK;
  assign \DFF_1471.CK  = CK;
  assign \DFF_1472.CK  = CK;
  assign \DFF_1473.CK  = CK;
  assign \DFF_1474.CK  = CK;
  assign \DFF_1475.CK  = CK;
  assign \DFF_1476.CK  = CK;
  assign \DFF_1477.CK  = CK;
  assign \DFF_1478.CK  = CK;
  assign \DFF_1479.CK  = CK;
  assign \DFF_148.CK  = CK;
  assign \DFF_148.D  = \DFF_159.D ;
  assign \DFF_148.Q  = \DFF_159.Q ;
  assign \DFF_1480.CK  = CK;
  assign \DFF_1481.CK  = CK;
  assign \DFF_1482.CK  = CK;
  assign \DFF_1482.D  = \DFF_1452.Q ;
  assign \DFF_1483.CK  = CK;
  assign \DFF_1484.CK  = CK;
  assign \DFF_1485.CK  = CK;
  assign \DFF_1486.CK  = CK;
  assign \DFF_1487.CK  = CK;
  assign \DFF_1488.CK  = CK;
  assign \DFF_1489.CK  = CK;
  assign \DFF_149.CK  = CK;
  assign \DFF_149.D  = \DFF_156.D ;
  assign \DFF_149.Q  = \DFF_156.Q ;
  assign \DFF_1490.CK  = CK;
  assign \DFF_1491.CK  = CK;
  assign \DFF_1492.CK  = CK;
  assign \DFF_1493.CK  = CK;
  assign \DFF_1493.D  = \DFF_1492.Q ;
  assign \DFF_1494.CK  = CK;
  assign \DFF_1495.CK  = CK;
  assign \DFF_1496.CK  = CK;
  assign \DFF_1497.CK  = CK;
  assign \DFF_1498.CK  = CK;
  assign \DFF_1499.CK  = CK;
  assign \DFF_15.CK  = CK;
  assign \DFF_150.CK  = CK;
  assign \DFF_1500.CK  = CK;
  assign \DFF_1501.CK  = CK;
  assign \DFF_1502.CK  = CK;
  assign \DFF_1503.CK  = CK;
  assign \DFF_1504.CK  = CK;
  assign \DFF_1504.D  = \DFF_1563.Q ;
  assign \DFF_1505.CK  = CK;
  assign \DFF_1505.D  = \DFF_1504.Q ;
  assign \DFF_1506.CK  = CK;
  assign \DFF_1506.D  = \DFF_1505.Q ;
  assign \DFF_1507.CK  = CK;
  assign \DFF_1508.CK  = CK;
  assign \DFF_1509.CK  = CK;
  assign \DFF_151.CK  = CK;
  assign \DFF_1510.CK  = CK;
  assign \DFF_1511.CK  = CK;
  assign \DFF_1512.CK  = CK;
  assign \DFF_1513.CK  = CK;
  assign \DFF_1514.CK  = CK;
  assign \DFF_1515.CK  = CK;
  assign \DFF_1516.CK  = CK;
  assign \DFF_1517.CK  = CK;
  assign \DFF_1518.CK  = CK;
  assign \DFF_1519.CK  = CK;
  assign \DFF_152.CK  = CK;
  assign \DFF_1520.CK  = CK;
  assign \DFF_1521.CK  = CK;
  assign \DFF_1522.CK  = CK;
  assign \DFF_1523.CK  = CK;
  assign \DFF_1524.CK  = CK;
  assign \DFF_1525.CK  = CK;
  assign \DFF_1526.CK  = CK;
  assign \DFF_1527.CK  = CK;
  assign \DFF_1528.CK  = CK;
  assign \DFF_1529.CK  = CK;
  assign \DFF_153.CK  = CK;
  assign \DFF_153.D  = \DFF_157.D ;
  assign \DFF_153.Q  = \DFF_157.Q ;
  assign \DFF_1530.CK  = CK;
  assign \DFF_1531.CK  = CK;
  assign \DFF_1532.CK  = CK;
  assign \DFF_1533.CK  = CK;
  assign \DFF_1534.CK  = CK;
  assign \DFF_1535.CK  = CK;
  assign \DFF_1536.CK  = CK;
  assign \DFF_1537.CK  = CK;
  assign \DFF_1538.CK  = CK;
  assign \DFF_1539.CK  = CK;
  assign \DFF_154.CK  = CK;
  assign \DFF_154.D  = \DFF_158.D ;
  assign \DFF_154.Q  = \DFF_158.Q ;
  assign \DFF_1540.CK  = CK;
  assign \DFF_1541.CK  = CK;
  assign \DFF_1542.CK  = CK;
  assign \DFF_1543.CK  = CK;
  assign \DFF_1544.CK  = CK;
  assign \DFF_1545.CK  = CK;
  assign \DFF_1546.CK  = CK;
  assign \DFF_1547.CK  = CK;
  assign \DFF_1548.CK  = CK;
  assign \DFF_1549.CK  = CK;
  assign \DFF_155.CK  = CK;
  assign \DFF_155.D  = \DFF_159.D ;
  assign \DFF_155.Q  = \DFF_159.Q ;
  assign \DFF_1550.CK  = CK;
  assign \DFF_1551.CK  = CK;
  assign \DFF_1552.CK  = CK;
  assign \DFF_1553.CK  = CK;
  assign \DFF_1554.CK  = CK;
  assign \DFF_1555.CK  = CK;
  assign \DFF_1556.CK  = CK;
  assign \DFF_1557.CK  = CK;
  assign \DFF_1558.CK  = CK;
  assign \DFF_1559.CK  = CK;
  assign \DFF_156.CK  = CK;
  assign \DFF_1560.CK  = CK;
  assign \DFF_1561.CK  = CK;
  assign \DFF_1562.CK  = CK;
  assign \DFF_1563.CK  = CK;
  assign \DFF_1564.CK  = CK;
  assign \DFF_1565.CK  = CK;
  assign \DFF_1566.CK  = CK;
  assign \DFF_1567.CK  = CK;
  assign \DFF_1568.CK  = CK;
  assign \DFF_1569.CK  = CK;
  assign \DFF_157.CK  = CK;
  assign \DFF_1570.CK  = CK;
  assign \DFF_1571.CK  = CK;
  assign \DFF_1572.CK  = CK;
  assign \DFF_1573.CK  = CK;
  assign \DFF_1574.CK  = CK;
  assign \DFF_1575.CK  = CK;
  assign \DFF_1576.CK  = CK;
  assign \DFF_1577.CK  = CK;
  assign \DFF_1578.CK  = CK;
  assign \DFF_1579.CK  = CK;
  assign \DFF_158.CK  = CK;
  assign \DFF_1580.CK  = CK;
  assign \DFF_1581.CK  = CK;
  assign \DFF_1582.CK  = CK;
  assign \DFF_1583.CK  = CK;
  assign \DFF_1584.CK  = CK;
  assign \DFF_1585.CK  = CK;
  assign \DFF_1586.CK  = CK;
  assign \DFF_1587.CK  = CK;
  assign \DFF_1588.CK  = CK;
  assign \DFF_1589.CK  = CK;
  assign \DFF_159.CK  = CK;
  assign \DFF_1590.CK  = CK;
  assign \DFF_1591.CK  = CK;
  assign \DFF_1592.CK  = CK;
  assign \DFF_1593.CK  = CK;
  assign \DFF_1594.CK  = CK;
  assign \DFF_1595.CK  = CK;
  assign \DFF_1596.CK  = CK;
  assign \DFF_1597.CK  = CK;
  assign \DFF_1598.CK  = CK;
  assign \DFF_1599.CK  = CK;
  assign \DFF_16.CK  = CK;
  assign \DFF_160.CK  = CK;
  assign \DFF_1600.CK  = CK;
  assign \DFF_1601.CK  = CK;
  assign \DFF_1602.CK  = CK;
  assign \DFF_1603.CK  = CK;
  assign \DFF_1604.CK  = CK;
  assign \DFF_1605.CK  = CK;
  assign \DFF_1606.CK  = CK;
  assign \DFF_1607.CK  = CK;
  assign \DFF_1608.CK  = CK;
  assign \DFF_1609.CK  = CK;
  assign \DFF_161.CK  = CK;
  assign \DFF_161.D  = \DFF_3.Q ;
  assign \DFF_161.Q  = \DFF_1427.Q ;
  assign \DFF_1610.CK  = CK;
  assign \DFF_1611.CK  = CK;
  assign \DFF_1611.D  = g3234;
  assign \DFF_1612.CK  = CK;
  assign \DFF_1612.D  = \DFF_1611.Q ;
  assign \DFF_1613.CK  = CK;
  assign \DFF_1614.CK  = CK;
  assign \DFF_1615.CK  = CK;
  assign \DFF_1616.CK  = CK;
  assign \DFF_1617.CK  = CK;
  assign \DFF_1618.CK  = CK;
  assign \DFF_1619.CK  = CK;
  assign \DFF_162.CK  = CK;
  assign \DFF_162.D  = \DFF_1427.Q ;
  assign \DFF_162.Q  = \DFF_1428.Q ;
  assign \DFF_1620.CK  = CK;
  assign \DFF_1621.CK  = CK;
  assign \DFF_1622.CK  = CK;
  assign \DFF_1623.CK  = CK;
  assign \DFF_1624.CK  = CK;
  assign \DFF_1625.CK  = CK;
  assign \DFF_1626.CK  = CK;
  assign \DFF_1627.CK  = CK;
  assign \DFF_1628.CK  = CK;
  assign \DFF_1629.CK  = CK;
  assign \DFF_163.CK  = CK;
  assign \DFF_163.D  = \DFF_1428.Q ;
  assign \DFF_163.Q  = \DFF_1429.Q ;
  assign \DFF_1630.CK  = CK;
  assign \DFF_1631.CK  = CK;
  assign \DFF_1632.CK  = CK;
  assign \DFF_1633.CK  = CK;
  assign \DFF_1634.CK  = CK;
  assign \DFF_1635.CK  = CK;
  assign \DFF_164.CK  = CK;
  assign \DFF_165.CK  = CK;
  assign \DFF_166.CK  = CK;
  assign \DFF_167.CK  = CK;
  assign \DFF_168.CK  = CK;
  assign \DFF_169.CK  = CK;
  assign \DFF_17.CK  = CK;
  assign \DFF_17.D  = g51;
  assign \DFF_170.CK  = CK;
  assign \DFF_171.CK  = CK;
  assign \DFF_172.CK  = CK;
  assign \DFF_173.CK  = CK;
  assign \DFF_174.CK  = CK;
  assign \DFF_175.CK  = CK;
  assign \DFF_176.CK  = CK;
  assign \DFF_177.CK  = CK;
  assign \DFF_178.CK  = CK;
  assign \DFF_179.CK  = CK;
  assign \DFF_18.CK  = CK;
  assign \DFF_18.D  = \DFF_17.Q ;
  assign \DFF_180.CK  = CK;
  assign \DFF_181.CK  = CK;
  assign \DFF_182.CK  = CK;
  assign \DFF_183.CK  = CK;
  assign \DFF_184.CK  = CK;
  assign \DFF_185.CK  = CK;
  assign \DFF_186.CK  = CK;
  assign \DFF_187.CK  = CK;
  assign \DFF_188.CK  = CK;
  assign \DFF_189.CK  = CK;
  assign \DFF_19.CK  = CK;
  assign \DFF_190.CK  = CK;
  assign \DFF_191.CK  = CK;
  assign \DFF_192.CK  = CK;
  assign \DFF_193.CK  = CK;
  assign \DFF_194.CK  = CK;
  assign \DFF_195.CK  = CK;
  assign \DFF_196.CK  = CK;
  assign \DFF_197.CK  = CK;
  assign \DFF_198.CK  = CK;
  assign \DFF_199.CK  = CK;
  assign \DFF_2.CK  = CK;
  assign \DFF_20.CK  = CK;
  assign \DFF_20.D  = g3212;
  assign \DFF_200.CK  = CK;
  assign \DFF_201.CK  = CK;
  assign \DFF_202.CK  = CK;
  assign \DFF_203.CK  = CK;
  assign \DFF_204.CK  = CK;
  assign \DFF_205.CK  = CK;
  assign \DFF_206.CK  = CK;
  assign \DFF_207.CK  = CK;
  assign \DFF_208.CK  = CK;
  assign \DFF_209.CK  = CK;
  assign \DFF_21.CK  = CK;
  assign \DFF_21.D  = g3228;
  assign \DFF_210.CK  = CK;
  assign \DFF_211.CK  = CK;
  assign \DFF_212.CK  = CK;
  assign \DFF_213.CK  = CK;
  assign \DFF_214.CK  = CK;
  assign \DFF_215.CK  = CK;
  assign \DFF_216.CK  = CK;
  assign \DFF_217.CK  = CK;
  assign \DFF_218.CK  = CK;
  assign \DFF_219.CK  = CK;
  assign \DFF_22.CK  = CK;
  assign \DFF_22.D  = g3227;
  assign \DFF_220.CK  = CK;
  assign \DFF_221.CK  = CK;
  assign \DFF_222.CK  = CK;
  assign \DFF_223.CK  = CK;
  assign \DFF_224.CK  = CK;
  assign \DFF_225.CK  = CK;
  assign \DFF_226.CK  = CK;
  assign \DFF_227.CK  = CK;
  assign \DFF_228.CK  = CK;
  assign \DFF_229.CK  = CK;
  assign \DFF_23.CK  = CK;
  assign \DFF_23.D  = g3226;
  assign \DFF_230.CK  = CK;
  assign \DFF_231.CK  = CK;
  assign \DFF_232.CK  = CK;
  assign \DFF_233.CK  = CK;
  assign \DFF_234.CK  = CK;
  assign \DFF_235.CK  = CK;
  assign \DFF_236.CK  = CK;
  assign \DFF_237.CK  = CK;
  assign \DFF_238.CK  = CK;
  assign \DFF_239.CK  = CK;
  assign \DFF_24.CK  = CK;
  assign \DFF_24.D  = g3225;
  assign \DFF_240.CK  = CK;
  assign \DFF_241.CK  = CK;
  assign \DFF_242.CK  = CK;
  assign \DFF_243.CK  = CK;
  assign \DFF_244.CK  = CK;
  assign \DFF_245.CK  = CK;
  assign \DFF_246.CK  = CK;
  assign \DFF_246.D  = \DFF_1296.D ;
  assign \DFF_246.Q  = \DFF_1296.Q ;
  assign \DFF_247.CK  = CK;
  assign \DFF_247.D  = \DFF_1296.Q ;
  assign \DFF_247.Q  = \DFF_1297.Q ;
  assign \DFF_248.CK  = CK;
  assign \DFF_248.D  = \DFF_1297.Q ;
  assign \DFF_248.Q  = \DFF_1302.Q ;
  assign \DFF_249.CK  = CK;
  assign \DFF_249.D  = \DFF_3.Q ;
  assign \DFF_249.Q  = \DFF_1427.Q ;
  assign \DFF_25.CK  = CK;
  assign \DFF_25.D  = g3224;
  assign \DFF_250.CK  = CK;
  assign \DFF_250.D  = \DFF_1427.Q ;
  assign \DFF_250.Q  = \DFF_1428.Q ;
  assign \DFF_251.CK  = CK;
  assign \DFF_251.D  = \DFF_1428.Q ;
  assign \DFF_251.Q  = \DFF_1429.Q ;
  assign \DFF_252.CK  = CK;
  assign \DFF_252.D  = \DFF_1297.Q ;
  assign \DFF_252.Q  = \DFF_1302.Q ;
  assign \DFF_253.CK  = CK;
  assign \DFF_254.CK  = CK;
  assign \DFF_255.CK  = CK;
  assign \DFF_256.CK  = CK;
  assign \DFF_257.CK  = CK;
  assign \DFF_258.CK  = CK;
  assign \DFF_259.CK  = CK;
  assign \DFF_26.CK  = CK;
  assign \DFF_26.D  = g3223;
  assign \DFF_260.CK  = CK;
  assign \DFF_261.CK  = CK;
  assign \DFF_262.CK  = CK;
  assign \DFF_263.CK  = CK;
  assign \DFF_264.CK  = CK;
  assign \DFF_265.CK  = CK;
  assign \DFF_266.CK  = CK;
  assign \DFF_267.CK  = CK;
  assign \DFF_268.CK  = CK;
  assign \DFF_269.CK  = CK;
  assign \DFF_27.CK  = CK;
  assign \DFF_27.D  = g3222;
  assign \DFF_270.CK  = CK;
  assign \DFF_271.CK  = CK;
  assign \DFF_272.CK  = CK;
  assign \DFF_273.CK  = CK;
  assign \DFF_274.CK  = CK;
  assign \DFF_275.CK  = CK;
  assign \DFF_276.CK  = CK;
  assign \DFF_277.CK  = CK;
  assign \DFF_278.CK  = CK;
  assign \DFF_279.CK  = CK;
  assign \DFF_28.CK  = CK;
  assign \DFF_28.D  = g3221;
  assign \DFF_280.CK  = CK;
  assign \DFF_281.CK  = CK;
  assign \DFF_282.CK  = CK;
  assign \DFF_283.CK  = CK;
  assign \DFF_284.CK  = CK;
  assign \DFF_285.CK  = CK;
  assign \DFF_286.CK  = CK;
  assign \DFF_287.CK  = CK;
  assign \DFF_288.CK  = CK;
  assign \DFF_289.CK  = CK;
  assign \DFF_29.CK  = CK;
  assign \DFF_29.D  = g3232;
  assign \DFF_290.CK  = CK;
  assign \DFF_291.CK  = CK;
  assign \DFF_292.CK  = CK;
  assign \DFF_293.CK  = CK;
  assign \DFF_294.CK  = CK;
  assign \DFF_295.CK  = CK;
  assign \DFF_296.CK  = CK;
  assign \DFF_297.CK  = CK;
  assign \DFF_298.CK  = CK;
  assign \DFF_299.CK  = CK;
  assign \DFF_299.D  = \DFF_298.Q ;
  assign \DFF_3.CK  = CK;
  assign \DFF_30.CK  = CK;
  assign \DFF_30.D  = g3220;
  assign \DFF_300.CK  = CK;
  assign \DFF_301.CK  = CK;
  assign \DFF_301.D  = \DFF_300.Q ;
  assign \DFF_302.CK  = CK;
  assign \DFF_303.CK  = CK;
  assign \DFF_303.D  = \DFF_302.Q ;
  assign \DFF_304.CK  = CK;
  assign \DFF_305.CK  = CK;
  assign \DFF_305.D  = \DFF_304.Q ;
  assign \DFF_306.CK  = CK;
  assign \DFF_307.CK  = CK;
  assign \DFF_307.D  = \DFF_306.Q ;
  assign \DFF_308.CK  = CK;
  assign \DFF_309.CK  = CK;
  assign \DFF_309.D  = \DFF_308.Q ;
  assign \DFF_31.CK  = CK;
  assign \DFF_31.D  = g3219;
  assign \DFF_310.CK  = CK;
  assign \DFF_311.CK  = CK;
  assign \DFF_311.D  = \DFF_310.Q ;
  assign \DFF_312.CK  = CK;
  assign \DFF_313.CK  = CK;
  assign \DFF_313.D  = \DFF_312.Q ;
  assign \DFF_314.CK  = CK;
  assign \DFF_314.D  = \DFF_82.Q ;
  assign \DFF_315.CK  = CK;
  assign \DFF_315.D  = \DFF_314.Q ;
  assign \DFF_316.CK  = CK;
  assign \DFF_317.CK  = CK;
  assign \DFF_318.CK  = CK;
  assign \DFF_319.CK  = CK;
  assign \DFF_32.CK  = CK;
  assign \DFF_32.D  = g3218;
  assign \DFF_320.CK  = CK;
  assign \DFF_321.CK  = CK;
  assign \DFF_322.CK  = CK;
  assign \DFF_323.CK  = CK;
  assign \DFF_324.CK  = CK;
  assign \DFF_325.CK  = CK;
  assign \DFF_326.CK  = CK;
  assign \DFF_327.CK  = CK;
  assign \DFF_328.CK  = CK;
  assign \DFF_329.CK  = CK;
  assign \DFF_329.D  = \DFF_253.Q ;
  assign \DFF_33.CK  = CK;
  assign \DFF_33.D  = g3217;
  assign \DFF_330.CK  = CK;
  assign \DFF_330.D  = \DFF_329.Q ;
  assign \DFF_331.CK  = CK;
  assign \DFF_331.D  = \DFF_254.Q ;
  assign \DFF_332.CK  = CK;
  assign \DFF_332.D  = \DFF_331.Q ;
  assign \DFF_333.CK  = CK;
  assign \DFF_333.D  = \DFF_255.Q ;
  assign \DFF_334.CK  = CK;
  assign \DFF_334.D  = \DFF_333.Q ;
  assign \DFF_335.CK  = CK;
  assign \DFF_335.D  = \DFF_256.Q ;
  assign \DFF_336.CK  = CK;
  assign \DFF_336.D  = \DFF_335.Q ;
  assign \DFF_337.CK  = CK;
  assign \DFF_337.D  = \DFF_257.Q ;
  assign \DFF_338.CK  = CK;
  assign \DFF_338.D  = \DFF_337.Q ;
  assign \DFF_339.CK  = CK;
  assign \DFF_339.D  = \DFF_258.Q ;
  assign \DFF_34.CK  = CK;
  assign \DFF_34.D  = g3216;
  assign \DFF_340.CK  = CK;
  assign \DFF_340.D  = \DFF_339.Q ;
  assign \DFF_341.CK  = CK;
  assign \DFF_341.D  = \DFF_259.Q ;
  assign \DFF_342.CK  = CK;
  assign \DFF_342.D  = \DFF_341.Q ;
  assign \DFF_343.CK  = CK;
  assign \DFF_343.D  = \DFF_260.Q ;
  assign \DFF_344.CK  = CK;
  assign \DFF_344.D  = \DFF_343.Q ;
  assign \DFF_345.CK  = CK;
  assign \DFF_345.D  = \DFF_261.Q ;
  assign \DFF_346.CK  = CK;
  assign \DFF_346.D  = \DFF_345.Q ;
  assign \DFF_347.CK  = CK;
  assign \DFF_347.D  = \DFF_262.Q ;
  assign \DFF_348.CK  = CK;
  assign \DFF_348.D  = \DFF_347.Q ;
  assign \DFF_349.CK  = CK;
  assign \DFF_349.D  = \DFF_263.Q ;
  assign \DFF_35.CK  = CK;
  assign \DFF_35.D  = g3215;
  assign \DFF_350.CK  = CK;
  assign \DFF_350.D  = \DFF_349.Q ;
  assign \DFF_351.CK  = CK;
  assign \DFF_351.D  = \DFF_264.Q ;
  assign \DFF_352.CK  = CK;
  assign \DFF_352.D  = \DFF_351.Q ;
  assign \DFF_353.CK  = CK;
  assign \DFF_353.D  = \DFF_1563.Q ;
  assign \DFF_353.Q  = \DFF_1504.Q ;
  assign \DFF_354.CK  = CK;
  assign \DFF_354.D  = \DFF_1504.Q ;
  assign \DFF_354.Q  = \DFF_1505.Q ;
  assign \DFF_355.CK  = CK;
  assign \DFF_355.D  = \DFF_1505.Q ;
  assign \DFF_355.Q  = \DFF_1506.Q ;
  assign \DFF_356.CK  = CK;
  assign \DFF_356.D  = \DFF_1563.Q ;
  assign \DFF_356.Q  = \DFF_1504.Q ;
  assign \DFF_357.CK  = CK;
  assign \DFF_357.D  = \DFF_1504.Q ;
  assign \DFF_357.Q  = \DFF_1505.Q ;
  assign \DFF_358.CK  = CK;
  assign \DFF_358.D  = \DFF_1505.Q ;
  assign \DFF_358.Q  = \DFF_1506.Q ;
  assign \DFF_359.CK  = CK;
  assign \DFF_36.CK  = CK;
  assign \DFF_36.D  = g3214;
  assign \DFF_360.CK  = CK;
  assign \DFF_361.CK  = CK;
  assign \DFF_362.CK  = CK;
  assign \DFF_363.CK  = CK;
  assign \DFF_363.D  = \DFF_362.Q ;
  assign \DFF_364.CK  = CK;
  assign \DFF_364.D  = \DFF_363.Q ;
  assign \DFF_365.CK  = CK;
  assign \DFF_365.D  = \DFF_383.Q ;
  assign \DFF_366.CK  = CK;
  assign \DFF_366.D  = \DFF_365.Q ;
  assign \DFF_367.CK  = CK;
  assign \DFF_367.D  = \DFF_384.Q ;
  assign \DFF_368.CK  = CK;
  assign \DFF_368.D  = \DFF_367.Q ;
  assign \DFF_369.CK  = CK;
  assign \DFF_369.D  = \DFF_385.Q ;
  assign \DFF_37.CK  = CK;
  assign \DFF_37.D  = g3213;
  assign \DFF_370.CK  = CK;
  assign \DFF_370.D  = \DFF_369.Q ;
  assign \DFF_371.CK  = CK;
  assign \DFF_371.D  = \DFF_392.Q ;
  assign \DFF_372.CK  = CK;
  assign \DFF_372.D  = \DFF_371.Q ;
  assign \DFF_373.CK  = CK;
  assign \DFF_373.D  = \DFF_393.Q ;
  assign \DFF_374.CK  = CK;
  assign \DFF_374.D  = \DFF_373.Q ;
  assign \DFF_375.CK  = CK;
  assign \DFF_375.D  = \DFF_394.Q ;
  assign \DFF_376.CK  = CK;
  assign \DFF_376.D  = \DFF_375.Q ;
  assign \DFF_377.CK  = CK;
  assign \DFF_377.D  = \DFF_3.Q ;
  assign \DFF_377.Q  = \DFF_1427.Q ;
  assign \DFF_378.CK  = CK;
  assign \DFF_378.D  = \DFF_1427.Q ;
  assign \DFF_378.Q  = \DFF_1428.Q ;
  assign \DFF_379.CK  = CK;
  assign \DFF_379.D  = \DFF_1428.Q ;
  assign \DFF_379.Q  = \DFF_1429.Q ;
  assign \DFF_38.CK  = CK;
  assign \DFF_380.CK  = CK;
  assign \DFF_381.CK  = CK;
  assign \DFF_382.CK  = CK;
  assign \DFF_383.CK  = CK;
  assign \DFF_384.CK  = CK;
  assign \DFF_385.CK  = CK;
  assign \DFF_386.CK  = CK;
  assign \DFF_387.CK  = CK;
  assign \DFF_388.CK  = CK;
  assign \DFF_389.CK  = CK;
  assign \DFF_39.CK  = CK;
  assign \DFF_390.CK  = CK;
  assign \DFF_391.CK  = CK;
  assign \DFF_392.CK  = CK;
  assign \DFF_393.CK  = CK;
  assign \DFF_394.CK  = CK;
  assign \DFF_395.CK  = CK;
  assign \DFF_396.CK  = CK;
  assign \DFF_396.D  = \DFF_395.Q ;
  assign \DFF_397.CK  = CK;
  assign \DFF_397.D  = \DFF_396.Q ;
  assign \DFF_398.CK  = CK;
  assign \DFF_399.CK  = CK;
  assign \DFF_399.D  = \DFF_398.Q ;
  assign \DFF_4.CK  = CK;
  assign \DFF_40.CK  = CK;
  assign \DFF_400.CK  = CK;
  assign \DFF_401.CK  = CK;
  assign \DFF_402.CK  = CK;
  assign \DFF_402.D  = \DFF_401.Q ;
  assign \DFF_403.CK  = CK;
  assign \DFF_404.CK  = CK;
  assign \DFF_404.D  = \DFF_403.Q ;
  assign \DFF_405.CK  = CK;
  assign \DFF_406.CK  = CK;
  assign \DFF_407.CK  = CK;
  assign \DFF_408.CK  = CK;
  assign \DFF_409.CK  = CK;
  assign \DFF_41.CK  = CK;
  assign \DFF_410.CK  = CK;
  assign \DFF_411.CK  = CK;
  assign \DFF_412.CK  = CK;
  assign \DFF_413.CK  = CK;
  assign \DFF_414.CK  = CK;
  assign \DFF_415.CK  = CK;
  assign \DFF_416.CK  = CK;
  assign \DFF_417.CK  = CK;
  assign \DFF_418.CK  = CK;
  assign \DFF_419.CK  = CK;
  assign \DFF_42.CK  = CK;
  assign \DFF_420.CK  = CK;
  assign \DFF_421.CK  = CK;
  assign \DFF_422.CK  = CK;
  assign \DFF_423.CK  = CK;
  assign \DFF_424.CK  = CK;
  assign \DFF_425.CK  = CK;
  assign \DFF_426.CK  = CK;
  assign \DFF_427.CK  = CK;
  assign \DFF_428.CK  = CK;
  assign \DFF_429.CK  = CK;
  assign \DFF_43.CK  = CK;
  assign \DFF_430.CK  = CK;
  assign \DFF_431.CK  = CK;
  assign \DFF_432.CK  = CK;
  assign \DFF_432.D  = \DFF_402.Q ;
  assign \DFF_433.CK  = CK;
  assign \DFF_434.CK  = CK;
  assign \DFF_435.CK  = CK;
  assign \DFF_436.CK  = CK;
  assign \DFF_437.CK  = CK;
  assign \DFF_438.CK  = CK;
  assign \DFF_439.CK  = CK;
  assign \DFF_44.CK  = CK;
  assign \DFF_440.CK  = CK;
  assign \DFF_441.CK  = CK;
  assign \DFF_442.CK  = CK;
  assign \DFF_443.CK  = CK;
  assign \DFF_443.D  = \DFF_442.Q ;
  assign \DFF_444.CK  = CK;
  assign \DFF_445.CK  = CK;
  assign \DFF_446.CK  = CK;
  assign \DFF_447.CK  = CK;
  assign \DFF_448.CK  = CK;
  assign \DFF_449.CK  = CK;
  assign \DFF_45.CK  = CK;
  assign \DFF_450.CK  = CK;
  assign \DFF_451.CK  = CK;
  assign \DFF_452.CK  = CK;
  assign \DFF_453.CK  = CK;
  assign \DFF_454.CK  = CK;
  assign \DFF_454.D  = \DFF_1563.Q ;
  assign \DFF_454.Q  = \DFF_1504.Q ;
  assign \DFF_455.CK  = CK;
  assign \DFF_455.D  = \DFF_1504.Q ;
  assign \DFF_455.Q  = \DFF_1505.Q ;
  assign \DFF_456.CK  = CK;
  assign \DFF_456.D  = \DFF_1505.Q ;
  assign \DFF_456.Q  = \DFF_1506.Q ;
  assign \DFF_457.CK  = CK;
  assign \DFF_458.CK  = CK;
  assign \DFF_459.CK  = CK;
  assign \DFF_46.CK  = CK;
  assign \DFF_460.CK  = CK;
  assign \DFF_461.CK  = CK;
  assign \DFF_462.CK  = CK;
  assign \DFF_463.CK  = CK;
  assign \DFF_464.CK  = CK;
  assign \DFF_465.CK  = CK;
  assign \DFF_466.CK  = CK;
  assign \DFF_467.CK  = CK;
  assign \DFF_468.CK  = CK;
  assign \DFF_469.CK  = CK;
  assign \DFF_47.CK  = CK;
  assign \DFF_470.CK  = CK;
  assign \DFF_471.CK  = CK;
  assign \DFF_472.CK  = CK;
  assign \DFF_473.CK  = CK;
  assign \DFF_474.CK  = CK;
  assign \DFF_475.CK  = CK;
  assign \DFF_476.CK  = CK;
  assign \DFF_477.CK  = CK;
  assign \DFF_478.CK  = CK;
  assign \DFF_479.CK  = CK;
  assign \DFF_48.CK  = CK;
  assign \DFF_48.D  = \DFF_47.Q ;
  assign \DFF_480.CK  = CK;
  assign \DFF_481.CK  = CK;
  assign \DFF_482.CK  = CK;
  assign \DFF_483.CK  = CK;
  assign \DFF_484.CK  = CK;
  assign \DFF_485.CK  = CK;
  assign \DFF_486.CK  = CK;
  assign \DFF_487.CK  = CK;
  assign \DFF_488.CK  = CK;
  assign \DFF_489.CK  = CK;
  assign \DFF_49.CK  = CK;
  assign \DFF_490.CK  = CK;
  assign \DFF_491.CK  = CK;
  assign \DFF_492.CK  = CK;
  assign \DFF_493.CK  = CK;
  assign \DFF_494.CK  = CK;
  assign \DFF_495.CK  = CK;
  assign \DFF_496.CK  = CK;
  assign \DFF_497.CK  = CK;
  assign \DFF_498.CK  = CK;
  assign \DFF_499.CK  = CK;
  assign \DFF_5.CK  = CK;
  assign \DFF_50.CK  = CK;
  assign \DFF_50.D  = \DFF_49.Q ;
  assign \DFF_500.CK  = CK;
  assign \DFF_501.CK  = CK;
  assign \DFF_502.CK  = CK;
  assign \DFF_503.CK  = CK;
  assign \DFF_504.CK  = CK;
  assign \DFF_505.CK  = CK;
  assign \DFF_506.CK  = CK;
  assign \DFF_507.CK  = CK;
  assign \DFF_508.CK  = CK;
  assign \DFF_509.CK  = CK;
  assign \DFF_51.CK  = CK;
  assign \DFF_510.CK  = CK;
  assign \DFF_511.CK  = CK;
  assign \DFF_511.D  = \DFF_3.Q ;
  assign \DFF_511.Q  = \DFF_1427.Q ;
  assign \DFF_512.CK  = CK;
  assign \DFF_512.D  = \DFF_1427.Q ;
  assign \DFF_512.Q  = \DFF_1428.Q ;
  assign \DFF_513.CK  = CK;
  assign \DFF_513.D  = \DFF_1428.Q ;
  assign \DFF_513.Q  = \DFF_1429.Q ;
  assign \DFF_514.CK  = CK;
  assign \DFF_515.CK  = CK;
  assign \DFF_516.CK  = CK;
  assign \DFF_517.CK  = CK;
  assign \DFF_518.CK  = CK;
  assign \DFF_519.CK  = CK;
  assign \DFF_52.CK  = CK;
  assign \DFF_52.D  = \DFF_51.Q ;
  assign \DFF_520.CK  = CK;
  assign \DFF_521.CK  = CK;
  assign \DFF_522.CK  = CK;
  assign \DFF_523.CK  = CK;
  assign \DFF_524.CK  = CK;
  assign \DFF_525.CK  = CK;
  assign \DFF_526.CK  = CK;
  assign \DFF_527.CK  = CK;
  assign \DFF_528.CK  = CK;
  assign \DFF_529.CK  = CK;
  assign \DFF_53.CK  = CK;
  assign \DFF_530.CK  = CK;
  assign \DFF_531.CK  = CK;
  assign \DFF_532.CK  = CK;
  assign \DFF_533.CK  = CK;
  assign \DFF_534.CK  = CK;
  assign \DFF_535.CK  = CK;
  assign \DFF_536.CK  = CK;
  assign \DFF_537.CK  = CK;
  assign \DFF_538.CK  = CK;
  assign \DFF_539.CK  = CK;
  assign \DFF_54.CK  = CK;
  assign \DFF_54.D  = \DFF_53.Q ;
  assign \DFF_540.CK  = CK;
  assign \DFF_541.CK  = CK;
  assign \DFF_542.CK  = CK;
  assign \DFF_543.CK  = CK;
  assign \DFF_544.CK  = CK;
  assign \DFF_545.CK  = CK;
  assign \DFF_546.CK  = CK;
  assign \DFF_547.CK  = CK;
  assign \DFF_548.CK  = CK;
  assign \DFF_549.CK  = CK;
  assign \DFF_55.CK  = CK;
  assign \DFF_550.CK  = CK;
  assign \DFF_551.CK  = CK;
  assign \DFF_552.CK  = CK;
  assign \DFF_553.CK  = CK;
  assign \DFF_554.CK  = CK;
  assign \DFF_555.CK  = CK;
  assign \DFF_556.CK  = CK;
  assign \DFF_557.CK  = CK;
  assign \DFF_558.CK  = CK;
  assign \DFF_559.CK  = CK;
  assign \DFF_56.CK  = CK;
  assign \DFF_56.D  = \DFF_55.Q ;
  assign \DFF_560.CK  = CK;
  assign \DFF_561.CK  = CK;
  assign \DFF_562.CK  = CK;
  assign \DFF_563.CK  = CK;
  assign \DFF_564.CK  = CK;
  assign \DFF_565.CK  = CK;
  assign \DFF_566.CK  = CK;
  assign \DFF_567.CK  = CK;
  assign \DFF_568.CK  = CK;
  assign \DFF_569.CK  = CK;
  assign \DFF_57.CK  = CK;
  assign \DFF_570.CK  = CK;
  assign \DFF_571.CK  = CK;
  assign \DFF_572.CK  = CK;
  assign \DFF_573.CK  = CK;
  assign \DFF_574.CK  = CK;
  assign \DFF_575.CK  = CK;
  assign \DFF_576.CK  = CK;
  assign \DFF_577.CK  = CK;
  assign \DFF_578.CK  = CK;
  assign \DFF_579.CK  = CK;
  assign \DFF_58.CK  = CK;
  assign \DFF_58.D  = \DFF_57.Q ;
  assign \DFF_580.CK  = CK;
  assign \DFF_581.CK  = CK;
  assign \DFF_582.CK  = CK;
  assign \DFF_583.CK  = CK;
  assign \DFF_584.CK  = CK;
  assign \DFF_585.CK  = CK;
  assign \DFF_586.CK  = CK;
  assign \DFF_587.CK  = CK;
  assign \DFF_588.CK  = CK;
  assign \DFF_589.CK  = CK;
  assign \DFF_59.CK  = CK;
  assign \DFF_590.CK  = CK;
  assign \DFF_591.CK  = CK;
  assign \DFF_592.CK  = CK;
  assign \DFF_593.CK  = CK;
  assign \DFF_594.CK  = CK;
  assign \DFF_595.CK  = CK;
  assign \DFF_596.CK  = CK;
  assign \DFF_596.D  = \DFF_1296.D ;
  assign \DFF_596.Q  = \DFF_1296.Q ;
  assign \DFF_597.CK  = CK;
  assign \DFF_597.D  = \DFF_1296.Q ;
  assign \DFF_597.Q  = \DFF_1297.Q ;
  assign \DFF_598.CK  = CK;
  assign \DFF_598.D  = \DFF_1297.Q ;
  assign \DFF_598.Q  = \DFF_1302.Q ;
  assign \DFF_599.CK  = CK;
  assign \DFF_599.D  = \DFF_3.Q ;
  assign \DFF_599.Q  = \DFF_1427.Q ;
  assign \DFF_6.CK  = CK;
  assign \DFF_60.CK  = CK;
  assign \DFF_60.D  = \DFF_59.Q ;
  assign \DFF_600.CK  = CK;
  assign \DFF_600.D  = \DFF_1427.Q ;
  assign \DFF_600.Q  = \DFF_1428.Q ;
  assign \DFF_601.CK  = CK;
  assign \DFF_601.D  = \DFF_1428.Q ;
  assign \DFF_601.Q  = \DFF_1429.Q ;
  assign \DFF_602.CK  = CK;
  assign \DFF_602.D  = \DFF_1297.Q ;
  assign \DFF_602.Q  = \DFF_1302.Q ;
  assign \DFF_603.CK  = CK;
  assign \DFF_604.CK  = CK;
  assign \DFF_605.CK  = CK;
  assign \DFF_606.CK  = CK;
  assign \DFF_607.CK  = CK;
  assign \DFF_608.CK  = CK;
  assign \DFF_609.CK  = CK;
  assign \DFF_61.CK  = CK;
  assign \DFF_610.CK  = CK;
  assign \DFF_611.CK  = CK;
  assign \DFF_612.CK  = CK;
  assign \DFF_613.CK  = CK;
  assign \DFF_614.CK  = CK;
  assign \DFF_615.CK  = CK;
  assign \DFF_616.CK  = CK;
  assign \DFF_617.CK  = CK;
  assign \DFF_618.CK  = CK;
  assign \DFF_619.CK  = CK;
  assign \DFF_62.CK  = CK;
  assign \DFF_62.D  = \DFF_61.Q ;
  assign \DFF_620.CK  = CK;
  assign \DFF_621.CK  = CK;
  assign \DFF_622.CK  = CK;
  assign \DFF_623.CK  = CK;
  assign \DFF_624.CK  = CK;
  assign \DFF_625.CK  = CK;
  assign \DFF_626.CK  = CK;
  assign \DFF_627.CK  = CK;
  assign \DFF_628.CK  = CK;
  assign \DFF_629.CK  = CK;
  assign \DFF_63.CK  = CK;
  assign \DFF_630.CK  = CK;
  assign \DFF_631.CK  = CK;
  assign \DFF_632.CK  = CK;
  assign \DFF_633.CK  = CK;
  assign \DFF_634.CK  = CK;
  assign \DFF_635.CK  = CK;
  assign \DFF_636.CK  = CK;
  assign \DFF_637.CK  = CK;
  assign \DFF_638.CK  = CK;
  assign \DFF_639.CK  = CK;
  assign \DFF_64.CK  = CK;
  assign \DFF_64.D  = \DFF_63.Q ;
  assign \DFF_640.CK  = CK;
  assign \DFF_641.CK  = CK;
  assign \DFF_642.CK  = CK;
  assign \DFF_643.CK  = CK;
  assign \DFF_644.CK  = CK;
  assign \DFF_645.CK  = CK;
  assign \DFF_646.CK  = CK;
  assign \DFF_647.CK  = CK;
  assign \DFF_648.CK  = CK;
  assign \DFF_649.CK  = CK;
  assign \DFF_649.D  = \DFF_648.Q ;
  assign \DFF_65.CK  = CK;
  assign \DFF_650.CK  = CK;
  assign \DFF_651.CK  = CK;
  assign \DFF_651.D  = \DFF_650.Q ;
  assign \DFF_652.CK  = CK;
  assign \DFF_653.CK  = CK;
  assign \DFF_653.D  = \DFF_652.Q ;
  assign \DFF_654.CK  = CK;
  assign \DFF_655.CK  = CK;
  assign \DFF_655.D  = \DFF_654.Q ;
  assign \DFF_656.CK  = CK;
  assign \DFF_657.CK  = CK;
  assign \DFF_657.D  = \DFF_656.Q ;
  assign \DFF_658.CK  = CK;
  assign \DFF_659.CK  = CK;
  assign \DFF_659.D  = \DFF_658.Q ;
  assign \DFF_66.CK  = CK;
  assign \DFF_66.D  = \DFF_65.Q ;
  assign \DFF_660.CK  = CK;
  assign \DFF_661.CK  = CK;
  assign \DFF_661.D  = \DFF_660.Q ;
  assign \DFF_662.CK  = CK;
  assign \DFF_663.CK  = CK;
  assign \DFF_663.D  = \DFF_662.Q ;
  assign \DFF_664.CK  = CK;
  assign \DFF_664.D  = \DFF_64.Q ;
  assign \DFF_665.CK  = CK;
  assign \DFF_665.D  = \DFF_664.Q ;
  assign \DFF_666.CK  = CK;
  assign \DFF_667.CK  = CK;
  assign \DFF_668.CK  = CK;
  assign \DFF_669.CK  = CK;
  assign \DFF_67.CK  = CK;
  assign \DFF_670.CK  = CK;
  assign \DFF_671.CK  = CK;
  assign \DFF_672.CK  = CK;
  assign \DFF_673.CK  = CK;
  assign \DFF_674.CK  = CK;
  assign \DFF_675.CK  = CK;
  assign \DFF_676.CK  = CK;
  assign \DFF_677.CK  = CK;
  assign \DFF_678.CK  = CK;
  assign \DFF_679.CK  = CK;
  assign \DFF_679.D  = \DFF_603.Q ;
  assign \DFF_68.CK  = CK;
  assign \DFF_68.D  = \DFF_67.Q ;
  assign \DFF_680.CK  = CK;
  assign \DFF_680.D  = \DFF_679.Q ;
  assign \DFF_681.CK  = CK;
  assign \DFF_681.D  = \DFF_604.Q ;
  assign \DFF_682.CK  = CK;
  assign \DFF_682.D  = \DFF_681.Q ;
  assign \DFF_683.CK  = CK;
  assign \DFF_683.D  = \DFF_605.Q ;
  assign \DFF_684.CK  = CK;
  assign \DFF_684.D  = \DFF_683.Q ;
  assign \DFF_685.CK  = CK;
  assign \DFF_685.D  = \DFF_606.Q ;
  assign \DFF_686.CK  = CK;
  assign \DFF_686.D  = \DFF_685.Q ;
  assign \DFF_687.CK  = CK;
  assign \DFF_687.D  = \DFF_607.Q ;
  assign \DFF_688.CK  = CK;
  assign \DFF_688.D  = \DFF_687.Q ;
  assign \DFF_689.CK  = CK;
  assign \DFF_689.D  = \DFF_608.Q ;
  assign \DFF_69.CK  = CK;
  assign \DFF_690.CK  = CK;
  assign \DFF_690.D  = \DFF_689.Q ;
  assign \DFF_691.CK  = CK;
  assign \DFF_691.D  = \DFF_609.Q ;
  assign \DFF_692.CK  = CK;
  assign \DFF_692.D  = \DFF_691.Q ;
  assign \DFF_693.CK  = CK;
  assign \DFF_693.D  = \DFF_610.Q ;
  assign \DFF_694.CK  = CK;
  assign \DFF_694.D  = \DFF_693.Q ;
  assign \DFF_695.CK  = CK;
  assign \DFF_695.D  = \DFF_611.Q ;
  assign \DFF_696.CK  = CK;
  assign \DFF_696.D  = \DFF_695.Q ;
  assign \DFF_697.CK  = CK;
  assign \DFF_697.D  = \DFF_612.Q ;
  assign \DFF_698.CK  = CK;
  assign \DFF_698.D  = \DFF_697.Q ;
  assign \DFF_699.CK  = CK;
  assign \DFF_699.D  = \DFF_613.Q ;
  assign \DFF_7.CK  = CK;
  assign \DFF_70.CK  = CK;
  assign \DFF_70.D  = \DFF_69.Q ;
  assign \DFF_700.CK  = CK;
  assign \DFF_700.D  = \DFF_699.Q ;
  assign \DFF_701.CK  = CK;
  assign \DFF_701.D  = \DFF_614.Q ;
  assign \DFF_702.CK  = CK;
  assign \DFF_702.D  = \DFF_701.Q ;
  assign \DFF_703.CK  = CK;
  assign \DFF_703.D  = \DFF_1563.Q ;
  assign \DFF_703.Q  = \DFF_1504.Q ;
  assign \DFF_704.CK  = CK;
  assign \DFF_704.D  = \DFF_1504.Q ;
  assign \DFF_704.Q  = \DFF_1505.Q ;
  assign \DFF_705.CK  = CK;
  assign \DFF_705.D  = \DFF_1505.Q ;
  assign \DFF_705.Q  = \DFF_1506.Q ;
  assign \DFF_706.CK  = CK;
  assign \DFF_706.D  = \DFF_1563.Q ;
  assign \DFF_706.Q  = \DFF_1504.Q ;
  assign \DFF_707.CK  = CK;
  assign \DFF_707.D  = \DFF_1504.Q ;
  assign \DFF_707.Q  = \DFF_1505.Q ;
  assign \DFF_708.CK  = CK;
  assign \DFF_708.D  = \DFF_1505.Q ;
  assign \DFF_708.Q  = \DFF_1506.Q ;
  assign \DFF_709.CK  = CK;
  assign \DFF_71.CK  = CK;
  assign \DFF_710.CK  = CK;
  assign \DFF_711.CK  = CK;
  assign \DFF_712.CK  = CK;
  assign \DFF_713.CK  = CK;
  assign \DFF_713.D  = \DFF_712.Q ;
  assign \DFF_714.CK  = CK;
  assign \DFF_714.D  = \DFF_713.Q ;
  assign \DFF_715.CK  = CK;
  assign \DFF_715.D  = \DFF_733.Q ;
  assign \DFF_716.CK  = CK;
  assign \DFF_716.D  = \DFF_715.Q ;
  assign \DFF_717.CK  = CK;
  assign \DFF_717.D  = \DFF_734.Q ;
  assign \DFF_718.CK  = CK;
  assign \DFF_718.D  = \DFF_717.Q ;
  assign \DFF_719.CK  = CK;
  assign \DFF_719.D  = \DFF_735.Q ;
  assign \DFF_72.CK  = CK;
  assign \DFF_72.D  = \DFF_71.Q ;
  assign \DFF_720.CK  = CK;
  assign \DFF_720.D  = \DFF_719.Q ;
  assign \DFF_721.CK  = CK;
  assign \DFF_721.D  = \DFF_742.Q ;
  assign \DFF_722.CK  = CK;
  assign \DFF_722.D  = \DFF_721.Q ;
  assign \DFF_723.CK  = CK;
  assign \DFF_723.D  = \DFF_743.Q ;
  assign \DFF_724.CK  = CK;
  assign \DFF_724.D  = \DFF_723.Q ;
  assign \DFF_725.CK  = CK;
  assign \DFF_725.D  = \DFF_744.Q ;
  assign \DFF_726.CK  = CK;
  assign \DFF_726.D  = \DFF_725.Q ;
  assign \DFF_727.CK  = CK;
  assign \DFF_727.D  = \DFF_3.Q ;
  assign \DFF_727.Q  = \DFF_1427.Q ;
  assign \DFF_728.CK  = CK;
  assign \DFF_728.D  = \DFF_1427.Q ;
  assign \DFF_728.Q  = \DFF_1428.Q ;
  assign \DFF_729.CK  = CK;
  assign \DFF_729.D  = \DFF_1428.Q ;
  assign \DFF_729.Q  = \DFF_1429.Q ;
  assign \DFF_73.CK  = CK;
  assign \DFF_730.CK  = CK;
  assign \DFF_731.CK  = CK;
  assign \DFF_732.CK  = CK;
  assign \DFF_733.CK  = CK;
  assign \DFF_734.CK  = CK;
  assign \DFF_735.CK  = CK;
  assign \DFF_736.CK  = CK;
  assign \DFF_737.CK  = CK;
  assign \DFF_738.CK  = CK;
  assign \DFF_739.CK  = CK;
  assign \DFF_74.CK  = CK;
  assign \DFF_74.D  = \DFF_73.Q ;
  assign \DFF_740.CK  = CK;
  assign \DFF_741.CK  = CK;
  assign \DFF_742.CK  = CK;
  assign \DFF_743.CK  = CK;
  assign \DFF_744.CK  = CK;
  assign \DFF_745.CK  = CK;
  assign \DFF_746.CK  = CK;
  assign \DFF_746.D  = \DFF_745.Q ;
  assign \DFF_747.CK  = CK;
  assign \DFF_747.D  = \DFF_746.Q ;
  assign \DFF_748.CK  = CK;
  assign \DFF_749.CK  = CK;
  assign \DFF_749.D  = \DFF_748.Q ;
  assign \DFF_75.CK  = CK;
  assign \DFF_750.CK  = CK;
  assign \DFF_751.CK  = CK;
  assign \DFF_752.CK  = CK;
  assign \DFF_752.D  = \DFF_751.Q ;
  assign \DFF_753.CK  = CK;
  assign \DFF_754.CK  = CK;
  assign \DFF_754.D  = \DFF_753.Q ;
  assign \DFF_755.CK  = CK;
  assign \DFF_756.CK  = CK;
  assign \DFF_757.CK  = CK;
  assign \DFF_758.CK  = CK;
  assign \DFF_759.CK  = CK;
  assign \DFF_76.CK  = CK;
  assign \DFF_76.D  = \DFF_75.Q ;
  assign \DFF_760.CK  = CK;
  assign \DFF_761.CK  = CK;
  assign \DFF_762.CK  = CK;
  assign \DFF_763.CK  = CK;
  assign \DFF_764.CK  = CK;
  assign \DFF_765.CK  = CK;
  assign \DFF_766.CK  = CK;
  assign \DFF_767.CK  = CK;
  assign \DFF_768.CK  = CK;
  assign \DFF_769.CK  = CK;
  assign \DFF_77.CK  = CK;
  assign \DFF_770.CK  = CK;
  assign \DFF_771.CK  = CK;
  assign \DFF_772.CK  = CK;
  assign \DFF_773.CK  = CK;
  assign \DFF_774.CK  = CK;
  assign \DFF_775.CK  = CK;
  assign \DFF_776.CK  = CK;
  assign \DFF_777.CK  = CK;
  assign \DFF_778.CK  = CK;
  assign \DFF_779.CK  = CK;
  assign \DFF_78.CK  = CK;
  assign \DFF_78.D  = \DFF_77.Q ;
  assign \DFF_780.CK  = CK;
  assign \DFF_781.CK  = CK;
  assign \DFF_782.CK  = CK;
  assign \DFF_782.D  = \DFF_752.Q ;
  assign \DFF_783.CK  = CK;
  assign \DFF_784.CK  = CK;
  assign \DFF_785.CK  = CK;
  assign \DFF_786.CK  = CK;
  assign \DFF_787.CK  = CK;
  assign \DFF_788.CK  = CK;
  assign \DFF_789.CK  = CK;
  assign \DFF_79.CK  = CK;
  assign \DFF_790.CK  = CK;
  assign \DFF_791.CK  = CK;
  assign \DFF_792.CK  = CK;
  assign \DFF_793.CK  = CK;
  assign \DFF_793.D  = \DFF_792.Q ;
  assign \DFF_794.CK  = CK;
  assign \DFF_795.CK  = CK;
  assign \DFF_796.CK  = CK;
  assign \DFF_797.CK  = CK;
  assign \DFF_798.CK  = CK;
  assign \DFF_799.CK  = CK;
  assign \DFF_8.CK  = CK;
  assign \DFF_80.CK  = CK;
  assign \DFF_80.D  = \DFF_79.Q ;
  assign \DFF_800.CK  = CK;
  assign \DFF_801.CK  = CK;
  assign \DFF_802.CK  = CK;
  assign \DFF_803.CK  = CK;
  assign \DFF_804.CK  = CK;
  assign \DFF_804.D  = \DFF_1563.Q ;
  assign \DFF_804.Q  = \DFF_1504.Q ;
  assign \DFF_805.CK  = CK;
  assign \DFF_805.D  = \DFF_1504.Q ;
  assign \DFF_805.Q  = \DFF_1505.Q ;
  assign \DFF_806.CK  = CK;
  assign \DFF_806.D  = \DFF_1505.Q ;
  assign \DFF_806.Q  = \DFF_1506.Q ;
  assign \DFF_807.CK  = CK;
  assign \DFF_808.CK  = CK;
  assign \DFF_809.CK  = CK;
  assign \DFF_81.CK  = CK;
  assign \DFF_810.CK  = CK;
  assign \DFF_811.CK  = CK;
  assign \DFF_812.CK  = CK;
  assign \DFF_813.CK  = CK;
  assign \DFF_814.CK  = CK;
  assign \DFF_815.CK  = CK;
  assign \DFF_816.CK  = CK;
  assign \DFF_817.CK  = CK;
  assign \DFF_818.CK  = CK;
  assign \DFF_819.CK  = CK;
  assign \DFF_82.CK  = CK;
  assign \DFF_82.D  = \DFF_81.Q ;
  assign \DFF_820.CK  = CK;
  assign \DFF_821.CK  = CK;
  assign \DFF_822.CK  = CK;
  assign \DFF_823.CK  = CK;
  assign \DFF_824.CK  = CK;
  assign \DFF_825.CK  = CK;
  assign \DFF_826.CK  = CK;
  assign \DFF_827.CK  = CK;
  assign \DFF_828.CK  = CK;
  assign \DFF_829.CK  = CK;
  assign \DFF_83.CK  = CK;
  assign \DFF_830.CK  = CK;
  assign \DFF_831.CK  = CK;
  assign \DFF_832.CK  = CK;
  assign \DFF_833.CK  = CK;
  assign \DFF_834.CK  = CK;
  assign \DFF_835.CK  = CK;
  assign \DFF_836.CK  = CK;
  assign \DFF_837.CK  = CK;
  assign \DFF_838.CK  = CK;
  assign \DFF_839.CK  = CK;
  assign \DFF_84.CK  = CK;
  assign \DFF_840.CK  = CK;
  assign \DFF_841.CK  = CK;
  assign \DFF_842.CK  = CK;
  assign \DFF_843.CK  = CK;
  assign \DFF_844.CK  = CK;
  assign \DFF_845.CK  = CK;
  assign \DFF_846.CK  = CK;
  assign \DFF_847.CK  = CK;
  assign \DFF_848.CK  = CK;
  assign \DFF_849.CK  = CK;
  assign \DFF_85.CK  = CK;
  assign \DFF_850.CK  = CK;
  assign \DFF_851.CK  = CK;
  assign \DFF_852.CK  = CK;
  assign \DFF_853.CK  = CK;
  assign \DFF_854.CK  = CK;
  assign \DFF_855.CK  = CK;
  assign \DFF_856.CK  = CK;
  assign \DFF_857.CK  = CK;
  assign \DFF_858.CK  = CK;
  assign \DFF_859.CK  = CK;
  assign \DFF_86.CK  = CK;
  assign \DFF_860.CK  = CK;
  assign \DFF_861.CK  = CK;
  assign \DFF_861.D  = \DFF_3.Q ;
  assign \DFF_861.Q  = \DFF_1427.Q ;
  assign \DFF_862.CK  = CK;
  assign \DFF_862.D  = \DFF_1427.Q ;
  assign \DFF_862.Q  = \DFF_1428.Q ;
  assign \DFF_863.CK  = CK;
  assign \DFF_863.D  = \DFF_1428.Q ;
  assign \DFF_863.Q  = \DFF_1429.Q ;
  assign \DFF_864.CK  = CK;
  assign \DFF_865.CK  = CK;
  assign \DFF_866.CK  = CK;
  assign \DFF_867.CK  = CK;
  assign \DFF_868.CK  = CK;
  assign \DFF_869.CK  = CK;
  assign \DFF_87.CK  = CK;
  assign \DFF_870.CK  = CK;
  assign \DFF_871.CK  = CK;
  assign \DFF_872.CK  = CK;
  assign \DFF_873.CK  = CK;
  assign \DFF_874.CK  = CK;
  assign \DFF_875.CK  = CK;
  assign \DFF_876.CK  = CK;
  assign \DFF_877.CK  = CK;
  assign \DFF_878.CK  = CK;
  assign \DFF_879.CK  = CK;
  assign \DFF_88.CK  = CK;
  assign \DFF_880.CK  = CK;
  assign \DFF_881.CK  = CK;
  assign \DFF_882.CK  = CK;
  assign \DFF_883.CK  = CK;
  assign \DFF_884.CK  = CK;
  assign \DFF_885.CK  = CK;
  assign \DFF_886.CK  = CK;
  assign \DFF_887.CK  = CK;
  assign \DFF_888.CK  = CK;
  assign \DFF_889.CK  = CK;
  assign \DFF_89.CK  = CK;
  assign \DFF_890.CK  = CK;
  assign \DFF_891.CK  = CK;
  assign \DFF_892.CK  = CK;
  assign \DFF_893.CK  = CK;
  assign \DFF_894.CK  = CK;
  assign \DFF_895.CK  = CK;
  assign \DFF_896.CK  = CK;
  assign \DFF_897.CK  = CK;
  assign \DFF_898.CK  = CK;
  assign \DFF_899.CK  = CK;
  assign \DFF_9.CK  = CK;
  assign \DFF_90.CK  = CK;
  assign \DFF_900.CK  = CK;
  assign \DFF_901.CK  = CK;
  assign \DFF_902.CK  = CK;
  assign \DFF_903.CK  = CK;
  assign \DFF_904.CK  = CK;
  assign \DFF_905.CK  = CK;
  assign \DFF_906.CK  = CK;
  assign \DFF_907.CK  = CK;
  assign \DFF_908.CK  = CK;
  assign \DFF_909.CK  = CK;
  assign \DFF_91.CK  = CK;
  assign \DFF_910.CK  = CK;
  assign \DFF_911.CK  = CK;
  assign \DFF_912.CK  = CK;
  assign \DFF_913.CK  = CK;
  assign \DFF_914.CK  = CK;
  assign \DFF_915.CK  = CK;
  assign \DFF_916.CK  = CK;
  assign \DFF_917.CK  = CK;
  assign \DFF_918.CK  = CK;
  assign \DFF_919.CK  = CK;
  assign \DFF_92.CK  = CK;
  assign \DFF_92.D  = \DFF_1563.Q ;
  assign \DFF_92.Q  = \DFF_1504.Q ;
  assign \DFF_920.CK  = CK;
  assign \DFF_921.CK  = CK;
  assign \DFF_922.CK  = CK;
  assign \DFF_923.CK  = CK;
  assign \DFF_924.CK  = CK;
  assign \DFF_925.CK  = CK;
  assign \DFF_926.CK  = CK;
  assign \DFF_927.CK  = CK;
  assign \DFF_928.CK  = CK;
  assign \DFF_929.CK  = CK;
  assign \DFF_93.CK  = CK;
  assign \DFF_93.D  = \DFF_1504.Q ;
  assign \DFF_93.Q  = \DFF_1505.Q ;
  assign \DFF_930.CK  = CK;
  assign \DFF_931.CK  = CK;
  assign \DFF_932.CK  = CK;
  assign \DFF_933.CK  = CK;
  assign \DFF_934.CK  = CK;
  assign \DFF_935.CK  = CK;
  assign \DFF_936.CK  = CK;
  assign \DFF_937.CK  = CK;
  assign \DFF_938.CK  = CK;
  assign \DFF_939.CK  = CK;
  assign \DFF_94.CK  = CK;
  assign \DFF_94.D  = \DFF_1505.Q ;
  assign \DFF_94.Q  = \DFF_1506.Q ;
  assign \DFF_940.CK  = CK;
  assign \DFF_941.CK  = CK;
  assign \DFF_942.CK  = CK;
  assign \DFF_943.CK  = CK;
  assign \DFF_944.CK  = CK;
  assign \DFF_945.CK  = CK;
  assign \DFF_946.CK  = CK;
  assign \DFF_946.D  = \DFF_1296.D ;
  assign \DFF_946.Q  = \DFF_1296.Q ;
  assign \DFF_947.CK  = CK;
  assign \DFF_947.D  = \DFF_1296.Q ;
  assign \DFF_947.Q  = \DFF_1297.Q ;
  assign \DFF_948.CK  = CK;
  assign \DFF_948.D  = \DFF_1297.Q ;
  assign \DFF_948.Q  = \DFF_1302.Q ;
  assign \DFF_949.CK  = CK;
  assign \DFF_949.D  = \DFF_3.Q ;
  assign \DFF_949.Q  = \DFF_1427.Q ;
  assign \DFF_95.CK  = CK;
  assign \DFF_950.CK  = CK;
  assign \DFF_950.D  = \DFF_1427.Q ;
  assign \DFF_950.Q  = \DFF_1428.Q ;
  assign \DFF_951.CK  = CK;
  assign \DFF_951.D  = \DFF_1428.Q ;
  assign \DFF_951.Q  = \DFF_1429.Q ;
  assign \DFF_952.CK  = CK;
  assign \DFF_952.D  = \DFF_1297.Q ;
  assign \DFF_952.Q  = \DFF_1302.Q ;
  assign \DFF_953.CK  = CK;
  assign \DFF_954.CK  = CK;
  assign \DFF_955.CK  = CK;
  assign \DFF_956.CK  = CK;
  assign \DFF_957.CK  = CK;
  assign \DFF_958.CK  = CK;
  assign \DFF_959.CK  = CK;
  assign \DFF_96.CK  = CK;
  assign \DFF_960.CK  = CK;
  assign \DFF_961.CK  = CK;
  assign \DFF_962.CK  = CK;
  assign \DFF_963.CK  = CK;
  assign \DFF_964.CK  = CK;
  assign \DFF_965.CK  = CK;
  assign \DFF_966.CK  = CK;
  assign \DFF_967.CK  = CK;
  assign \DFF_968.CK  = CK;
  assign \DFF_969.CK  = CK;
  assign \DFF_97.CK  = CK;
  assign \DFF_970.CK  = CK;
  assign \DFF_971.CK  = CK;
  assign \DFF_972.CK  = CK;
  assign \DFF_973.CK  = CK;
  assign \DFF_974.CK  = CK;
  assign \DFF_975.CK  = CK;
  assign \DFF_976.CK  = CK;
  assign \DFF_977.CK  = CK;
  assign \DFF_978.CK  = CK;
  assign \DFF_979.CK  = CK;
  assign \DFF_98.CK  = CK;
  assign \DFF_980.CK  = CK;
  assign \DFF_981.CK  = CK;
  assign \DFF_982.CK  = CK;
  assign \DFF_983.CK  = CK;
  assign \DFF_984.CK  = CK;
  assign \DFF_985.CK  = CK;
  assign \DFF_986.CK  = CK;
  assign \DFF_987.CK  = CK;
  assign \DFF_988.CK  = CK;
  assign \DFF_989.CK  = CK;
  assign \DFF_99.CK  = CK;
  assign \DFF_990.CK  = CK;
  assign \DFF_991.CK  = CK;
  assign \DFF_992.CK  = CK;
  assign \DFF_993.CK  = CK;
  assign \DFF_994.CK  = CK;
  assign \DFF_995.CK  = CK;
  assign \DFF_996.CK  = CK;
  assign \DFF_997.CK  = CK;
  assign \DFF_998.CK  = CK;
  assign \DFF_999.CK  = CK;
  assign \DFF_999.D  = \DFF_998.Q ;
  assign II13430 = \DFF_310.D ;
  assign II13433 = \DFF_308.D ;
  assign II13501 = \DFF_660.D ;
  assign II13504 = \DFF_658.D ;
  assign II13575 = \DFF_1010.D ;
  assign II13578 = \DFF_1008.D ;
  assign II13601 = \DFF_300.D ;
  assign II13604 = \DFF_298.D ;
  assign II13652 = \DFF_1360.D ;
  assign II13655 = \DFF_1358.D ;
  assign II13677 = \DFF_650.D ;
  assign II13680 = \DFF_648.D ;
  assign II13742 = \DFF_1000.D ;
  assign II13745 = \DFF_998.D ;
  assign II13775 = \DFF_306.D ;
  assign II13801 = \DFF_1350.D ;
  assign II13804 = \DFF_1348.D ;
  assign II13820 = \DFF_656.D ;
  assign II13849 = \DFF_1006.D ;
  assign II13868 = \DFF_1356.D ;
  assign II14163 = \DFF_304.D ;
  assign II14219 = \DFF_654.D ;
  assign II14280 = \DFF_1004.D ;
  assign II14306 = \DFF_312.D ;
  assign II14338 = \DFF_1354.D ;
  assign II14357 = \DFF_662.D ;
  assign II14402 = \DFF_1012.D ;
  assign II14424 = \DFF_302.D ;
  assign II14442 = \DFF_1362.D ;
  assign II14459 = \DFF_652.D ;
  assign II14489 = \DFF_1002.D ;
  assign II14513 = \DFF_1352.D ;
  assign II15562 = \DFF_1016.Q ;
  assign II15580 = \DFF_1366.Q ;
  assign II15629 = \DFF_1366.Q ;
  assign II15850 = \DFF_66.Q ;
  assign II15873 = \DFF_48.Q ;
  assign II15887 = \DFF_38.Q ;
  assign II15899 = \DFF_68.Q ;
  assign II15909 = \DFF_83.Q ;
  assign II15922 = \DFF_50.Q ;
  assign II15932 = \DFF_19.Q ;
  assign II15946 = \DFF_39.Q ;
  assign II15964 = \DFF_70.Q ;
  assign II15975 = \DFF_84.Q ;
  assign II15995 = \DFF_52.Q ;
  assign II16024 = \DFF_40.Q ;
  assign II16056 = \DFF_85.Q ;
  assign II17632 = \DFF_315.Q ;
  assign II17637 = \DFF_313.Q ;
  assign II17641 = \DFF_665.Q ;
  assign II17645 = \DFF_311.Q ;
  assign II17649 = \DFF_663.Q ;
  assign II17653 = \DFF_1015.Q ;
  assign II17658 = \DFF_309.Q ;
  assign II17662 = \DFF_661.Q ;
  assign II17666 = \DFF_1013.Q ;
  assign II17670 = \DFF_1365.Q ;
  assign II17677 = \DFF_307.Q ;
  assign II17681 = \DFF_659.Q ;
  assign II17685 = \DFF_1011.Q ;
  assign II17689 = \DFF_1363.Q ;
  assign II17698 = \DFF_305.Q ;
  assign II17701 = \DFF_657.Q ;
  assign II17705 = \DFF_1009.Q ;
  assign II17709 = \DFF_1361.Q ;
  assign II17721 = \DFF_72.Q ;
  assign II17724 = \DFF_303.Q ;
  assign II17727 = \DFF_655.Q ;
  assign II17730 = \DFF_1007.Q ;
  assign II17734 = \DFF_1359.Q ;
  assign II17750 = \DFF_301.Q ;
  assign II17753 = \DFF_54.Q ;
  assign II17756 = \DFF_653.Q ;
  assign II17759 = \DFF_1005.Q ;
  assign II17762 = \DFF_1357.Q ;
  assign II17780 = \DFF_299.Q ;
  assign II17783 = \DFF_651.Q ;
  assign II17786 = \DFF_41.Q ;
  assign II17789 = \DFF_1003.Q ;
  assign II17792 = \DFF_1355.Q ;
  assign II17813 = \DFF_74.Q ;
  assign II17816 = \DFF_80.Q ;
  assign II17822 = \DFF_649.Q ;
  assign II17825 = \DFF_1001.Q ;
  assign II17828 = \DFF_86.Q ;
  assign II17831 = \DFF_1353.Q ;
  assign II17849 = \DFF_160.Q ;
  assign II17860 = \DFF_56.Q ;
  assign II17863 = \DFF_62.Q ;
  assign II17869 = \DFF_999.Q ;
  assign II17872 = \DFF_1351.Q ;
  assign II17907 = \DFF_42.Q ;
  assign II17910 = \DFF_45.Q ;
  assign II17916 = \DFF_1349.Q ;
  assign II17942 = \DFF_76.Q ;
  assign II17945 = \DFF_316.Q ;
  assign II17969 = \DFF_87.Q ;
  assign II17972 = \DFF_90.Q ;
  assign II17998 = \DFF_316.Q ;
  assign II18013 = \DFF_58.Q ;
  assign II18016 = \DFF_666.Q ;
  assign II18055 = \DFF_316.Q ;
  assign II18070 = \DFF_666.Q ;
  assign II18085 = \DFF_43.Q ;
  assign II18088 = \DFF_1016.Q ;
  assign II18130 = \DFF_78.Q ;
  assign II18136 = \DFF_316.Q ;
  assign II18151 = \DFF_666.Q ;
  assign II18166 = \DFF_1016.Q ;
  assign II18181 = \DFF_88.Q ;
  assign II18184 = \DFF_1366.Q ;
  assign II18226 = \DFF_316.Q ;
  assign II18238 = \DFF_60.Q ;
  assign II18244 = \DFF_666.Q ;
  assign II18259 = \DFF_1016.Q ;
  assign II18274 = \DFF_1366.Q ;
  assign II18311 = \DFF_316.Q ;
  assign II18329 = \DFF_666.Q ;
  assign II18341 = \DFF_44.Q ;
  assign II18347 = \DFF_1016.Q ;
  assign II18362 = \DFF_1366.Q ;
  assign II18405 = \DFF_666.Q ;
  assign II18423 = \DFF_1016.Q ;
  assign II18435 = \DFF_89.Q ;
  assign II18441 = \DFF_1366.Q ;
  assign II18449 = \DFF_72.Q ;
  assign II18452 = \DFF_74.Q ;
  assign II18455 = \DFF_76.Q ;
  assign II18458 = \DFF_78.Q ;
  assign II18461 = \DFF_80.Q ;
  assign II18503 = \DFF_66.Q ;
  assign II18506 = \DFF_68.Q ;
  assign II18509 = \DFF_70.Q ;
  assign II18530 = \DFF_54.Q ;
  assign II18533 = \DFF_56.Q ;
  assign II18536 = \DFF_58.Q ;
  assign II18539 = \DFF_60.Q ;
  assign II18542 = \DFF_62.Q ;
  assign II18584 = \DFF_48.Q ;
  assign II18587 = \DFF_50.Q ;
  assign II18590 = \DFF_52.Q ;
  assign II18611 = \DFF_41.Q ;
  assign II18614 = \DFF_42.Q ;
  assign II18617 = \DFF_43.Q ;
  assign II18620 = \DFF_44.Q ;
  assign II18623 = \DFF_45.Q ;
  assign II18665 = \DFF_38.Q ;
  assign II18668 = \DFF_39.Q ;
  assign II18671 = \DFF_40.Q ;
  assign II18692 = \DFF_86.Q ;
  assign II18695 = \DFF_87.Q ;
  assign II18698 = \DFF_88.Q ;
  assign II18701 = \DFF_89.Q ;
  assign II18704 = \DFF_90.Q ;
  assign II18746 = \DFF_83.Q ;
  assign II18749 = \DFF_84.Q ;
  assign II18752 = \DFF_85.Q ;
  assign II18773 = \DFF_307.Q ;
  assign II18780 = \DFF_655.Q ;
  assign II18787 = \DFF_1003.Q ;
  assign II18794 = \DFF_1351.Q ;
  assign II18810 = \DFF_309.Q ;
  assign II18813 = \DFF_657.Q ;
  assign II18820 = \DFF_1005.Q ;
  assign II18827 = \DFF_1353.Q ;
  assign II18835 = \DFF_659.Q ;
  assign II18838 = \DFF_1007.Q ;
  assign II18845 = \DFF_1355.Q ;
  assign II18854 = \DFF_1009.Q ;
  assign II18857 = \DFF_1357.Q ;
  assign II18866 = \DFF_1359.Q ;
  assign II18969 = \DFF_19.Q ;
  assign II19030 = \DFF_19.Q ;
  assign II19105 = \DFF_19.Q ;
  assign II19195 = \DFF_19.Q ;
  assign II19307 = \DFF_19.Q ;
  assign II19718 = \DFF_19.Q ;
  assign II19727 = \DFF_19.Q ;
  assign II19733 = \DFF_19.Q ;
  assign II19747 = \DFF_19.Q ;
  assign II19750 = \DFF_19.Q ;
  assign II19767 = \DFF_19.Q ;
  assign II19784 = \DFF_19.Q ;
  assign II19787 = \DFF_19.Q ;
  assign II19808 = \DFF_19.Q ;
  assign II19833 = \DFF_19.Q ;
  assign II19836 = \DFF_19.Q ;
  assign II19869 = \DFF_19.Q ;
  assign II19905 = \DFF_19.Q ;
  assign II20299 = \DFF_311.Q ;
  assign II20320 = \DFF_313.Q ;
  assign II20328 = \DFF_661.Q ;
  assign II20347 = \DFF_315.Q ;
  assign II20351 = \DFF_663.Q ;
  assign II20359 = \DFF_1011.Q ;
  assign II20382 = \DFF_299.Q ;
  assign II20386 = \DFF_665.Q ;
  assign II20390 = \DFF_1013.Q ;
  assign II20398 = \DFF_1361.Q ;
  assign II20410 = \DFF_301.Q ;
  assign II20417 = \DFF_649.Q ;
  assign II20421 = \DFF_1015.Q ;
  assign II20425 = \DFF_1363.Q ;
  assign II20444 = \DFF_303.Q ;
  assign II20451 = \DFF_651.Q ;
  assign II20458 = \DFF_999.Q ;
  assign II20462 = \DFF_1365.Q ;
  assign II20479 = \DFF_305.Q ;
  assign II20486 = \DFF_653.Q ;
  assign II20493 = \DFF_1001.Q ;
  assign II20500 = \DFF_1349.Q ;
  assign II20529 = \DFF_299.Q ;
  assign II20532 = \DFF_301.Q ;
  assign II20535 = \DFF_303.Q ;
  assign II20538 = \DFF_305.Q ;
  assign II20541 = \DFF_307.Q ;
  assign II20544 = \DFF_309.Q ;
  assign II20547 = \DFF_311.Q ;
  assign II20550 = \DFF_313.Q ;
  assign II20553 = \DFF_315.Q ;
  assign II20577 = \DFF_649.Q ;
  assign II20580 = \DFF_651.Q ;
  assign II20583 = \DFF_653.Q ;
  assign II20586 = \DFF_655.Q ;
  assign II20589 = \DFF_657.Q ;
  assign II20592 = \DFF_659.Q ;
  assign II20595 = \DFF_661.Q ;
  assign II20598 = \DFF_663.Q ;
  assign II20601 = \DFF_665.Q ;
  assign II20625 = \DFF_999.Q ;
  assign II20628 = \DFF_1001.Q ;
  assign II20631 = \DFF_1003.Q ;
  assign II20634 = \DFF_1005.Q ;
  assign II20637 = \DFF_1007.Q ;
  assign II20640 = \DFF_1009.Q ;
  assign II20643 = \DFF_1011.Q ;
  assign II20646 = \DFF_1013.Q ;
  assign II20649 = \DFF_1015.Q ;
  assign II20673 = \DFF_1349.Q ;
  assign II20676 = \DFF_1351.Q ;
  assign II20679 = \DFF_1353.Q ;
  assign II20682 = \DFF_1355.Q ;
  assign II20685 = \DFF_1357.Q ;
  assign II20688 = \DFF_1359.Q ;
  assign II20691 = \DFF_1361.Q ;
  assign II20694 = \DFF_1363.Q ;
  assign II20697 = \DFF_1365.Q ;
  assign II21381 = \DFF_157.Q ;
  assign II21420 = \DFF_157.Q ;
  assign II24913 = g3234;
  assign II25258 = g3229;
  assign II25308 = g3229;
  assign II25315 = g3229;
  assign II25320 = g3229;
  assign II25325 = g3229;
  assign II26960 = g3229;
  assign II26972 = g3229;
  assign II26985 = g3229;
  assign II32248 = \DFF_146.D ;
  assign II32251 = \DFF_146.D ;
  assign II33257 = \DFF_144.D ;
  assign II33260 = \DFF_144.D ;
  assign II34029 = \DFF_141.D ;
  assign II34032 = \DFF_141.D ;
  assign II35373 = \DFF_146.D ;
  assign II35708 = \DFF_160.D ;
  assign II35711 = \DFF_160.D ;
  assign II35723 = \DFF_146.D ;
  assign II36046 = \DFF_144.D ;
  assign II36162 = \DFF_146.D ;
  assign II36224 = \DFF_131.D ;
  assign II36234 = \DFF_144.D ;
  assign II36362 = \DFF_144.D ;
  assign II36864 = \DFF_141.D ;
  assign II37182 = \DFF_144.D ;
  assign II37188 = \DFF_131.D ;
  assign II37200 = \DFF_144.D ;
  assign II37232 = \DFF_141.D ;
  assign II37252 = \DFF_141.D ;
  assign II37266 = \DFF_141.D ;
  assign II37319 = \DFF_151.D ;
  assign II37400 = \DFF_141.D ;
  assign II37629 = \DFF_141.D ;
  assign II37635 = \DFF_151.D ;
  assign II37647 = \DFF_141.D ;
  assign II37653 = \DFF_141.D ;
  assign II37662 = \DFF_141.D ;
  assign II37793 = \DFF_159.D ;
  assign II38128 = \DFF_160.D ;
  assign II38241 = \DFF_159.D ;
  assign II38330 = \DFF_160.D ;
  assign II38339 = \DFF_160.D ;
  assign II38462 = \DFF_160.D ;
  assign II38764 = \DFF_160.D ;
  assign II38767 = \DFF_160.D ;
  assign II38770 = \DFF_160.D ;
  assign II38801 = \DFF_157.D ;
  assign II38807 = \DFF_157.D ;
  assign II39086 = \DFF_157.D ;
  assign II39089 = \DFF_157.D ;
  assign g1 = \DFF_1635.Q ;
  assign g1000 = \DFF_634.Q ;
  assign g10004 = \DFF_1613.Q ;
  assign g1001 = \DFF_635.Q ;
  assign g10015 = \DFF_82.Q ;
  assign g10016 = \DFF_3.Q ;
  assign g10017 = \DFF_392.Q ;
  assign g10018 = \DFF_1506.Q ;
  assign g1002 = \DFF_636.Q ;
  assign g10021 = \DFF_1505.Q ;
  assign g1003 = \DFF_637.Q ;
  assign g1004 = \DFF_638.Q ;
  assign g10049 = \DFF_1505.Q ;
  assign g1005 = \DFF_639.Q ;
  assign g10052 = \DFF_1504.Q ;
  assign g1006 = \DFF_640.Q ;
  assign g10067 = \DFF_1506.Q ;
  assign g1007 = \DFF_641.Q ;
  assign g10070 = \DFF_1504.Q ;
  assign g1008 = \DFF_644.Q ;
  assign g10086 = \DFF_1435.Q ;
  assign g10087 = \DFF_1506.Q ;
  assign g1009 = \DFF_642.Q ;
  assign g10090 = \DFF_1505.Q ;
  assign g10096 = \DFF_1613.Q ;
  assign g10099 = \DFF_106.Q ;
  assign g101 = \DFF_78.Q ;
  assign g1010 = \DFF_643.Q ;
  assign g10109 = \DFF_1506.Q ;
  assign g1011 = \DFF_702.Q ;
  assign g1012 = \DFF_1504.Q ;
  assign g10124 = \DFF_64.Q ;
  assign g10125 = \DFF_3.Q ;
  assign g10126 = \DFF_742.Q ;
  assign g10127 = \DFF_1506.Q ;
  assign g10130 = \DFF_1505.Q ;
  assign g10158 = \DFF_1505.Q ;
  assign g10161 = \DFF_1504.Q ;
  assign g10176 = \DFF_1506.Q ;
  assign g10179 = \DFF_1504.Q ;
  assign g1018 = \DFF_1505.Q ;
  assign g10189 = \DFF_1613.Q ;
  assign g10214 = \DFF_1506.Q ;
  assign g10229 = \DFF_46.Q ;
  assign g10230 = \DFF_3.Q ;
  assign g10231 = \DFF_1092.Q ;
  assign g10232 = \DFF_1506.Q ;
  assign g10235 = \DFF_1505.Q ;
  assign g1024 = \DFF_1506.Q ;
  assign g10263 = \DFF_1505.Q ;
  assign g10266 = \DFF_1504.Q ;
  assign g10273 = \DFF_1613.Q ;
  assign g10276 = \DFF_1613.Q ;
  assign g1029 = \DFF_679.Q ;
  assign g1030 = \DFF_604.Q ;
  assign g10316 = \DFF_1506.Q ;
  assign g1033 = \DFF_605.Q ;
  assign g10331 = \DFF_91.Q ;
  assign g10332 = \DFF_3.Q ;
  assign g10333 = \DFF_1442.Q ;
  assign g10334 = \DFF_1506.Q ;
  assign g10337 = \DFF_1505.Q ;
  assign g10357 = \DFF_1613.Q ;
  assign g1036 = \DFF_680.Q ;
  assign g1037 = \DFF_681.Q ;
  assign g1038 = \DFF_682.Q ;
  assign g1039 = \DFF_683.Q ;
  assign g1040 = \DFF_684.Q ;
  assign g10409 = \DFF_1506.Q ;
  assign g1041 = \DFF_603.Q ;
  assign g10416 = \DFF_1613.Q ;
  assign g10419 = \DFF_1613.Q ;
  assign g10424 = \DFF_1427.Q ;
  assign g1044 = \DFF_685.Q ;
  assign g1045 = \DFF_607.Q ;
  assign g1048 = \DFF_608.Q ;
  assign g10481 = \DFF_1613.Q ;
  assign g10482 = \DFF_1613.Q ;
  assign g10486 = \DFF_1428.Q ;
  assign g105 = \DFF_76.Q ;
  assign g10500 = \DFF_1427.Q ;
  assign g1051 = \DFF_686.Q ;
  assign g1052 = \DFF_687.Q ;
  assign g1053 = \DFF_688.Q ;
  assign g1054 = \DFF_689.Q ;
  assign g10542 = \DFF_1613.Q ;
  assign g10545 = \DFF_1613.Q ;
  assign g10549 = \DFF_1429.Q ;
  assign g1055 = \DFF_690.Q ;
  assign g1056 = \DFF_606.Q ;
  assign g10560 = \DFF_1428.Q ;
  assign g10574 = \DFF_1427.Q ;
  assign g1059 = \DFF_691.Q ;
  assign g1060 = \DFF_610.Q ;
  assign g10601 = \DFF_1613.Q ;
  assign g10606 = \DFF_1429.Q ;
  assign g10617 = \DFF_1428.Q ;
  assign g1063 = \DFF_611.Q ;
  assign g10631 = \DFF_1427.Q ;
  assign g10646 = \DFF_1613.Q ;
  assign g10653 = \DFF_1429.Q ;
  assign g1066 = \DFF_692.Q ;
  assign g10664 = \DFF_1428.Q ;
  assign g1067 = \DFF_693.Q ;
  assign g1068 = \DFF_694.Q ;
  assign g10683 = \DFF_1429.Q ;
  assign g1069 = \DFF_695.Q ;
  assign g10694 = \DFF_1302.Q ;
  assign g1070 = \DFF_696.Q ;
  assign g1071 = \DFF_609.Q ;
  assign g10714 = \DFF_1302.Q ;
  assign g10730 = \DFF_360.Q ;
  assign g10735 = \DFF_1302.Q ;
  assign g1074 = \DFF_697.Q ;
  assign g10749 = \DFF_710.Q ;
  assign g1075 = \DFF_613.Q ;
  assign g10754 = \DFF_1302.Q ;
  assign g10766 = \DFF_404.Q ;
  assign g10767 = \DFF_1060.Q ;
  assign g10772 = \DFF_754.Q ;
  assign g10773 = \DFF_1410.Q ;
  assign g1078 = \DFF_614.Q ;
  assign g10783 = \DFF_1104.Q ;
  assign g10787 = \DFF_453.D ;
  assign g10788 = \DFF_1454.Q ;
  assign g10792 = \DFF_451.D ;
  assign g10796 = \DFF_803.D ;
  assign g10800 = \DFF_450.D ;
  assign g10804 = \DFF_801.D ;
  assign g10808 = \DFF_1153.D ;
  assign g1081 = \DFF_698.Q ;
  assign g10813 = \DFF_449.D ;
  assign g10817 = \DFF_800.D ;
  assign g1082 = \DFF_699.Q ;
  assign g10821 = \DFF_1151.D ;
  assign g10825 = \DFF_1503.D ;
  assign g10826 = \DFF_1504.Q ;
  assign g1083 = \DFF_700.Q ;
  assign g10830 = \DFF_448.D ;
  assign g10834 = \DFF_799.D ;
  assign g10838 = \DFF_1150.D ;
  assign g1084 = \DFF_701.Q ;
  assign g10842 = \DFF_1501.D ;
  assign g10843 = \DFF_1504.Q ;
  assign g10849 = \DFF_447.D ;
  assign g1085 = \DFF_612.Q ;
  assign g10850 = \DFF_798.D ;
  assign g10854 = \DFF_1149.D ;
  assign g10858 = \DFF_1500.D ;
  assign g10859 = \DFF_1505.Q ;
  assign g10862 = \DFF_1504.Q ;
  assign g10868 = \DFF_304.D ;
  assign g10869 = \DFF_446.D ;
  assign g10870 = \DFF_797.D ;
  assign g10871 = \DFF_1148.D ;
  assign g10875 = \DFF_1499.D ;
  assign g10876 = \DFF_1563.Q ;
  assign g10877 = \DFF_1505.Q ;
  assign g1088 = \DFF_1429.Q ;
  assign g10880 = \DFF_1504.Q ;
  assign g10883 = \DFF_1504.Q ;
  assign g10887 = \DFF_445.D ;
  assign g10888 = \DFF_654.D ;
  assign g10889 = \DFF_796.D ;
  assign g1089 = \DFF_647.Q ;
  assign g10890 = \DFF_1147.D ;
  assign g10891 = \DFF_1498.D ;
  assign g10892 = \DFF_1506.Q ;
  assign g10895 = \DFF_1505.Q ;
  assign g10898 = \DFF_1504.Q ;
  assign g109 = \DFF_74.Q ;
  assign g1090 = \DFF_645.Q ;
  assign g10901 = \DFF_1504.Q ;
  assign g10907 = \DFF_444.D ;
  assign g10908 = \DFF_795.D ;
  assign g10909 = \DFF_1004.D ;
  assign g1091 = \DFF_646.Q ;
  assign g10910 = \DFF_1146.D ;
  assign g10911 = \DFF_1497.D ;
  assign g10912 = \DFF_1506.Q ;
  assign g10915 = \DFF_1505.Q ;
  assign g10918 = \DFF_1504.Q ;
  assign g1092 = \DFF_1428.Q ;
  assign g10921 = \DFF_1505.Q ;
  assign g10924 = \DFF_1504.Q ;
  assign g10930 = \DFF_306.D ;
  assign g10931 = \DFF_312.D ;
  assign g10932 = \DFF_1428.Q ;
  assign g10933 = \DFF_794.D ;
  assign g10934 = \DFF_1145.D ;
  assign g10935 = \DFF_1354.D ;
  assign g10936 = \DFF_1496.D ;
  assign g10937 = \DFF_1506.Q ;
  assign g10940 = \DFF_1505.Q ;
  assign g10943 = \DFF_1504.Q ;
  assign g10946 = \DFF_1505.Q ;
  assign g10949 = \DFF_1504.Q ;
  assign g1095 = \DFF_615.Q ;
  assign g10963 = \DFF_1427.Q ;
  assign g10966 = \DFF_1428.Q ;
  assign g10967 = \DFF_656.D ;
  assign g10968 = \DFF_662.D ;
  assign g10969 = \DFF_1428.Q ;
  assign g10972 = \DFF_1144.D ;
  assign g10973 = \DFF_1495.D ;
  assign g10974 = \DFF_1506.Q ;
  assign g10977 = \DFF_1505.Q ;
  assign g1098 = \DFF_616.Q ;
  assign g10980 = \DFF_1506.Q ;
  assign g10983 = \DFF_1505.Q ;
  assign g10988 = \DFF_1428.Q ;
  assign g10991 = \DFF_1427.Q ;
  assign g10994 = \DFF_1428.Q ;
  assign g10995 = \DFF_1505.Q ;
  assign g10996 = \DFF_1427.Q ;
  assign g10999 = \DFF_1428.Q ;
  assign g11 = \DFF_1628.Q ;
  assign g11002 = \DFF_1006.D ;
  assign g11003 = \DFF_1012.D ;
  assign g11004 = \DFF_1428.Q ;
  assign g11007 = \DFF_1494.D ;
  assign g11008 = \DFF_1506.Q ;
  assign g1101 = \DFF_617.Q ;
  assign g11011 = \DFF_1505.Q ;
  assign g11014 = \DFF_1506.Q ;
  assign g11017 = \DFF_1505.Q ;
  assign g11022 = \DFF_1429.Q ;
  assign g11025 = \DFF_1428.Q ;
  assign g11028 = \DFF_1427.Q ;
  assign g11031 = \DFF_308.D ;
  assign g11035 = \DFF_1505.Q ;
  assign g11036 = \DFF_1428.Q ;
  assign g11039 = \DFF_1427.Q ;
  assign g1104 = \DFF_618.Q ;
  assign g11042 = \DFF_1428.Q ;
  assign g11045 = \DFF_1505.Q ;
  assign g11048 = \DFF_1427.Q ;
  assign g11051 = \DFF_1428.Q ;
  assign g11054 = \DFF_1356.D ;
  assign g11055 = \DFF_1362.D ;
  assign g11056 = \DFF_1428.Q ;
  assign g11063 = \DFF_1506.Q ;
  assign g11066 = \DFF_1506.Q ;
  assign g11069 = \DFF_156.Q ;
  assign g1107 = \DFF_619.Q ;
  assign g11079 = \DFF_1429.Q ;
  assign g11082 = \DFF_1428.Q ;
  assign g11085 = \DFF_1427.Q ;
  assign g11091 = \DFF_1505.Q ;
  assign g11092 = \DFF_1429.Q ;
  assign g11095 = \DFF_1428.Q ;
  assign g11098 = \DFF_1427.Q ;
  assign g1110 = \DFF_620.Q ;
  assign g11101 = \DFF_658.D ;
  assign g11105 = \DFF_1505.Q ;
  assign g11108 = \DFF_1428.Q ;
  assign g11111 = \DFF_1427.Q ;
  assign g11114 = \DFF_1428.Q ;
  assign g11117 = \DFF_1505.Q ;
  assign g11120 = \DFF_1427.Q ;
  assign g11123 = \DFF_1428.Q ;
  assign g11126 = \DFF_1506.Q ;
  assign g11129 = \DFF_1506.Q ;
  assign g1113 = \DFF_623.Q ;
  assign g11132 = \DFF_1429.Q ;
  assign g11135 = \DFF_1428.Q ;
  assign g11138 = \DFF_1427.Q ;
  assign g1114 = \DFF_621.Q ;
  assign g11144 = \DFF_1505.Q ;
  assign g11145 = \DFF_1429.Q ;
  assign g11148 = \DFF_1428.Q ;
  assign g1115 = \DFF_622.Q ;
  assign g11151 = \DFF_1427.Q ;
  assign g11157 = \DFF_1505.Q ;
  assign g1116 = \DFF_624.Q ;
  assign g11160 = \DFF_1429.Q ;
  assign g11163 = \DFF_1428.Q ;
  assign g11166 = \DFF_1427.Q ;
  assign g11169 = \DFF_1008.D ;
  assign g11173 = \DFF_1505.Q ;
  assign g11176 = \DFF_1428.Q ;
  assign g11179 = \DFF_1427.Q ;
  assign g11182 = \DFF_1428.Q ;
  assign g11185 = \DFF_1505.Q ;
  assign g1119 = \DFF_625.Q ;
  assign g11190 = \DFF_159.Q ;
  assign g11199 = \DFF_1429.Q ;
  assign g11202 = \DFF_1428.Q ;
  assign g11205 = \DFF_1427.Q ;
  assign g11208 = \DFF_310.D ;
  assign g11209 = \DFF_1428.Q ;
  assign g11213 = \DFF_1505.Q ;
  assign g11216 = \DFF_1429.Q ;
  assign g11219 = \DFF_1428.Q ;
  assign g1122 = \DFF_626.Q ;
  assign g11222 = \DFF_1427.Q ;
  assign g11228 = \DFF_1505.Q ;
  assign g11231 = \DFF_1429.Q ;
  assign g11234 = \DFF_1428.Q ;
  assign g11237 = \DFF_1427.Q ;
  assign g11243 = \DFF_1505.Q ;
  assign g11246 = \DFF_1429.Q ;
  assign g11249 = \DFF_1428.Q ;
  assign g1125 = \DFF_627.Q ;
  assign g11252 = \DFF_1427.Q ;
  assign g11255 = \DFF_1358.D ;
  assign g11259 = \DFF_1505.Q ;
  assign g11265 = \DFF_1427.Q ;
  assign g11268 = \DFF_1429.Q ;
  assign g11271 = \DFF_1428.Q ;
  assign g11274 = \DFF_1427.Q ;
  assign g11277 = \DFF_1428.Q ;
  assign g1128 = \DFF_628.Q ;
  assign g11281 = \DFF_1429.Q ;
  assign g11284 = \DFF_1428.Q ;
  assign g11287 = \DFF_1427.Q ;
  assign g11290 = \DFF_660.D ;
  assign g11291 = \DFF_1428.Q ;
  assign g11297 = \DFF_1505.Q ;
  assign g113 = \DFF_72.Q ;
  assign g11300 = \DFF_1429.Q ;
  assign g11303 = \DFF_1428.Q ;
  assign g11306 = \DFF_1427.Q ;
  assign g1131 = \DFF_629.Q ;
  assign g11312 = \DFF_1505.Q ;
  assign g11315 = \DFF_1429.Q ;
  assign g11318 = \DFF_1428.Q ;
  assign g11321 = \DFF_1427.Q ;
  assign g11327 = \DFF_1505.Q ;
  assign g11332 = \DFF_158.Q ;
  assign g1134 = \DFF_632.Q ;
  assign g11341 = \DFF_1428.Q ;
  assign g11344 = \DFF_1427.Q ;
  assign g11348 = \DFF_1429.Q ;
  assign g1135 = \DFF_630.Q ;
  assign g11351 = \DFF_1428.Q ;
  assign g11354 = \DFF_1428.Q ;
  assign g11358 = \DFF_1427.Q ;
  assign g1136 = \DFF_631.Q ;
  assign g11361 = \DFF_1429.Q ;
  assign g11364 = \DFF_1428.Q ;
  assign g11367 = \DFF_1427.Q ;
  assign g1137 = \DFF_648.Q ;
  assign g11370 = \DFF_1428.Q ;
  assign g11376 = \DFF_1429.Q ;
  assign g11379 = \DFF_1428.Q ;
  assign g1138 = \DFF_649.Q ;
  assign g11382 = \DFF_1427.Q ;
  assign g11385 = \DFF_1010.D ;
  assign g11386 = \DFF_1428.Q ;
  assign g1139 = \DFF_650.Q ;
  assign g11392 = \DFF_1505.Q ;
  assign g11395 = \DFF_1429.Q ;
  assign g11398 = \DFF_1428.Q ;
  assign g1140 = \DFF_651.Q ;
  assign g11401 = \DFF_1427.Q ;
  assign g11407 = \DFF_1505.Q ;
  assign g1141 = \DFF_652.Q ;
  assign g11411 = \DFF_1429.Q ;
  assign g11414 = \DFF_1428.Q ;
  assign g11417 = \DFF_1427.Q ;
  assign g1142 = \DFF_733.Q ;
  assign g11422 = \DFF_1429.Q ;
  assign g11425 = \DFF_1428.Q ;
  assign g11428 = \DFF_1427.Q ;
  assign g11432 = \DFF_1429.Q ;
  assign g11435 = \DFF_1428.Q ;
  assign g11438 = \DFF_1428.Q ;
  assign g11444 = \DFF_1427.Q ;
  assign g11447 = \DFF_1429.Q ;
  assign g1145 = \DFF_734.Q ;
  assign g11450 = \DFF_1428.Q ;
  assign g11453 = \DFF_1427.Q ;
  assign g11456 = \DFF_1428.Q ;
  assign g11462 = \DFF_1429.Q ;
  assign g11465 = \DFF_1428.Q ;
  assign g11468 = \DFF_1427.Q ;
  assign g11471 = \DFF_1360.D ;
  assign g11472 = \DFF_1428.Q ;
  assign g11478 = \DFF_1505.Q ;
  assign g1148 = \DFF_735.Q ;
  assign g11481 = \DFF_157.Q ;
  assign g11490 = g51;
  assign g11491 = \DFF_304.D ;
  assign g11492 = \DFF_306.D ;
  assign g11493 = \DFF_308.D ;
  assign g11494 = \DFF_310.D ;
  assign g11495 = \DFF_312.D ;
  assign g11496 = \DFF_1297.Q ;
  assign g11497 = \DFF_253.Q ;
  assign g11498 = \DFF_254.Q ;
  assign g11499 = \DFF_255.Q ;
  assign g11500 = \DFF_256.Q ;
  assign g11501 = \DFF_257.Q ;
  assign g11502 = \DFF_258.Q ;
  assign g11503 = \DFF_259.Q ;
  assign g11504 = \DFF_260.Q ;
  assign g11505 = \DFF_261.Q ;
  assign g11506 = \DFF_262.Q ;
  assign g11507 = \DFF_263.Q ;
  assign g11508 = \DFF_264.Q ;
  assign g11509 = \DFF_298.D ;
  assign g1151 = \DFF_741.Q ;
  assign g11510 = \DFF_300.D ;
  assign g11511 = \DFF_302.D ;
  assign g11512 = \DFF_383.Q ;
  assign g11513 = \DFF_393.Q ;
  assign g11514 = \DFF_394.Q ;
  assign g11515 = \DFF_384.Q ;
  assign g11516 = \DFF_385.Q ;
  assign g11517 = \DFF_392.Q ;
  assign g11518 = \DFF_654.D ;
  assign g11519 = \DFF_656.D ;
  assign g1152 = \DFF_742.Q ;
  assign g11520 = \DFF_658.D ;
  assign g11521 = \DFF_660.D ;
  assign g11522 = \DFF_662.D ;
  assign g11523 = \DFF_1297.Q ;
  assign g11524 = \DFF_603.Q ;
  assign g11525 = \DFF_604.Q ;
  assign g11526 = \DFF_605.Q ;
  assign g11527 = \DFF_606.Q ;
  assign g11528 = \DFF_607.Q ;
  assign g11529 = \DFF_608.Q ;
  assign g11530 = \DFF_609.Q ;
  assign g11531 = \DFF_610.Q ;
  assign g11532 = \DFF_611.Q ;
  assign g11533 = \DFF_612.Q ;
  assign g11534 = \DFF_613.Q ;
  assign g11535 = \DFF_614.Q ;
  assign g11536 = \DFF_648.D ;
  assign g11537 = \DFF_650.D ;
  assign g11538 = \DFF_652.D ;
  assign g11539 = \DFF_733.Q ;
  assign g11540 = \DFF_743.Q ;
  assign g11541 = \DFF_744.Q ;
  assign g11542 = \DFF_734.Q ;
  assign g11543 = \DFF_735.Q ;
  assign g11544 = \DFF_742.Q ;
  assign g11545 = \DFF_1004.D ;
  assign g11546 = \DFF_1006.D ;
  assign g11547 = \DFF_1008.D ;
  assign g11548 = \DFF_1010.D ;
  assign g11549 = \DFF_1012.D ;
  assign g1155 = \DFF_743.Q ;
  assign g11550 = \DFF_1297.Q ;
  assign g11551 = \DFF_953.Q ;
  assign g11552 = \DFF_954.Q ;
  assign g11553 = \DFF_955.Q ;
  assign g11554 = \DFF_956.Q ;
  assign g11555 = \DFF_957.Q ;
  assign g11556 = \DFF_958.Q ;
  assign g11557 = \DFF_959.Q ;
  assign g11558 = \DFF_960.Q ;
  assign g11559 = \DFF_961.Q ;
  assign g11560 = \DFF_962.Q ;
  assign g11561 = \DFF_963.Q ;
  assign g11562 = \DFF_964.Q ;
  assign g11563 = \DFF_998.D ;
  assign g11564 = \DFF_1000.D ;
  assign g11565 = \DFF_1002.D ;
  assign g11566 = \DFF_1083.Q ;
  assign g11567 = \DFF_1093.Q ;
  assign g11568 = \DFF_1094.Q ;
  assign g11569 = \DFF_1084.Q ;
  assign g11570 = \DFF_1085.Q ;
  assign g11571 = \DFF_1092.Q ;
  assign g11572 = \DFF_1354.D ;
  assign g11573 = \DFF_1356.D ;
  assign g11574 = \DFF_1358.D ;
  assign g11575 = \DFF_1360.D ;
  assign g11576 = \DFF_1362.D ;
  assign g11577 = \DFF_1297.Q ;
  assign g11578 = \DFF_1303.Q ;
  assign g11579 = \DFF_1304.Q ;
  assign g1158 = \DFF_744.Q ;
  assign g11580 = \DFF_1305.Q ;
  assign g11581 = \DFF_1306.Q ;
  assign g11582 = \DFF_1307.Q ;
  assign g11583 = \DFF_1308.Q ;
  assign g11584 = \DFF_1309.Q ;
  assign g11585 = \DFF_1310.Q ;
  assign g11586 = \DFF_1311.Q ;
  assign g11587 = \DFF_1312.Q ;
  assign g11588 = \DFF_1313.Q ;
  assign g11589 = \DFF_1314.Q ;
  assign g11590 = \DFF_1348.D ;
  assign g11591 = \DFF_1350.D ;
  assign g11592 = \DFF_1352.D ;
  assign g11593 = \DFF_1433.Q ;
  assign g11594 = \DFF_1443.Q ;
  assign g11595 = \DFF_1444.Q ;
  assign g11596 = \DFF_1434.Q ;
  assign g11597 = \DFF_1435.Q ;
  assign g11598 = \DFF_1442.Q ;
  assign g11599 = \DFF_448.D ;
  assign g11603 = \DFF_782.Q ;
  assign g11606 = \DFF_797.D ;
  assign g11608 = \DFF_1132.Q ;
  assign g1161 = \DFF_1427.Q ;
  assign g11611 = \DFF_1146.D ;
  assign g11613 = \DFF_1482.Q ;
  assign g11616 = \DFF_1495.D ;
  assign g11623 = g3230;
  assign g11628 = \DFF_449.D ;
  assign g11629 = \DFF_798.D ;
  assign g11633 = \DFF_1132.Q ;
  assign g11636 = \DFF_1147.D ;
  assign g11638 = \DFF_1482.Q ;
  assign g1164 = \DFF_736.Q ;
  assign g11641 = \DFF_1496.D ;
  assign g1165 = \DFF_737.Q ;
  assign g11651 = \DFF_799.D ;
  assign g11652 = \DFF_1148.D ;
  assign g11656 = \DFF_1482.Q ;
  assign g11659 = \DFF_1497.D ;
  assign g1166 = \DFF_738.Q ;
  assign g1167 = \DFF_739.Q ;
  assign g11670 = \DFF_1149.D ;
  assign g11671 = \DFF_1498.D ;
  assign g1168 = \DFF_1428.Q ;
  assign g11682 = \DFF_1499.D ;
  assign g117 = \DFF_70.Q ;
  assign g11706 = g3233;
  assign g1171 = \DFF_740.Q ;
  assign g11713 = \DFF_1613.D ;
  assign g1172 = \DFF_1429.Q ;
  assign g1173 = \DFF_730.Q ;
  assign g11737 = g3231;
  assign g1174 = \DFF_731.Q ;
  assign g11743 = g3232;
  assign g1175 = \DFF_732.Q ;
  assign g11758 = g3220;
  assign g1176 = \DFF_726.Q ;
  assign g11766 = g3219;
  assign g11769 = \DFF_3.Q ;
  assign g1177 = \DFF_779.Q ;
  assign g11779 = g3218;
  assign g11786 = \DFF_3.Q ;
  assign g11798 = g3217;
  assign g1180 = \DFF_780.Q ;
  assign g11812 = \DFF_3.Q ;
  assign g11821 = g3216;
  assign g11827 = \DFF_316.Q ;
  assign g1183 = \DFF_781.Q ;
  assign g11845 = \DFF_3.Q ;
  assign g11854 = g3215;
  assign g11859 = \DFF_316.Q ;
  assign g1186 = \DFF_752.Q ;
  assign g11869 = \DFF_666.Q ;
  assign g11888 = g3214;
  assign g11894 = \DFF_316.Q ;
  assign g11901 = \DFF_666.Q ;
  assign g11911 = \DFF_1016.Q ;
  assign g1192 = \DFF_782.Q ;
  assign g11927 = g3213;
  assign g1193 = \DFF_783.Q ;
  assign g11933 = \DFF_316.Q ;
  assign g11937 = \DFF_1563.Q ;
  assign g11944 = \DFF_666.Q ;
  assign g11951 = \DFF_1016.Q ;
  assign g1196 = \DFF_711.Q ;
  assign g11961 = \DFF_1366.Q ;
  assign g11973 = \DFF_316.Q ;
  assign g11976 = \DFF_1429.Q ;
  assign g11986 = \DFF_666.Q ;
  assign g1199 = \DFF_712.Q ;
  assign g11990 = \DFF_1563.Q ;
  assign g11997 = \DFF_1016.Q ;
  assign g12004 = \DFF_1366.Q ;
  assign g12025 = \DFF_316.Q ;
  assign g12027 = \DFF_1427.Q ;
  assign g12030 = \DFF_1428.Q ;
  assign g12042 = \DFF_666.Q ;
  assign g12045 = \DFF_1429.Q ;
  assign g12055 = \DFF_1016.Q ;
  assign g12059 = \DFF_1563.Q ;
  assign g1206 = \DFF_792.Q ;
  assign g12066 = \DFF_1366.Q ;
  assign g12089 = \DFF_666.Q ;
  assign g1209 = \DFF_713.Q ;
  assign g12091 = \DFF_1427.Q ;
  assign g12094 = \DFF_1428.Q ;
  assign g121 = \DFF_68.Q ;
  assign g1210 = \DFF_714.Q ;
  assign g12106 = \DFF_1016.Q ;
  assign g12109 = \DFF_1429.Q ;
  assign g1211 = \DFF_793.Q ;
  assign g12119 = \DFF_1366.Q ;
  assign g12123 = \DFF_1563.Q ;
  assign g12136 = \DFF_1427.Q ;
  assign g12139 = \DFF_1428.Q ;
  assign g1214 = \DFF_745.Q ;
  assign g12142 = \DFF_1429.Q ;
  assign g1215 = \DFF_794.Q ;
  assign g1216 = \DFF_795.Q ;
  assign g12161 = \DFF_1016.Q ;
  assign g12163 = \DFF_1427.Q ;
  assign g12166 = \DFF_1428.Q ;
  assign g1217 = \DFF_796.Q ;
  assign g12178 = \DFF_1366.Q ;
  assign g1218 = \DFF_797.Q ;
  assign g12181 = \DFF_1429.Q ;
  assign g1219 = \DFF_798.Q ;
  assign g12198 = \DFF_1427.Q ;
  assign g1220 = \DFF_799.Q ;
  assign g12201 = \DFF_1428.Q ;
  assign g12204 = \DFF_1429.Q ;
  assign g1221 = \DFF_746.Q ;
  assign g1222 = \DFF_800.Q ;
  assign g12223 = \DFF_1366.Q ;
  assign g12225 = \DFF_1427.Q ;
  assign g12228 = \DFF_1428.Q ;
  assign g1223 = \DFF_801.Q ;
  assign g12239 = \DFF_1428.Q ;
  assign g1224 = \DFF_802.Q ;
  assign g12242 = \DFF_1429.Q ;
  assign g12253 = \DFF_1427.Q ;
  assign g12256 = \DFF_1428.Q ;
  assign g12259 = \DFF_1429.Q ;
  assign g1227 = \DFF_803.Q ;
  assign g12279 = \DFF_1427.Q ;
  assign g1228 = \DFF_747.Q ;
  assign g12282 = \DFF_1428.Q ;
  assign g12285 = \DFF_1429.Q ;
  assign g1229 = \DFF_748.Q ;
  assign g12296 = \DFF_1427.Q ;
  assign g12299 = \DFF_1428.Q ;
  assign g1230 = \DFF_749.Q ;
  assign g12302 = \DFF_1429.Q ;
  assign g1231 = \DFF_1504.Q ;
  assign g12312 = \DFF_1429.Q ;
  assign g12315 = \DFF_1427.Q ;
  assign g12318 = \DFF_1428.Q ;
  assign g12321 = \DFF_1429.Q ;
  assign g12332 = g3212;
  assign g12333 = \DFF_1427.Q ;
  assign g12336 = \DFF_1428.Q ;
  assign g1234 = \DFF_750.Q ;
  assign g12340 = \DFF_1429.Q ;
  assign g12343 = \DFF_1427.Q ;
  assign g12346 = \DFF_1428.Q ;
  assign g12349 = \DFF_1429.Q ;
  assign g1235 = \DFF_751.Q ;
  assign g1236 = \DFF_1506.Q ;
  assign g12362 = g3228;
  assign g12363 = \DFF_1427.Q ;
  assign g12366 = \DFF_1428.Q ;
  assign g1237 = \DFF_1505.Q ;
  assign g12370 = \DFF_1429.Q ;
  assign g12373 = \DFF_1427.Q ;
  assign g12378 = g3227;
  assign g12379 = \DFF_1429.Q ;
  assign g12382 = \DFF_1427.Q ;
  assign g12385 = \DFF_1428.Q ;
  assign g12389 = \DFF_1429.Q ;
  assign g1240 = \DFF_709.Q ;
  assign g12408 = g3226;
  assign g12409 = \DFF_1429.Q ;
  assign g12412 = \DFF_1427.Q ;
  assign g12415 = \DFF_1428.Q ;
  assign g12420 = g3225;
  assign g12421 = \DFF_1429.Q ;
  assign g12424 = g3224;
  assign g12425 = \DFF_3.Q ;
  assign g12426 = \DFF_1429.Q ;
  assign g1243 = \DFF_710.Q ;
  assign g12430 = g3223;
  assign g12432 = \DFF_3.Q ;
  assign g12433 = \DFF_19.D ;
  assign g12434 = g3222;
  assign g12435 = \DFF_1563.Q ;
  assign g12437 = \DFF_3.Q ;
  assign g12438 = g3221;
  assign g1244 = \DFF_753.Q ;
  assign g12440 = \DFF_1563.Q ;
  assign g12442 = \DFF_3.Q ;
  assign g12445 = \DFF_1563.Q ;
  assign g1245 = \DFF_754.Q ;
  assign g12450 = \DFF_1563.Q ;
  assign g12457 = \DFF_395.D ;
  assign g12467 = \DFF_745.D ;
  assign g1248 = g1249;
  assign g12482 = \DFF_1095.D ;
  assign g12487 = \DFF_362.D ;
  assign g12499 = \DFF_1445.D ;
  assign g125 = \DFF_66.Q ;
  assign g1250 = \DFF_715.Q ;
  assign g12507 = \DFF_712.D ;
  assign g1251 = \DFF_722.Q ;
  assign g12519 = \DFF_3.Q ;
  assign g1252 = \DFF_723.Q ;
  assign g12524 = \DFF_1062.D ;
  assign g1253 = \DFF_724.Q ;
  assign g12534 = \DFF_3.Q ;
  assign g12539 = \DFF_1412.D ;
  assign g1254 = \DFF_725.Q ;
  assign g12543 = \DFF_3.Q ;
  assign g1255 = \DFF_716.Q ;
  assign g12552 = \DFF_3.Q ;
  assign g1256 = \DFF_717.Q ;
  assign g12564 = \DFF_157.Q ;
  assign g12565 = \DFF_1302.Q ;
  assign g1257 = \DFF_718.Q ;
  assign g1258 = \DFF_719.Q ;
  assign g1259 = \DFF_720.Q ;
  assign g1260 = \DFF_721.Q ;
  assign g12607 = \DFF_157.Q ;
  assign g12608 = \DFF_1427.Q ;
  assign g1261 = \DFF_757.Q ;
  assign g12611 = \DFF_1302.Q ;
  assign g1262 = \DFF_755.Q ;
  assign g1263 = \DFF_756.Q ;
  assign g1264 = \DFF_760.Q ;
  assign g1265 = \DFF_758.Q ;
  assign g12654 = \DFF_1427.Q ;
  assign g12657 = \DFF_1302.Q ;
  assign g1266 = \DFF_759.Q ;
  assign g1267 = \DFF_763.Q ;
  assign g1268 = \DFF_761.Q ;
  assign g1269 = \DFF_762.Q ;
  assign g12699 = \DFF_1428.Q ;
  assign g1270 = \DFF_766.Q ;
  assign g12708 = \DFF_1427.Q ;
  assign g1271 = \DFF_764.Q ;
  assign g12711 = \DFF_1302.Q ;
  assign g1272 = \DFF_765.Q ;
  assign g1273 = \DFF_767.Q ;
  assign g12756 = \DFF_1428.Q ;
  assign g1276 = \DFF_768.Q ;
  assign g12765 = \DFF_1427.Q ;
  assign g1279 = \DFF_769.Q ;
  assign g12798 = \DFF_1428.Q ;
  assign g12811 = \DFF_1563.Q ;
  assign g1282 = \DFF_770.Q ;
  assign g12837 = \DFF_1428.Q ;
  assign g1285 = \DFF_771.Q ;
  assign g1288 = \DFF_772.Q ;
  assign g129 = \DFF_166.Q ;
  assign g12909 = g3234;
  assign g1291 = \DFF_776.Q ;
  assign g1294 = \DFF_777.Q ;
  assign g12962 = \DFF_3.Q ;
  assign g1297 = \DFF_778.Q ;
  assign g130 = \DFF_164.Q ;
  assign g1300 = \DFF_773.Q ;
  assign g1303 = \DFF_774.Q ;
  assign g1306 = \DFF_775.Q ;
  assign g13070 = \DFF_1563.Q ;
  assign g1309 = \DFF_1504.Q ;
  assign g131 = \DFF_165.Q ;
  assign g13110 = \DFF_1296.D ;
  assign g13111 = \DFF_401.D ;
  assign g1312 = \DFF_1505.Q ;
  assign g13124 = \DFF_751.D ;
  assign g13135 = \DFF_1101.D ;
  assign g13143 = \DFF_1451.D ;
  assign g13149 = \DFF_398.D ;
  assign g1315 = \DFF_1506.Q ;
  assign g13155 = \DFF_748.D ;
  assign g1316 = \DFF_807.Q ;
  assign g13160 = \DFF_403.D ;
  assign g13164 = \DFF_1098.D ;
  assign g13171 = \DFF_753.D ;
  assign g13175 = \DFF_1448.D ;
  assign g13182 = \DFF_1103.D ;
  assign g1319 = \DFF_810.Q ;
  assign g13194 = \DFF_1453.D ;
  assign g132 = \DFF_169.Q ;
  assign g13215 = \DFF_432.Q ;
  assign g13229 = \DFF_432.Q ;
  assign g13234 = \DFF_782.Q ;
  assign g13246 = \DFF_82.Q ;
  assign g13248 = \DFF_450.D ;
  assign g13252 = \DFF_782.Q ;
  assign g13257 = \DFF_1132.Q ;
  assign g1326 = \DFF_809.Q ;
  assign g13265 = g3229;
  assign g13267 = \DFF_451.D ;
  assign g13269 = \DFF_64.Q ;
  assign g13271 = \DFF_800.D ;
  assign g13275 = \DFF_1132.Q ;
  assign g13280 = \DFF_1482.Q ;
  assign g13290 = \DFF_453.D ;
  assign g13292 = \DFF_801.D ;
  assign g13294 = \DFF_46.Q ;
  assign g13296 = \DFF_1150.D ;
  assign g133 = \DFF_167.Q ;
  assign g13300 = \DFF_1482.Q ;
  assign g13317 = \DFF_1563.Q ;
  assign g13318 = \DFF_1505.Q ;
  assign g13319 = \DFF_444.D ;
  assign g1332 = \DFF_812.Q ;
  assign g13321 = \DFF_803.D ;
  assign g13323 = \DFF_1151.D ;
  assign g13325 = \DFF_91.Q ;
  assign g13327 = \DFF_1500.D ;
  assign g13336 = \DFF_432.Q ;
  assign g13339 = \DFF_445.D ;
  assign g13341 = \DFF_1563.Q ;
  assign g13342 = \DFF_794.D ;
  assign g13344 = \DFF_1153.D ;
  assign g13346 = \DFF_1501.D ;
  assign g13356 = \DFF_432.Q ;
  assign g13359 = \DFF_446.D ;
  assign g13361 = \DFF_782.Q ;
  assign g13364 = \DFF_795.D ;
  assign g13366 = \DFF_1563.Q ;
  assign g13367 = \DFF_1144.D ;
  assign g13369 = \DFF_1503.D ;
  assign g13381 = \DFF_432.Q ;
  assign g13384 = \DFF_447.D ;
  assign g13386 = \DFF_782.Q ;
  assign g13389 = \DFF_796.D ;
  assign g1339 = \DFF_811.Q ;
  assign g13391 = \DFF_1132.Q ;
  assign g13394 = \DFF_1145.D ;
  assign g13396 = \DFF_1563.Q ;
  assign g13397 = \DFF_1494.D ;
  assign g134 = \DFF_168.Q ;
  assign g13405 = \DFF_3.Q ;
  assign g13406 = \DFF_3.Q ;
  assign g13407 = \DFF_82.Q ;
  assign g13408 = \DFF_1563.Q ;
  assign g13409 = \DFF_3.Q ;
  assign g13410 = \DFF_444.D ;
  assign g13411 = \DFF_445.D ;
  assign g13412 = \DFF_446.D ;
  assign g13413 = \DFF_447.D ;
  assign g13414 = \DFF_448.D ;
  assign g13415 = \DFF_449.D ;
  assign g13416 = \DFF_450.D ;
  assign g13417 = \DFF_451.D ;
  assign g13418 = \DFF_453.D ;
  assign g13419 = \DFF_1563.Q ;
  assign g13420 = \DFF_1563.Q ;
  assign g13421 = \DFF_3.Q ;
  assign g13422 = \DFF_3.Q ;
  assign g13423 = \DFF_64.Q ;
  assign g13424 = \DFF_1563.Q ;
  assign g13425 = \DFF_3.Q ;
  assign g13426 = \DFF_794.D ;
  assign g13427 = \DFF_795.D ;
  assign g13428 = \DFF_796.D ;
  assign g13429 = \DFF_797.D ;
  assign g13430 = \DFF_798.D ;
  assign g13431 = \DFF_799.D ;
  assign g13432 = \DFF_800.D ;
  assign g13433 = \DFF_801.D ;
  assign g13434 = \DFF_803.D ;
  assign g13435 = \DFF_1563.Q ;
  assign g13436 = \DFF_1563.Q ;
  assign g13437 = \DFF_3.Q ;
  assign g13438 = \DFF_3.Q ;
  assign g13439 = \DFF_46.Q ;
  assign g13440 = \DFF_1563.Q ;
  assign g13441 = \DFF_3.Q ;
  assign g13442 = \DFF_1144.D ;
  assign g13443 = \DFF_1145.D ;
  assign g13444 = \DFF_1146.D ;
  assign g13445 = \DFF_1147.D ;
  assign g13446 = \DFF_1148.D ;
  assign g13447 = \DFF_1149.D ;
  assign g13448 = \DFF_1150.D ;
  assign g13449 = \DFF_1151.D ;
  assign g1345 = \DFF_808.Q ;
  assign g13450 = \DFF_1153.D ;
  assign g13451 = \DFF_1563.Q ;
  assign g13452 = \DFF_1563.Q ;
  assign g13453 = \DFF_3.Q ;
  assign g13454 = \DFF_3.Q ;
  assign g13455 = \DFF_91.Q ;
  assign g13456 = \DFF_1563.Q ;
  assign g13457 = \DFF_3.Q ;
  assign g13458 = \DFF_1494.D ;
  assign g13459 = \DFF_1495.D ;
  assign g1346 = \DFF_813.Q ;
  assign g13460 = \DFF_1496.D ;
  assign g13461 = \DFF_1497.D ;
  assign g13462 = \DFF_1498.D ;
  assign g13463 = \DFF_1499.D ;
  assign g13464 = \DFF_1500.D ;
  assign g13465 = \DFF_1501.D ;
  assign g13466 = \DFF_1503.D ;
  assign g13467 = \DFF_1563.Q ;
  assign g13468 = \DFF_1563.Q ;
  assign g13469 = g51;
  assign g13475 = \DFF_1563.Q ;
  assign g135 = \DFF_1428.Q ;
  assign g1352 = \DFF_815.Q ;
  assign g13571 = \DFF_398.D ;
  assign g13572 = \DFF_401.D ;
  assign g13579 = \DFF_748.D ;
  assign g1358 = \DFF_814.Q ;
  assign g13580 = \DFF_403.D ;
  assign g13581 = \DFF_751.D ;
  assign g13588 = \DFF_1098.D ;
  assign g13589 = g3229;
  assign g13598 = \DFF_362.D ;
  assign g13600 = \DFF_753.D ;
  assign g13601 = \DFF_1101.D ;
  assign g13608 = \DFF_1448.D ;
  assign g13610 = \DFF_712.D ;
  assign g13612 = \DFF_1103.D ;
  assign g13613 = \DFF_1451.D ;
  assign g13620 = \DFF_1062.D ;
  assign g13622 = \DFF_1453.D ;
  assign g13624 = \DFF_395.D ;
  assign g13632 = \DFF_1412.D ;
  assign g13635 = \DFF_745.D ;
  assign g13647 = \DFF_1095.D ;
  assign g1365 = \DFF_816.Q ;
  assign g13673 = \DFF_1445.D ;
  assign g1372 = \DFF_817.Q ;
  assign g1378 = \DFF_818.Q ;
  assign g138 = \DFF_1427.Q ;
  assign g1384 = \DFF_821.Q ;
  assign g1385 = \DFF_819.Q ;
  assign g1386 = \DFF_820.Q ;
  assign g13863 = \DFF_1613.D ;
  assign g1387 = \DFF_824.Q ;
  assign g1388 = \DFF_822.Q ;
  assign g1389 = \DFF_823.Q ;
  assign g1390 = \DFF_827.Q ;
  assign g1391 = \DFF_825.Q ;
  assign g1392 = \DFF_826.Q ;
  assign g1393 = \DFF_830.Q ;
  assign g1394 = \DFF_828.Q ;
  assign g1395 = \DFF_829.Q ;
  assign g1396 = \DFF_833.Q ;
  assign g1397 = \DFF_831.Q ;
  assign g1398 = \DFF_832.Q ;
  assign g1399 = \DFF_836.Q ;
  assign g14 = \DFF_1629.Q ;
  assign g1400 = \DFF_834.Q ;
  assign g1401 = \DFF_835.Q ;
  assign g1402 = \DFF_839.Q ;
  assign g1403 = \DFF_837.Q ;
  assign g1404 = \DFF_838.Q ;
  assign g1405 = \DFF_842.Q ;
  assign g1406 = \DFF_840.Q ;
  assign g1407 = \DFF_841.Q ;
  assign g1408 = \DFF_845.Q ;
  assign g1409 = \DFF_843.Q ;
  assign g141 = \DFF_172.Q ;
  assign g1410 = \DFF_844.Q ;
  assign g1411 = \DFF_848.Q ;
  assign g1412 = \DFF_846.Q ;
  assign g1413 = \DFF_847.Q ;
  assign g1414 = \DFF_851.Q ;
  assign g1415 = \DFF_849.Q ;
  assign g1416 = \DFF_850.Q ;
  assign g1417 = \DFF_854.Q ;
  assign g1418 = \DFF_852.Q ;
  assign g1419 = \DFF_853.Q ;
  assign g142 = \DFF_170.Q ;
  assign g1420 = \DFF_857.Q ;
  assign g1421 = \DFF_855.Q ;
  assign g1422 = \DFF_856.Q ;
  assign g1423 = \DFF_860.Q ;
  assign g1424 = \DFF_858.Q ;
  assign g1425 = \DFF_859.Q ;
  assign g1426 = \DFF_945.Q ;
  assign g143 = \DFF_171.Q ;
  assign g1430 = \DFF_944.Q ;
  assign g14337 = \DFF_1296.D ;
  assign g1435 = \DFF_943.Q ;
  assign g1439 = \DFF_942.Q ;
  assign g144 = \DFF_175.Q ;
  assign g1444 = \DFF_941.Q ;
  assign g1448 = \DFF_940.Q ;
  assign g145 = \DFF_173.Q ;
  assign g1453 = \DFF_939.Q ;
  assign g1457 = \DFF_938.Q ;
  assign g146 = \DFF_174.Q ;
  assign g1462 = \DFF_937.Q ;
  assign g1466 = \DFF_936.Q ;
  assign g14684 = \DFF_1613.D ;
  assign g147 = \DFF_178.Q ;
  assign g1471 = \DFF_45.Q ;
  assign g14718 = g3223;
  assign g14745 = g3222;
  assign g14746 = g3214;
  assign g1476 = \DFF_44.Q ;
  assign g14764 = \DFF_19.Q ;
  assign g14765 = g3221;
  assign g14766 = g3213;
  assign g14774 = g3212;
  assign g14775 = g3232;
  assign g14794 = \DFF_19.Q ;
  assign g14795 = g3228;
  assign g14796 = g3220;
  assign g148 = \DFF_176.Q ;
  assign g1481 = \DFF_43.Q ;
  assign g14829 = g3227;
  assign g14830 = g3219;
  assign g1486 = \DFF_42.Q ;
  assign g14881 = \DFF_19.Q ;
  assign g14882 = g3226;
  assign g14883 = g3218;
  assign g14885 = \DFF_316.D ;
  assign g149 = \DFF_177.Q ;
  assign g1491 = \DFF_41.Q ;
  assign g14954 = g3225;
  assign g14955 = g3217;
  assign g1496 = \DFF_40.Q ;
  assign g14966 = \DFF_666.D ;
  assign g150 = \DFF_181.Q ;
  assign g1501 = \DFF_39.Q ;
  assign g15017 = \DFF_19.Q ;
  assign g15018 = g3224;
  assign g15019 = g3216;
  assign g15055 = \DFF_1016.D ;
  assign g1506 = \DFF_38.Q ;
  assign g15092 = g3215;
  assign g151 = \DFF_179.Q ;
  assign g1511 = \DFF_866.Q ;
  assign g1512 = \DFF_864.Q ;
  assign g1513 = \DFF_865.Q ;
  assign g1514 = \DFF_869.Q ;
  assign g1515 = \DFF_867.Q ;
  assign g15151 = \DFF_1366.D ;
  assign g1516 = \DFF_868.Q ;
  assign g1517 = \DFF_1428.Q ;
  assign g15170 = \DFF_19.Q ;
  assign g152 = \DFF_180.Q ;
  assign g1520 = \DFF_1427.Q ;
  assign g1523 = \DFF_872.Q ;
  assign g1524 = \DFF_870.Q ;
  assign g1525 = \DFF_871.Q ;
  assign g1526 = \DFF_875.Q ;
  assign g1527 = \DFF_873.Q ;
  assign g1528 = \DFF_874.Q ;
  assign g1529 = \DFF_878.Q ;
  assign g153 = \DFF_184.Q ;
  assign g1530 = \DFF_876.Q ;
  assign g1531 = \DFF_877.Q ;
  assign g1532 = \DFF_881.Q ;
  assign g1533 = \DFF_879.Q ;
  assign g1534 = \DFF_880.Q ;
  assign g1535 = \DFF_884.Q ;
  assign g1536 = \DFF_882.Q ;
  assign g1537 = \DFF_883.Q ;
  assign g1538 = \DFF_887.Q ;
  assign g1539 = \DFF_885.Q ;
  assign g154 = \DFF_182.Q ;
  assign g1540 = \DFF_886.Q ;
  assign g1541 = \DFF_890.Q ;
  assign g1542 = \DFF_888.Q ;
  assign g1543 = \DFF_889.Q ;
  assign g1544 = \DFF_893.Q ;
  assign g1545 = \DFF_891.Q ;
  assign g1546 = \DFF_892.Q ;
  assign g1547 = \DFF_1429.Q ;
  assign g155 = \DFF_183.Q ;
  assign g1550 = \DFF_896.Q ;
  assign g1551 = \DFF_894.Q ;
  assign g1552 = \DFF_895.Q ;
  assign g1553 = \DFF_899.Q ;
  assign g1554 = \DFF_897.Q ;
  assign g1555 = \DFF_898.Q ;
  assign g1556 = \DFF_902.Q ;
  assign g1557 = \DFF_900.Q ;
  assign g1558 = \DFF_901.Q ;
  assign g1559 = \DFF_905.Q ;
  assign g156 = \DFF_187.Q ;
  assign g1560 = \DFF_903.Q ;
  assign g1561 = \DFF_904.Q ;
  assign g1562 = \DFF_1296.Q ;
  assign g1563 = \DFF_1302.Q ;
  assign g1564 = \DFF_1297.Q ;
  assign g1567 = \DFF_906.Q ;
  assign g157 = \DFF_185.Q ;
  assign g1570 = \DFF_907.Q ;
  assign g1573 = \DFF_908.Q ;
  assign g1576 = \DFF_912.Q ;
  assign g1579 = \DFF_913.Q ;
  assign g158 = \DFF_186.Q ;
  assign g1582 = \DFF_914.Q ;
  assign g1585 = \DFF_918.Q ;
  assign g15876 = g3234;
  assign g1588 = \DFF_919.Q ;
  assign g159 = \DFF_190.Q ;
  assign g1591 = \DFF_920.Q ;
  assign g1594 = \DFF_924.Q ;
  assign g1597 = \DFF_925.Q ;
  assign g15989 = \DFF_19.D ;
  assign g15991 = \DFF_19.Q ;
  assign g15994 = \DFF_19.Q ;
  assign g15997 = \DFF_19.Q ;
  assign g160 = \DFF_188.Q ;
  assign g1600 = \DFF_926.Q ;
  assign g16001 = \DFF_19.Q ;
  assign g16002 = \DFF_19.Q ;
  assign g16007 = \DFF_19.Q ;
  assign g16013 = \DFF_19.Q ;
  assign g16014 = \DFF_19.Q ;
  assign g16027 = \DFF_19.Q ;
  assign g1603 = \DFF_930.Q ;
  assign g16043 = \DFF_19.Q ;
  assign g16044 = \DFF_19.Q ;
  assign g1606 = \DFF_931.Q ;
  assign g16064 = \DFF_19.Q ;
  assign g1609 = \DFF_932.Q ;
  assign g16099 = \DFF_19.Q ;
  assign g161 = \DFF_189.Q ;
  assign g1612 = \DFF_909.Q ;
  assign g16132 = \DFF_16.D ;
  assign g1615 = \DFF_910.Q ;
  assign g1618 = \DFF_911.Q ;
  assign g16181 = \DFF_15.D ;
  assign g162 = \DFF_193.Q ;
  assign g1621 = \DFF_915.Q ;
  assign g1624 = \DFF_916.Q ;
  assign g1627 = \DFF_917.Q ;
  assign g16297 = \DFF_442.Q ;
  assign g163 = \DFF_191.Q ;
  assign g1630 = \DFF_921.Q ;
  assign g1633 = \DFF_922.Q ;
  assign g16355 = \DFF_792.Q ;
  assign g1636 = \DFF_923.Q ;
  assign g1639 = \DFF_927.Q ;
  assign g16399 = \DFF_1142.Q ;
  assign g164 = \DFF_192.Q ;
  assign g1642 = \DFF_928.Q ;
  assign g16437 = \DFF_1492.Q ;
  assign g1645 = \DFF_929.Q ;
  assign g16467 = \DFF_362.D ;
  assign g16468 = \DFF_395.D ;
  assign g16469 = \DFF_712.D ;
  assign g16470 = \DFF_745.D ;
  assign g16471 = \DFF_1062.D ;
  assign g16472 = \DFF_1095.D ;
  assign g16473 = \DFF_1412.D ;
  assign g16474 = \DFF_1445.D ;
  assign g16475 = g51;
  assign g16476 = g3212;
  assign g16477 = g3228;
  assign g16478 = g3227;
  assign g16479 = g3226;
  assign g1648 = \DFF_933.Q ;
  assign g16480 = g3225;
  assign g16481 = g3224;
  assign g16482 = g3223;
  assign g16483 = g3222;
  assign g16484 = g3221;
  assign g16485 = g3232;
  assign g16486 = g3220;
  assign g16487 = g3219;
  assign g16488 = g3218;
  assign g16489 = g3217;
  assign g16490 = g3216;
  assign g16491 = g3215;
  assign g16492 = g3214;
  assign g16493 = g3213;
  assign g16494 = \DFF_19.D ;
  assign g16495 = \DFF_1613.D ;
  assign g16496 = \DFF_1613.D ;
  assign g16497 = g3234;
  assign g165 = \DFF_1429.Q ;
  assign g16506 = \DFF_666.D ;
  assign g1651 = \DFF_934.Q ;
  assign g16528 = \DFF_1016.D ;
  assign g1654 = \DFF_935.Q ;
  assign g16559 = \DFF_1366.D ;
  assign g16566 = \DFF_1623.D ;
  assign g1657 = \DFF_1427.Q ;
  assign g1660 = \DFF_1003.Q ;
  assign g1661 = \DFF_1004.Q ;
  assign g1662 = \DFF_1005.Q ;
  assign g1663 = \DFF_1006.Q ;
  assign g1664 = \DFF_1007.Q ;
  assign g1665 = \DFF_1008.Q ;
  assign g16654 = \DFF_457.D ;
  assign g1666 = \DFF_1009.Q ;
  assign g1667 = \DFF_1010.Q ;
  assign g16671 = \DFF_807.D ;
  assign g1668 = \DFF_1011.Q ;
  assign g1669 = \DFF_1012.Q ;
  assign g16692 = \DFF_1157.D ;
  assign g1670 = \DFF_1013.Q ;
  assign g1671 = \DFF_1014.Q ;
  assign g16718 = \DFF_1507.D ;
  assign g1672 = \DFF_1015.Q ;
  assign g1679 = \DFF_1028.Q ;
  assign g168 = \DFF_196.Q ;
  assign g1680 = \DFF_1016.Q ;
  assign g16802 = \DFF_1.D ;
  assign g16803 = \DFF_1618.D ;
  assign g16813 = \DFF_401.D ;
  assign g16823 = \DFF_2.D ;
  assign g16824 = \DFF_1614.D ;
  assign g16831 = \DFF_751.D ;
  assign g16835 = \DFF_1619.D ;
  assign g16843 = \DFF_1101.D ;
  assign g16844 = \DFF_1615.D ;
  assign g16845 = \DFF_1625.D ;
  assign g16849 = \DFF_1451.D ;
  assign g16851 = \DFF_1620.D ;
  assign g16853 = \DFF_1616.D ;
  assign g16854 = \DFF_1626.D ;
  assign g16857 = \DFF_1621.D ;
  assign g16858 = \DFF_398.D ;
  assign g1686 = \DFF_1017.Q ;
  assign g16860 = \DFF_1617.D ;
  assign g16861 = \DFF_1627.D ;
  assign g16862 = \DFF_403.D ;
  assign g16863 = \DFF_748.D ;
  assign g16866 = \DFF_1622.D ;
  assign g16877 = \DFF_753.D ;
  assign g16878 = \DFF_1098.D ;
  assign g16880 = \DFF_1628.D ;
  assign g16881 = \DFF_316.D ;
  assign g169 = \DFF_194.Q ;
  assign g1690 = \DFF_1302.Q ;
  assign g16905 = \DFF_1103.D ;
  assign g16906 = \DFF_1448.D ;
  assign g16910 = \DFF_666.D ;
  assign g1693 = \DFF_983.Q ;
  assign g16934 = \DFF_1453.D ;
  assign g1694 = \DFF_984.Q ;
  assign g16940 = \DFF_1016.D ;
  assign g1695 = \DFF_985.Q ;
  assign g1696 = \DFF_986.Q ;
  assign g1697 = \DFF_987.Q ;
  assign g16971 = \DFF_1366.D ;
  assign g1698 = \DFF_988.Q ;
  assign g1699 = \DFF_989.Q ;
  assign g17 = \DFF_1627.Q ;
  assign g170 = \DFF_195.Q ;
  assign g1700 = \DFF_990.Q ;
  assign g1701 = \DFF_991.Q ;
  assign g1702 = \DFF_994.Q ;
  assign g1703 = \DFF_992.Q ;
  assign g1704 = \DFF_993.Q ;
  assign g1705 = \DFF_1052.Q ;
  assign g1706 = \DFF_1504.Q ;
  assign g171 = \DFF_199.Q ;
  assign g1712 = \DFF_1505.Q ;
  assign g1718 = \DFF_1506.Q ;
  assign g172 = \DFF_197.Q ;
  assign g17222 = \DFF_98.D ;
  assign g17224 = \DFF_101.D ;
  assign g17225 = \DFF_99.D ;
  assign g17226 = \DFF_104.D ;
  assign g17227 = \DFF_16.D ;
  assign g17228 = \DFF_102.D ;
  assign g17229 = \DFF_119.D ;
  assign g1723 = \DFF_1029.Q ;
  assign g17233 = \DFF_15.D ;
  assign g17234 = \DFF_100.D ;
  assign g17235 = \DFF_105.D ;
  assign g17236 = \DFF_122.D ;
  assign g1724 = \DFF_954.Q ;
  assign g17246 = \DFF_103.D ;
  assign g17247 = \DFF_120.D ;
  assign g17248 = \DFF_125.D ;
  assign g17269 = \DFF_106.D ;
  assign g1727 = \DFF_955.Q ;
  assign g17270 = \DFF_123.D ;
  assign g17271 = \DFF_128.D ;
  assign g173 = \DFF_198.Q ;
  assign g1730 = \DFF_1030.Q ;
  assign g17300 = g51;
  assign g17302 = \DFF_121.D ;
  assign g17303 = \DFF_126.D ;
  assign g1731 = \DFF_1031.Q ;
  assign g1732 = \DFF_1032.Q ;
  assign g1733 = \DFF_1033.Q ;
  assign g1734 = \DFF_1034.Q ;
  assign g17340 = \DFF_124.D ;
  assign g17341 = \DFF_129.D ;
  assign g1735 = \DFF_953.Q ;
  assign g1738 = \DFF_1035.Q ;
  assign g17383 = \DFF_127.D ;
  assign g1739 = \DFF_957.Q ;
  assign g174 = \DFF_202.Q ;
  assign g1742 = \DFF_958.Q ;
  assign g17429 = \DFF_130.D ;
  assign g17442 = \DFF_316.D ;
  assign g1745 = \DFF_1036.Q ;
  assign g1746 = \DFF_1037.Q ;
  assign g1747 = \DFF_1038.Q ;
  assign g1748 = \DFF_1039.Q ;
  assign g1749 = \DFF_1040.Q ;
  assign g175 = \DFF_200.Q ;
  assign g1750 = \DFF_956.Q ;
  assign g17500 = \DFF_316.D ;
  assign g17503 = \DFF_316.D ;
  assign g17523 = \DFF_666.D ;
  assign g1753 = \DFF_1041.Q ;
  assign g1754 = \DFF_960.Q ;
  assign g1757 = \DFF_961.Q ;
  assign g17570 = \DFF_316.D ;
  assign g17591 = \DFF_666.D ;
  assign g17594 = \DFF_666.D ;
  assign g176 = \DFF_201.Q ;
  assign g1760 = \DFF_1042.Q ;
  assign g1761 = \DFF_1043.Q ;
  assign g17613 = \DFF_1016.D ;
  assign g1762 = \DFF_1044.Q ;
  assign g1763 = \DFF_1045.Q ;
  assign g1764 = \DFF_1046.Q ;
  assign g17645 = \DFF_1296.D ;
  assign g1765 = \DFF_959.Q ;
  assign g17667 = \DFF_666.D ;
  assign g1768 = \DFF_1047.Q ;
  assign g17688 = \DFF_1016.D ;
  assign g1769 = \DFF_963.Q ;
  assign g17691 = \DFF_1016.D ;
  assign g177 = \DFF_205.Q ;
  assign g17710 = \DFF_1366.D ;
  assign g1772 = \DFF_964.Q ;
  assign g17746 = \DFF_1296.D ;
  assign g1775 = \DFF_1048.Q ;
  assign g1776 = \DFF_1049.Q ;
  assign g17767 = \DFF_1016.D ;
  assign g1777 = \DFF_1050.Q ;
  assign g1778 = \DFF_1051.Q ;
  assign g17788 = \DFF_1366.D ;
  assign g1779 = \DFF_962.Q ;
  assign g17791 = \DFF_1366.D ;
  assign g178 = \DFF_203.Q ;
  assign g1782 = \DFF_1429.Q ;
  assign g1783 = \DFF_997.Q ;
  assign g1784 = \DFF_995.Q ;
  assign g17847 = \DFF_1296.D ;
  assign g1785 = \DFF_996.Q ;
  assign g1786 = \DFF_1428.Q ;
  assign g17868 = \DFF_1366.D ;
  assign g1789 = \DFF_965.Q ;
  assign g179 = \DFF_204.Q ;
  assign g1792 = \DFF_966.Q ;
  assign g1795 = \DFF_967.Q ;
  assign g17959 = \DFF_1296.D ;
  assign g1798 = \DFF_968.Q ;
  assign g180 = \DFF_1296.Q ;
  assign g1801 = \DFF_969.Q ;
  assign g1804 = \DFF_970.Q ;
  assign g1807 = \DFF_973.Q ;
  assign g1808 = \DFF_971.Q ;
  assign g1809 = \DFF_972.Q ;
  assign g181 = \DFF_1302.Q ;
  assign g1810 = \DFF_974.Q ;
  assign g1813 = \DFF_975.Q ;
  assign g1816 = \DFF_976.Q ;
  assign g1819 = \DFF_977.Q ;
  assign g182 = \DFF_1297.Q ;
  assign g1822 = \DFF_978.Q ;
  assign g1825 = \DFF_979.Q ;
  assign g1828 = \DFF_982.Q ;
  assign g1829 = \DFF_980.Q ;
  assign g1830 = \DFF_981.Q ;
  assign g1831 = \DFF_998.Q ;
  assign g1832 = \DFF_999.Q ;
  assign g1833 = \DFF_1000.Q ;
  assign g1834 = \DFF_1001.Q ;
  assign g1835 = \DFF_1002.Q ;
  assign g1836 = \DFF_1083.Q ;
  assign g1839 = \DFF_1084.Q ;
  assign g1842 = \DFF_1085.Q ;
  assign g1845 = \DFF_1091.Q ;
  assign g1846 = \DFF_1092.Q ;
  assign g1849 = \DFF_1093.Q ;
  assign g185 = \DFF_160.Q ;
  assign g1852 = \DFF_1094.Q ;
  assign g18542 = \DFF_1635.D ;
  assign g1855 = \DFF_1427.Q ;
  assign g1858 = \DFF_1086.Q ;
  assign g1859 = \DFF_1087.Q ;
  assign g186 = \DFF_206.Q ;
  assign g1860 = \DFF_1088.Q ;
  assign g1861 = \DFF_1089.Q ;
  assign g1862 = \DFF_1428.Q ;
  assign g1865 = \DFF_1090.Q ;
  assign g1866 = \DFF_1429.Q ;
  assign g18669 = \DFF_95.D ;
  assign g1867 = \DFF_1080.Q ;
  assign g18678 = \DFF_360.D ;
  assign g1868 = \DFF_1081.Q ;
  assign g1869 = \DFF_1082.Q ;
  assign g1870 = \DFF_1076.Q ;
  assign g18707 = \DFF_710.D ;
  assign g1871 = \DFF_1129.Q ;
  assign g18719 = \DFF_96.D ;
  assign g18726 = \DFF_361.D ;
  assign g1874 = \DFF_1130.Q ;
  assign g18743 = \DFF_1060.D ;
  assign g18754 = \DFF_38.D ;
  assign g18755 = \DFF_1629.D ;
  assign g18763 = \DFF_711.D ;
  assign g1877 = \DFF_1131.Q ;
  assign g18780 = \DFF_1410.D ;
  assign g18781 = \DFF_39.D ;
  assign g18782 = \DFF_97.D ;
  assign g18794 = \DFF_1061.D ;
  assign g1880 = \DFF_1102.Q ;
  assign g18803 = \DFF_40.D ;
  assign g18804 = \DFF_1630.D ;
  assign g18820 = \DFF_1411.D ;
  assign g18821 = \DFF_41.D ;
  assign g18835 = \DFF_42.D ;
  assign g18836 = \DFF_89.D ;
  assign g18837 = \DFF_1631.D ;
  assign g18852 = \DFF_43.D ;
  assign g1886 = \DFF_1132.Q ;
  assign g18866 = \DFF_44.D ;
  assign g18867 = \DFF_88.D ;
  assign g18868 = \DFF_1632.D ;
  assign g1887 = \DFF_1133.Q ;
  assign g18883 = \DFF_45.D ;
  assign g18885 = \DFF_83.D ;
  assign g189 = \DFF_207.Q ;
  assign g1890 = \DFF_1061.Q ;
  assign g18906 = \DFF_87.D ;
  assign g18907 = \DFF_1633.D ;
  assign g1893 = \DFF_1062.Q ;
  assign g18942 = \DFF_86.D ;
  assign g18957 = \DFF_90.D ;
  assign g18968 = \DFF_85.D ;
  assign g18975 = \DFF_84.D ;
  assign g1900 = \DFF_1142.Q ;
  assign g19000 = \DFF_316.D ;
  assign g19012 = \DFF_316.D ;
  assign g19021 = \DFF_398.D ;
  assign g19022 = \DFF_401.D ;
  assign g19023 = \DFF_403.D ;
  assign g19024 = \DFF_666.D ;
  assign g1903 = \DFF_1063.Q ;
  assign g19033 = \DFF_748.D ;
  assign g19034 = \DFF_751.D ;
  assign g19035 = \DFF_753.D ;
  assign g19036 = \DFF_1016.D ;
  assign g1904 = \DFF_1064.Q ;
  assign g19045 = \DFF_1098.D ;
  assign g19046 = \DFF_1101.D ;
  assign g19047 = \DFF_1103.D ;
  assign g19048 = \DFF_1366.D ;
  assign g1905 = \DFF_1143.Q ;
  assign g19057 = \DFF_1448.D ;
  assign g19058 = \DFF_1451.D ;
  assign g19059 = \DFF_1453.D ;
  assign g19060 = \DFF_16.D ;
  assign g19061 = \DFF_15.D ;
  assign g19062 = g51;
  assign g1908 = \DFF_1095.Q ;
  assign g1909 = \DFF_1144.Q ;
  assign g19096 = \DFF_1624.D ;
  assign g1910 = \DFF_1145.Q ;
  assign g1911 = \DFF_1146.Q ;
  assign g1912 = \DFF_1147.Q ;
  assign g1913 = \DFF_1148.Q ;
  assign g1914 = \DFF_1149.Q ;
  assign g19144 = \DFF_71.D ;
  assign g19145 = \DFF_1296.D ;
  assign g19147 = \DFF_1296.D ;
  assign g19149 = \DFF_73.D ;
  assign g1915 = \DFF_1096.Q ;
  assign g19151 = \DFF_1296.D ;
  assign g19152 = \DFF_3.D ;
  assign g19153 = \DFF_65.D ;
  assign g19154 = \DFF_47.D ;
  assign g19156 = \DFF_1296.D ;
  assign g19157 = \DFF_75.D ;
  assign g19158 = \DFF_95.D ;
  assign g19159 = \DFF_360.D ;
  assign g1916 = \DFF_1150.Q ;
  assign g19162 = \DFF_67.D ;
  assign g19163 = \DFF_49.D ;
  assign g19164 = \DFF_710.D ;
  assign g19167 = \DFF_77.D ;
  assign g19168 = \DFF_96.D ;
  assign g19169 = \DFF_361.D ;
  assign g1917 = \DFF_1151.Q ;
  assign g19170 = \DFF_1060.D ;
  assign g19172 = \DFF_69.D ;
  assign g19173 = \DFF_51.D ;
  assign g19174 = \DFF_1629.D ;
  assign g19175 = \DFF_711.D ;
  assign g19176 = \DFF_1410.D ;
  assign g19178 = \DFF_79.D ;
  assign g1918 = \DFF_1152.Q ;
  assign g19180 = \DFF_97.D ;
  assign g19182 = \DFF_1061.D ;
  assign g19183 = \DFF_41.D ;
  assign g19184 = \DFF_53.D ;
  assign g19185 = \DFF_1630.D ;
  assign g19189 = \DFF_1411.D ;
  assign g19190 = \DFF_42.D ;
  assign g19196 = \DFF_43.D ;
  assign g19197 = \DFF_89.D ;
  assign g19198 = \DFF_84.D ;
  assign g19199 = \DFF_1631.D ;
  assign g192 = \DFF_208.Q ;
  assign g19207 = \DFF_44.D ;
  assign g19208 = \DFF_85.D ;
  assign g1921 = \DFF_1153.Q ;
  assign g19217 = \DFF_45.D ;
  assign g19218 = \DFF_88.D ;
  assign g1922 = \DFF_1097.Q ;
  assign g19220 = \DFF_1632.D ;
  assign g19229 = \DFF_83.D ;
  assign g1923 = \DFF_1098.Q ;
  assign g19237 = \DFF_38.D ;
  assign g19238 = \DFF_87.D ;
  assign g19239 = \DFF_1633.D ;
  assign g1924 = \DFF_1099.Q ;
  assign g19247 = \DFF_39.D ;
  assign g19249 = \DFF_1635.D ;
  assign g1925 = \DFF_1504.Q ;
  assign g19258 = \DFF_40.D ;
  assign g19259 = \DFF_86.D ;
  assign g19270 = \DFF_90.D ;
  assign g1928 = \DFF_1100.Q ;
  assign g1929 = \DFF_1101.Q ;
  assign g1930 = \DFF_1506.Q ;
  assign g1931 = \DFF_1505.Q ;
  assign g1934 = \DFF_1059.Q ;
  assign g1937 = \DFF_1060.Q ;
  assign g1938 = \DFF_1103.Q ;
  assign g1939 = \DFF_1104.Q ;
  assign g1942 = g1943;
  assign g1944 = \DFF_1065.Q ;
  assign g1945 = \DFF_1072.Q ;
  assign g1946 = \DFF_1073.Q ;
  assign g1947 = \DFF_1074.Q ;
  assign g1948 = \DFF_1075.Q ;
  assign g19484 = g3229;
  assign g1949 = \DFF_1066.Q ;
  assign g195 = \DFF_212.Q ;
  assign g1950 = \DFF_1067.Q ;
  assign g19505 = g3229;
  assign g1951 = \DFF_1068.Q ;
  assign g1952 = \DFF_1069.Q ;
  assign g19524 = g3229;
  assign g1953 = \DFF_1070.Q ;
  assign g19534 = g3229;
  assign g1954 = \DFF_1071.Q ;
  assign g19543 = \DFF_457.D ;
  assign g19546 = \DFF_807.D ;
  assign g1955 = \DFF_1107.Q ;
  assign g19550 = \DFF_1157.D ;
  assign g19556 = \DFF_1507.D ;
  assign g1956 = \DFF_1105.Q ;
  assign g19563 = \DFF_1617.D ;
  assign g1957 = \DFF_1106.Q ;
  assign g19573 = \DFF_1622.D ;
  assign g19578 = g3229;
  assign g1958 = \DFF_1110.Q ;
  assign g1959 = \DFF_1108.Q ;
  assign g19595 = \DFF_1618.D ;
  assign g19596 = \DFF_1623.D ;
  assign g1960 = \DFF_1109.Q ;
  assign g19608 = g3229;
  assign g1961 = \DFF_1113.Q ;
  assign g1962 = \DFF_1111.Q ;
  assign g19622 = \DFF_1614.D ;
  assign g1963 = \DFF_1112.Q ;
  assign g1964 = \DFF_1116.Q ;
  assign g19641 = g3229;
  assign g1965 = \DFF_1114.Q ;
  assign g19652 = \DFF_1619.D ;
  assign g1966 = \DFF_1115.Q ;
  assign g1967 = \DFF_1117.Q ;
  assign g19681 = g3229;
  assign g19689 = \DFF_1615.D ;
  assign g19690 = \DFF_1625.D ;
  assign g19696 = \DFF_316.D ;
  assign g1970 = \DFF_1118.Q ;
  assign g19725 = \DFF_1620.D ;
  assign g1973 = \DFF_1119.Q ;
  assign g19740 = \DFF_666.D ;
  assign g1976 = \DFF_1120.Q ;
  assign g19762 = \DFF_1616.D ;
  assign g19763 = \DFF_1626.D ;
  assign g19783 = \DFF_1016.D ;
  assign g1979 = \DFF_1121.Q ;
  assign g19798 = \DFF_1621.D ;
  assign g198 = \DFF_213.Q ;
  assign g1982 = \DFF_1122.Q ;
  assign g19825 = \DFF_1366.D ;
  assign g19830 = g3234;
  assign g19838 = \DFF_1627.D ;
  assign g1985 = \DFF_1126.Q ;
  assign g1988 = \DFF_1127.Q ;
  assign g19893 = \DFF_1628.D ;
  assign g1991 = \DFF_1128.Q ;
  assign g1994 = \DFF_1123.Q ;
  assign g1997 = \DFF_1124.Q ;
  assign g2 = \DFF_1632.Q ;
  assign g20 = \DFF_1626.Q ;
  assign g2000 = \DFF_1125.Q ;
  assign g2003 = \DFF_1504.Q ;
  assign g2006 = \DFF_1505.Q ;
  assign g20082 = \DFF_1.D ;
  assign g20083 = \DFF_1634.D ;
  assign g2009 = \DFF_1506.Q ;
  assign g201 = \DFF_214.Q ;
  assign g2010 = \DFF_1157.Q ;
  assign g20105 = \DFF_2.D ;
  assign g2013 = \DFF_1160.Q ;
  assign g20164 = \DFF_1296.D ;
  assign g20193 = \DFF_316.D ;
  assign g20198 = \DFF_1296.D ;
  assign g2020 = \DFF_1159.Q ;
  assign g20223 = \DFF_666.D ;
  assign g20228 = \DFF_1296.D ;
  assign g20250 = \DFF_1016.D ;
  assign g20255 = \DFF_1296.D ;
  assign g2026 = \DFF_1162.Q ;
  assign g20273 = \DFF_1366.D ;
  assign g20310 = \DFF_55.D ;
  assign g20314 = \DFF_458.D ;
  assign g2033 = \DFF_1161.Q ;
  assign g20333 = \DFF_808.D ;
  assign g20343 = \DFF_57.D ;
  assign g20353 = \DFF_1158.D ;
  assign g20360 = \DFF_98.D ;
  assign g20375 = \DFF_1508.D ;
  assign g20376 = \DFF_59.D ;
  assign g20377 = \DFF_101.D ;
  assign g2039 = \DFF_1158.Q ;
  assign g20395 = \DFF_99.D ;
  assign g20396 = \DFF_104.D ;
  assign g204 = \DFF_218.Q ;
  assign g2040 = \DFF_1163.Q ;
  assign g20417 = \DFF_61.D ;
  assign g20418 = \DFF_102.D ;
  assign g20419 = \DFF_119.D ;
  assign g20439 = \DFF_100.D ;
  assign g20440 = \DFF_105.D ;
  assign g20441 = \DFF_122.D ;
  assign g20457 = \DFF_103.D ;
  assign g20458 = \DFF_120.D ;
  assign g20459 = \DFF_125.D ;
  assign g2046 = \DFF_1165.Q ;
  assign g20469 = \DFF_106.D ;
  assign g20470 = \DFF_123.D ;
  assign g20471 = \DFF_128.D ;
  assign g20478 = \DFF_121.D ;
  assign g20479 = \DFF_126.D ;
  assign g20484 = \DFF_124.D ;
  assign g20485 = \DFF_129.D ;
  assign g20491 = \DFF_127.D ;
  assign g20497 = \DFF_1563.D ;
  assign g20498 = \DFF_130.D ;
  assign g2052 = \DFF_1164.Q ;
  assign g20555 = \DFF_1296.D ;
  assign g20556 = \DFF_360.D ;
  assign g20557 = \DFF_361.D ;
  assign g20558 = \DFF_457.D ;
  assign g20559 = \DFF_1296.D ;
  assign g20560 = \DFF_710.D ;
  assign g20561 = \DFF_711.D ;
  assign g20562 = \DFF_807.D ;
  assign g20563 = \DFF_1296.D ;
  assign g20564 = \DFF_1060.D ;
  assign g20565 = \DFF_1061.D ;
  assign g20566 = \DFF_1157.D ;
  assign g20567 = \DFF_1296.D ;
  assign g20568 = \DFF_1410.D ;
  assign g20569 = \DFF_1411.D ;
  assign g20570 = \DFF_1507.D ;
  assign g20571 = \DFF_1.D ;
  assign g20572 = \DFF_38.D ;
  assign g20573 = \DFF_39.D ;
  assign g20574 = \DFF_40.D ;
  assign g20575 = \DFF_41.D ;
  assign g20576 = \DFF_42.D ;
  assign g20577 = \DFF_43.D ;
  assign g20578 = \DFF_44.D ;
  assign g20579 = \DFF_45.D ;
  assign g20580 = \DFF_90.D ;
  assign g20581 = \DFF_89.D ;
  assign g20582 = \DFF_88.D ;
  assign g20583 = \DFF_87.D ;
  assign g20584 = \DFF_86.D ;
  assign g20585 = \DFF_84.D ;
  assign g20586 = \DFF_85.D ;
  assign g20587 = \DFF_83.D ;
  assign g20588 = \DFF_2.D ;
  assign g20589 = \DFF_1629.D ;
  assign g2059 = \DFF_1166.Q ;
  assign g20590 = \DFF_1630.D ;
  assign g20591 = \DFF_1631.D ;
  assign g20592 = \DFF_1632.D ;
  assign g20593 = \DFF_1633.D ;
  assign g20594 = \DFF_1635.D ;
  assign g20595 = \DFF_1614.D ;
  assign g20596 = \DFF_1615.D ;
  assign g20597 = \DFF_1616.D ;
  assign g20598 = \DFF_1617.D ;
  assign g20599 = \DFF_1618.D ;
  assign g20600 = \DFF_1619.D ;
  assign g20601 = \DFF_1620.D ;
  assign g20602 = \DFF_1621.D ;
  assign g20603 = \DFF_1622.D ;
  assign g20604 = \DFF_1623.D ;
  assign g20605 = \DFF_1625.D ;
  assign g20606 = \DFF_1626.D ;
  assign g20607 = \DFF_1627.D ;
  assign g20608 = \DFF_1628.D ;
  assign g20609 = \DFF_98.D ;
  assign g20610 = \DFF_99.D ;
  assign g20611 = \DFF_100.D ;
  assign g20612 = \DFF_101.D ;
  assign g20613 = \DFF_102.D ;
  assign g20614 = \DFF_103.D ;
  assign g20615 = \DFF_104.D ;
  assign g20616 = \DFF_105.D ;
  assign g20617 = \DFF_106.D ;
  assign g20618 = \DFF_119.D ;
  assign g20619 = \DFF_120.D ;
  assign g20620 = \DFF_121.D ;
  assign g20621 = \DFF_122.D ;
  assign g20622 = \DFF_123.D ;
  assign g20623 = \DFF_124.D ;
  assign g20624 = \DFF_125.D ;
  assign g20625 = \DFF_126.D ;
  assign g20626 = \DFF_127.D ;
  assign g20627 = \DFF_128.D ;
  assign g20628 = \DFF_129.D ;
  assign g20629 = \DFF_130.D ;
  assign g20630 = \DFF_95.D ;
  assign g20631 = \DFF_96.D ;
  assign g20632 = \DFF_97.D ;
  assign g2066 = \DFF_1167.Q ;
  assign g20682 = \DFF_459.D ;
  assign g207 = \DFF_219.Q ;
  assign g20717 = \DFF_809.D ;
  assign g2072 = \DFF_1168.Q ;
  assign g20752 = \DFF_1159.D ;
  assign g2078 = \DFF_1171.Q ;
  assign g20789 = \DFF_1509.D ;
  assign g2079 = \DFF_1169.Q ;
  assign g2080 = \DFF_1170.Q ;
  assign g2081 = \DFF_1174.Q ;
  assign g2082 = \DFF_1172.Q ;
  assign g20825 = \DFF_4.D ;
  assign g2083 = \DFF_1173.Q ;
  assign g2084 = \DFF_1177.Q ;
  assign g2085 = \DFF_1175.Q ;
  assign g2086 = \DFF_1176.Q ;
  assign g2087 = \DFF_1180.Q ;
  assign g20874 = \DFF_81.D ;
  assign g20875 = \DFF_469.D ;
  assign g20876 = \DFF_496.D ;
  assign g20877 = \DFF_1561.D ;
  assign g20879 = \DFF_470.D ;
  assign g2088 = \DFF_1178.Q ;
  assign g20880 = \DFF_472.D ;
  assign g20881 = \DFF_497.D ;
  assign g20882 = \DFF_819.D ;
  assign g20883 = \DFF_846.D ;
  assign g20884 = \DFF_1562.D ;
  assign g2089 = \DFF_1179.Q ;
  assign g20891 = \DFF_471.D ;
  assign g20892 = \DFF_473.D ;
  assign g20893 = \DFF_475.D ;
  assign g20894 = \DFF_498.D ;
  assign g20896 = \DFF_820.D ;
  assign g20897 = \DFF_822.D ;
  assign g20898 = \DFF_847.D ;
  assign g20899 = \DFF_1169.D ;
  assign g2090 = \DFF_1183.Q ;
  assign g20900 = \DFF_1196.D ;
  assign g20901 = \DFF_474.D ;
  assign g20902 = \DFF_476.D ;
  assign g20903 = \DFF_478.D ;
  assign g2091 = \DFF_1181.Q ;
  assign g20910 = \DFF_821.D ;
  assign g20911 = \DFF_823.D ;
  assign g20912 = \DFF_825.D ;
  assign g20913 = \DFF_848.D ;
  assign g20915 = \DFF_1170.D ;
  assign g20916 = \DFF_1172.D ;
  assign g20917 = \DFF_1197.D ;
  assign g20918 = \DFF_1519.D ;
  assign g20919 = \DFF_1546.D ;
  assign g2092 = \DFF_1182.Q ;
  assign g20921 = \DFF_477.D ;
  assign g20922 = \DFF_479.D ;
  assign g20923 = \DFF_481.D ;
  assign g20924 = \DFF_499.D ;
  assign g20925 = \DFF_824.D ;
  assign g20926 = \DFF_826.D ;
  assign g20927 = \DFF_828.D ;
  assign g2093 = \DFF_1186.Q ;
  assign g20934 = \DFF_1171.D ;
  assign g20935 = \DFF_1173.D ;
  assign g20936 = \DFF_1175.D ;
  assign g20937 = \DFF_1198.D ;
  assign g20939 = \DFF_1520.D ;
  assign g2094 = \DFF_1184.Q ;
  assign g20940 = \DFF_1522.D ;
  assign g20941 = \DFF_1547.D ;
  assign g20942 = \DFF_55.D ;
  assign g20943 = \DFF_458.D ;
  assign g20944 = \DFF_480.D ;
  assign g20945 = \DFF_482.D ;
  assign g20946 = \DFF_484.D ;
  assign g20947 = \DFF_500.D ;
  assign g20948 = \DFF_502.D ;
  assign g20949 = \DFF_827.D ;
  assign g2095 = \DFF_1185.Q ;
  assign g20950 = \DFF_829.D ;
  assign g20951 = \DFF_831.D ;
  assign g20952 = \DFF_849.D ;
  assign g20953 = \DFF_1174.D ;
  assign g20954 = \DFF_1176.D ;
  assign g20955 = \DFF_1178.D ;
  assign g2096 = \DFF_1189.Q ;
  assign g20962 = \DFF_1521.D ;
  assign g20963 = \DFF_1523.D ;
  assign g20964 = \DFF_1525.D ;
  assign g20965 = \DFF_1548.D ;
  assign g20966 = \DFF_483.D ;
  assign g20967 = \DFF_485.D ;
  assign g20968 = \DFF_487.D ;
  assign g20969 = \DFF_501.D ;
  assign g2097 = \DFF_1187.Q ;
  assign g20970 = \DFF_503.D ;
  assign g20971 = \DFF_808.D ;
  assign g20972 = \DFF_830.D ;
  assign g20973 = \DFF_832.D ;
  assign g20974 = \DFF_834.D ;
  assign g20975 = \DFF_850.D ;
  assign g20976 = \DFF_852.D ;
  assign g20977 = \DFF_1177.D ;
  assign g20978 = \DFF_1179.D ;
  assign g20979 = \DFF_1181.D ;
  assign g2098 = \DFF_1188.Q ;
  assign g20980 = \DFF_1199.D ;
  assign g20981 = \DFF_1524.D ;
  assign g20982 = \DFF_1526.D ;
  assign g20983 = \DFF_1528.D ;
  assign g20984 = \DFF_57.D ;
  assign g20985 = \DFF_1634.D ;
  assign g20989 = \DFF_486.D ;
  assign g2099 = \DFF_1192.Q ;
  assign g20990 = \DFF_488.D ;
  assign g20991 = \DFF_490.D ;
  assign g20992 = \DFF_504.D ;
  assign g20993 = \DFF_833.D ;
  assign g20994 = \DFF_835.D ;
  assign g20995 = \DFF_837.D ;
  assign g20996 = \DFF_851.D ;
  assign g20997 = \DFF_853.D ;
  assign g20998 = \DFF_1158.D ;
  assign g20999 = \DFF_1180.D ;
  assign g210 = \DFF_220.Q ;
  assign g2100 = \DFF_1190.Q ;
  assign g21000 = \DFF_1182.D ;
  assign g21001 = \DFF_1184.D ;
  assign g21002 = \DFF_1200.D ;
  assign g21003 = \DFF_1202.D ;
  assign g21004 = \DFF_1527.D ;
  assign g21005 = \DFF_1529.D ;
  assign g21006 = \DFF_1531.D ;
  assign g21007 = \DFF_1549.D ;
  assign g21009 = \DFF_489.D ;
  assign g2101 = \DFF_1191.Q ;
  assign g21010 = \DFF_491.D ;
  assign g21011 = \DFF_493.D ;
  assign g21015 = \DFF_836.D ;
  assign g21016 = \DFF_838.D ;
  assign g21017 = \DFF_840.D ;
  assign g21018 = \DFF_854.D ;
  assign g21019 = \DFF_1183.D ;
  assign g2102 = \DFF_1195.Q ;
  assign g21020 = \DFF_1185.D ;
  assign g21021 = \DFF_1187.D ;
  assign g21022 = \DFF_1201.D ;
  assign g21023 = \DFF_1203.D ;
  assign g21024 = \DFF_1508.D ;
  assign g21025 = \DFF_1530.D ;
  assign g21026 = \DFF_1532.D ;
  assign g21027 = \DFF_1534.D ;
  assign g21028 = \DFF_1550.D ;
  assign g21029 = \DFF_1552.D ;
  assign g2103 = \DFF_1193.Q ;
  assign g21030 = \DFF_59.D ;
  assign g21031 = \DFF_492.D ;
  assign g21032 = \DFF_494.D ;
  assign g21033 = \DFF_839.D ;
  assign g21034 = \DFF_841.D ;
  assign g21035 = \DFF_843.D ;
  assign g21039 = \DFF_1186.D ;
  assign g2104 = \DFF_1194.Q ;
  assign g21040 = \DFF_1188.D ;
  assign g21041 = \DFF_1190.D ;
  assign g21042 = \DFF_1204.D ;
  assign g21043 = \DFF_1533.D ;
  assign g21044 = \DFF_1535.D ;
  assign g21045 = \DFF_1537.D ;
  assign g21046 = \DFF_1551.D ;
  assign g21047 = \DFF_1553.D ;
  assign g2105 = \DFF_1198.Q ;
  assign g21050 = g3229;
  assign g21051 = \DFF_495.D ;
  assign g21052 = \DFF_842.D ;
  assign g21053 = \DFF_844.D ;
  assign g21054 = \DFF_1189.D ;
  assign g21055 = \DFF_1191.D ;
  assign g21056 = \DFF_1193.D ;
  assign g2106 = \DFF_1196.Q ;
  assign g21060 = \DFF_1536.D ;
  assign g21061 = \DFF_1538.D ;
  assign g21062 = \DFF_1540.D ;
  assign g21063 = \DFF_1554.D ;
  assign g21064 = \DFF_61.D ;
  assign g21069 = g3229;
  assign g2107 = \DFF_1197.Q ;
  assign g21070 = \DFF_845.D ;
  assign g21071 = \DFF_1192.D ;
  assign g21072 = \DFF_1194.D ;
  assign g21073 = \DFF_1539.D ;
  assign g21074 = \DFF_1541.D ;
  assign g21075 = \DFF_1543.D ;
  assign g21079 = g3229;
  assign g2108 = \DFF_1201.Q ;
  assign g21080 = \DFF_1195.D ;
  assign g21081 = \DFF_1542.D ;
  assign g21082 = \DFF_1544.D ;
  assign g2109 = \DFF_1199.Q ;
  assign g21093 = g3229;
  assign g21094 = \DFF_1545.D ;
  assign g2110 = \DFF_1200.Q ;
  assign g2111 = \DFF_1204.Q ;
  assign g2112 = \DFF_1202.Q ;
  assign g2113 = \DFF_1203.Q ;
  assign g2114 = \DFF_1207.Q ;
  assign g2115 = \DFF_1205.Q ;
  assign g2116 = \DFF_1206.Q ;
  assign g2117 = \DFF_1210.Q ;
  assign g2118 = \DFF_1208.Q ;
  assign g21187 = g3229;
  assign g2119 = \DFF_1209.Q ;
  assign g2120 = \DFF_1295.Q ;
  assign g21202 = g3229;
  assign g21217 = g3229;
  assign g21225 = g3229;
  assign g2124 = \DFF_1294.Q ;
  assign g2129 = \DFF_1293.Q ;
  assign g213 = \DFF_224.Q ;
  assign g21327 = \DFF_71.D ;
  assign g2133 = \DFF_1292.Q ;
  assign g21346 = \DFF_317.D ;
  assign g21358 = \DFF_73.D ;
  assign g21359 = \DFF_1624.D ;
  assign g21376 = \DFF_65.D ;
  assign g21377 = \DFF_47.D ;
  assign g2138 = \DFF_1291.Q ;
  assign g21399 = \DFF_75.D ;
  assign g2142 = \DFF_1290.Q ;
  assign g21426 = \DFF_67.D ;
  assign g21427 = \DFF_49.D ;
  assign g21435 = \DFF_442.D ;
  assign g21457 = \DFF_77.D ;
  assign g2147 = \DFF_1289.Q ;
  assign g21495 = \DFF_69.D ;
  assign g21496 = \DFF_51.D ;
  assign g2151 = \DFF_1288.Q ;
  assign g21528 = \DFF_79.D ;
  assign g21557 = \DFF_53.D ;
  assign g2156 = \DFF_1287.Q ;
  assign g216 = \DFF_225.Q ;
  assign g2160 = \DFF_1286.Q ;
  assign g2165 = \DFF_90.Q ;
  assign g2170 = \DFF_89.Q ;
  assign g2175 = \DFF_88.Q ;
  assign g21795 = \DFF_3.D ;
  assign g2180 = \DFF_87.Q ;
  assign g21824 = \DFF_1563.D ;
  assign g21842 = \DFF_359.D ;
  assign g21843 = \DFF_709.D ;
  assign g21845 = \DFF_1059.D ;
  assign g21847 = \DFF_1409.D ;
  assign g2185 = \DFF_86.Q ;
  assign g21851 = \DFF_400.D ;
  assign g21878 = \DFF_63.D ;
  assign g21880 = \DFF_46.D ;
  assign g21882 = \DFF_91.D ;
  assign g219 = \DFF_226.Q ;
  assign g2190 = \DFF_85.Q ;
  assign g21943 = \DFF_458.D ;
  assign g21944 = \DFF_808.D ;
  assign g21945 = \DFF_1158.D ;
  assign g21946 = \DFF_1508.D ;
  assign g21947 = \DFF_55.D ;
  assign g21948 = \DFF_57.D ;
  assign g21949 = \DFF_59.D ;
  assign g2195 = \DFF_84.Q ;
  assign g21950 = \DFF_61.D ;
  assign g21951 = \DFF_3.D ;
  assign g21952 = \DFF_65.D ;
  assign g21953 = \DFF_67.D ;
  assign g21954 = \DFF_69.D ;
  assign g21955 = \DFF_71.D ;
  assign g21956 = \DFF_73.D ;
  assign g21957 = \DFF_75.D ;
  assign g21958 = \DFF_77.D ;
  assign g21959 = \DFF_79.D ;
  assign g21960 = \DFF_47.D ;
  assign g21961 = \DFF_49.D ;
  assign g21962 = \DFF_51.D ;
  assign g21963 = \DFF_53.D ;
  assign g21964 = \DFF_1634.D ;
  assign g21965 = \DFF_1563.D ;
  assign g21966 = \DFF_1624.D ;
  assign g21969 = \DFF_810.D ;
  assign g21970 = \DFF_1432.D ;
  assign g21972 = \DFF_1160.D ;
  assign g21974 = \DFF_1510.D ;
  assign g21989 = \DFF_11.D ;
  assign g2200 = \DFF_83.Q ;
  assign g22002 = \DFF_1607.D ;
  assign g22025 = \DFF_170.D ;
  assign g22026 = \DFF_5.D ;
  assign g22027 = \DFF_171.D ;
  assign g22028 = \DFF_173.D ;
  assign g22029 = \DFF_520.D ;
  assign g22030 = \DFF_172.D ;
  assign g22031 = \DFF_174.D ;
  assign g22032 = \DFF_176.D ;
  assign g22033 = \DFF_521.D ;
  assign g22034 = \DFF_523.D ;
  assign g22035 = \DFF_870.D ;
  assign g22037 = \DFF_175.D ;
  assign g22038 = \DFF_177.D ;
  assign g22039 = \DFF_179.D ;
  assign g22040 = \DFF_522.D ;
  assign g22041 = \DFF_524.D ;
  assign g22042 = \DFF_526.D ;
  assign g22043 = \DFF_871.D ;
  assign g22044 = \DFF_873.D ;
  assign g22045 = \DFF_1220.D ;
  assign g22047 = \DFF_178.D ;
  assign g22048 = \DFF_180.D ;
  assign g22049 = \DFF_182.D ;
  assign g2205 = \DFF_1216.Q ;
  assign g22054 = \DFF_525.D ;
  assign g22055 = \DFF_527.D ;
  assign g22056 = \DFF_529.D ;
  assign g22057 = \DFF_872.D ;
  assign g22058 = \DFF_874.D ;
  assign g22059 = \DFF_876.D ;
  assign g2206 = \DFF_1214.Q ;
  assign g22060 = \DFF_1221.D ;
  assign g22061 = \DFF_1223.D ;
  assign g22063 = \DFF_181.D ;
  assign g22064 = \DFF_183.D ;
  assign g22065 = \DFF_185.D ;
  assign g22066 = \DFF_528.D ;
  assign g22067 = \DFF_530.D ;
  assign g22068 = \DFF_532.D ;
  assign g2207 = \DFF_1215.Q ;
  assign g22073 = \DFF_875.D ;
  assign g22074 = \DFF_877.D ;
  assign g22075 = \DFF_879.D ;
  assign g22076 = \DFF_1222.D ;
  assign g22077 = \DFF_1224.D ;
  assign g22078 = \DFF_1226.D ;
  assign g22079 = \DFF_184.D ;
  assign g2208 = \DFF_1219.Q ;
  assign g22080 = \DFF_186.D ;
  assign g22081 = \DFF_188.D ;
  assign g22082 = \DFF_359.D ;
  assign g22087 = \DFF_531.D ;
  assign g22088 = \DFF_533.D ;
  assign g22089 = \DFF_535.D ;
  assign g2209 = \DFF_1217.Q ;
  assign g22090 = \DFF_878.D ;
  assign g22091 = \DFF_880.D ;
  assign g22092 = \DFF_882.D ;
  assign g22097 = \DFF_1225.D ;
  assign g22098 = \DFF_1227.D ;
  assign g22099 = \DFF_1229.D ;
  assign g2210 = \DFF_1218.Q ;
  assign g22100 = \DFF_164.D ;
  assign g22101 = \DFF_187.D ;
  assign g22102 = \DFF_189.D ;
  assign g22103 = \DFF_191.D ;
  assign g22104 = \DFF_534.D ;
  assign g22105 = \DFF_536.D ;
  assign g22106 = \DFF_538.D ;
  assign g22107 = \DFF_709.D ;
  assign g2211 = \DFF_1428.Q ;
  assign g22112 = \DFF_881.D ;
  assign g22113 = \DFF_883.D ;
  assign g22114 = \DFF_885.D ;
  assign g22115 = \DFF_1228.D ;
  assign g22116 = \DFF_1230.D ;
  assign g22117 = \DFF_1232.D ;
  assign g22122 = \DFF_165.D ;
  assign g22123 = \DFF_167.D ;
  assign g22124 = \DFF_190.D ;
  assign g22125 = \DFF_192.D ;
  assign g22126 = \DFF_514.D ;
  assign g22127 = \DFF_537.D ;
  assign g22128 = \DFF_539.D ;
  assign g22129 = \DFF_541.D ;
  assign g22130 = \DFF_884.D ;
  assign g22131 = \DFF_886.D ;
  assign g22132 = \DFF_888.D ;
  assign g22133 = \DFF_1059.D ;
  assign g22138 = \DFF_1231.D ;
  assign g22139 = \DFF_1233.D ;
  assign g2214 = \DFF_1427.Q ;
  assign g22140 = \DFF_1235.D ;
  assign g22141 = \DFF_166.D ;
  assign g22142 = \DFF_168.D ;
  assign g22143 = \DFF_193.D ;
  assign g22145 = \DFF_515.D ;
  assign g22146 = \DFF_517.D ;
  assign g22147 = \DFF_540.D ;
  assign g22148 = \DFF_542.D ;
  assign g22149 = \DFF_864.D ;
  assign g22150 = \DFF_887.D ;
  assign g22151 = \DFF_889.D ;
  assign g22152 = \DFF_891.D ;
  assign g22153 = \DFF_1234.D ;
  assign g22154 = \DFF_1236.D ;
  assign g22155 = \DFF_1238.D ;
  assign g22156 = \DFF_1409.D ;
  assign g22161 = \DFF_169.D ;
  assign g22162 = \DFF_516.D ;
  assign g22163 = \DFF_518.D ;
  assign g22164 = \DFF_543.D ;
  assign g22166 = \DFF_865.D ;
  assign g22167 = \DFF_867.D ;
  assign g22168 = \DFF_890.D ;
  assign g22169 = \DFF_892.D ;
  assign g2217 = \DFF_1222.Q ;
  assign g22170 = \DFF_1214.D ;
  assign g22171 = \DFF_1237.D ;
  assign g22172 = \DFF_1239.D ;
  assign g22173 = \DFF_1241.D ;
  assign g22176 = \DFF_400.D ;
  assign g22177 = \DFF_519.D ;
  assign g22178 = \DFF_866.D ;
  assign g22179 = \DFF_868.D ;
  assign g2218 = \DFF_1220.Q ;
  assign g22180 = \DFF_893.D ;
  assign g22182 = \DFF_1215.D ;
  assign g22183 = \DFF_1217.D ;
  assign g22184 = \DFF_1240.D ;
  assign g22185 = \DFF_1242.D ;
  assign g2219 = \DFF_1221.Q ;
  assign g22191 = \DFF_869.D ;
  assign g22192 = \DFF_1216.D ;
  assign g22193 = \DFF_1218.D ;
  assign g22194 = \DFF_1243.D ;
  assign g222 = \DFF_230.Q ;
  assign g2220 = \DFF_1225.Q ;
  assign g22200 = \DFF_1219.D ;
  assign g2221 = \DFF_1223.Q ;
  assign g22218 = \DFF_508.D ;
  assign g2222 = \DFF_1224.Q ;
  assign g22225 = \DFF_63.D ;
  assign g22226 = \DFF_46.D ;
  assign g2223 = \DFF_1228.Q ;
  assign g22231 = \DFF_509.D ;
  assign g22234 = \DFF_858.D ;
  assign g2224 = \DFF_1226.Q ;
  assign g22242 = \DFF_510.D ;
  assign g22247 = \DFF_859.D ;
  assign g22249 = \DFF_1208.D ;
  assign g2225 = \DFF_1227.Q ;
  assign g22253 = \DFF_91.D ;
  assign g2226 = \DFF_1231.Q ;
  assign g22263 = \DFF_860.D ;
  assign g22267 = \DFF_1209.D ;
  assign g22269 = \DFF_1558.D ;
  assign g2227 = \DFF_1229.Q ;
  assign g2228 = \DFF_1230.Q ;
  assign g22280 = \DFF_1210.D ;
  assign g22284 = \DFF_1559.D ;
  assign g2229 = \DFF_1234.Q ;
  assign g22299 = \DFF_1560.D ;
  assign g2230 = \DFF_1232.Q ;
  assign g2231 = \DFF_1233.Q ;
  assign g2232 = \DFF_1237.Q ;
  assign g2233 = \DFF_1235.Q ;
  assign g2234 = \DFF_1236.Q ;
  assign g2235 = \DFF_1240.Q ;
  assign g2236 = \DFF_1238.Q ;
  assign g2237 = \DFF_1239.Q ;
  assign g2238 = \DFF_1243.Q ;
  assign g2239 = \DFF_1241.Q ;
  assign g2240 = \DFF_1242.Q ;
  assign g2241 = \DFF_1429.Q ;
  assign g2244 = \DFF_1246.Q ;
  assign g22444 = \DFF_81.D ;
  assign g2245 = \DFF_1244.Q ;
  assign g2246 = \DFF_1245.Q ;
  assign g2247 = \DFF_1249.Q ;
  assign g2248 = \DFF_1247.Q ;
  assign g2249 = \DFF_1248.Q ;
  assign g225 = \DFF_231.Q ;
  assign g2250 = \DFF_1252.Q ;
  assign g2251 = \DFF_1250.Q ;
  assign g22518 = \DFF_469.D ;
  assign g22519 = \DFF_496.D ;
  assign g2252 = \DFF_1251.Q ;
  assign g2253 = \DFF_1255.Q ;
  assign g2254 = \DFF_1253.Q ;
  assign g22548 = \DFF_470.D ;
  assign g22549 = \DFF_472.D ;
  assign g2255 = \DFF_1254.Q ;
  assign g22550 = \DFF_497.D ;
  assign g22551 = \DFF_442.D ;
  assign g22558 = \DFF_819.D ;
  assign g22559 = \DFF_846.D ;
  assign g2256 = \DFF_1296.Q ;
  assign g2257 = \DFF_1302.Q ;
  assign g22578 = \DFF_433.D ;
  assign g2258 = \DFF_1297.Q ;
  assign g22582 = \DFF_459.D ;
  assign g22583 = \DFF_471.D ;
  assign g22584 = \DFF_473.D ;
  assign g22585 = \DFF_475.D ;
  assign g22586 = \DFF_498.D ;
  assign g22589 = \DFF_820.D ;
  assign g22590 = \DFF_822.D ;
  assign g22591 = \DFF_847.D ;
  assign g22598 = \DFF_1169.D ;
  assign g22599 = \DFF_1196.D ;
  assign g2261 = \DFF_1256.Q ;
  assign g22611 = \DFF_474.D ;
  assign g22612 = \DFF_476.D ;
  assign g22613 = \DFF_478.D ;
  assign g22615 = \DFF_783.D ;
  assign g22619 = \DFF_809.D ;
  assign g22620 = \DFF_821.D ;
  assign g22621 = \DFF_823.D ;
  assign g22622 = \DFF_825.D ;
  assign g22623 = \DFF_848.D ;
  assign g22626 = \DFF_1170.D ;
  assign g22627 = \DFF_1172.D ;
  assign g22628 = \DFF_1197.D ;
  assign g22635 = \DFF_1519.D ;
  assign g22636 = \DFF_1546.D ;
  assign g22639 = \DFF_477.D ;
  assign g2264 = \DFF_1257.Q ;
  assign g22640 = \DFF_479.D ;
  assign g22641 = \DFF_481.D ;
  assign g22642 = \DFF_499.D ;
  assign g22647 = \DFF_824.D ;
  assign g22648 = \DFF_826.D ;
  assign g22649 = \DFF_828.D ;
  assign g22651 = \DFF_1133.D ;
  assign g22655 = \DFF_1159.D ;
  assign g22656 = \DFF_1171.D ;
  assign g22657 = \DFF_1173.D ;
  assign g22658 = \DFF_1175.D ;
  assign g22659 = \DFF_1198.D ;
  assign g22662 = \DFF_1520.D ;
  assign g22663 = \DFF_1522.D ;
  assign g22664 = \DFF_1547.D ;
  assign g22669 = \DFF_480.D ;
  assign g2267 = \DFF_1258.Q ;
  assign g22670 = \DFF_482.D ;
  assign g22671 = \DFF_484.D ;
  assign g22672 = \DFF_500.D ;
  assign g22673 = \DFF_502.D ;
  assign g22675 = \DFF_827.D ;
  assign g22676 = \DFF_829.D ;
  assign g22677 = \DFF_831.D ;
  assign g22678 = \DFF_849.D ;
  assign g22683 = \DFF_1174.D ;
  assign g22684 = \DFF_1176.D ;
  assign g22685 = \DFF_1178.D ;
  assign g22687 = \DFF_1483.D ;
  assign g22691 = \DFF_1509.D ;
  assign g22692 = \DFF_1521.D ;
  assign g22693 = \DFF_1523.D ;
  assign g22694 = \DFF_1525.D ;
  assign g22695 = \DFF_1548.D ;
  assign g2270 = \DFF_1262.Q ;
  assign g22702 = \DFF_483.D ;
  assign g22703 = \DFF_485.D ;
  assign g22704 = \DFF_487.D ;
  assign g22705 = \DFF_501.D ;
  assign g22706 = \DFF_503.D ;
  assign g22709 = \DFF_830.D ;
  assign g22710 = \DFF_832.D ;
  assign g22711 = \DFF_834.D ;
  assign g22712 = \DFF_850.D ;
  assign g22713 = \DFF_852.D ;
  assign g22715 = \DFF_1177.D ;
  assign g22716 = \DFF_1179.D ;
  assign g22717 = \DFF_1181.D ;
  assign g22718 = \DFF_1199.D ;
  assign g22723 = \DFF_1524.D ;
  assign g22724 = \DFF_1526.D ;
  assign g22725 = \DFF_1528.D ;
  assign g22728 = \DFF_486.D ;
  assign g22729 = \DFF_488.D ;
  assign g2273 = \DFF_1263.Q ;
  assign g22730 = \DFF_490.D ;
  assign g22731 = \DFF_504.D ;
  assign g22733 = \DFF_833.D ;
  assign g22734 = \DFF_835.D ;
  assign g22735 = \DFF_837.D ;
  assign g22736 = \DFF_851.D ;
  assign g22737 = \DFF_853.D ;
  assign g22740 = \DFF_1180.D ;
  assign g22741 = \DFF_1182.D ;
  assign g22742 = \DFF_1184.D ;
  assign g22743 = \DFF_1200.D ;
  assign g22744 = \DFF_1202.D ;
  assign g22746 = \DFF_1527.D ;
  assign g22747 = \DFF_1529.D ;
  assign g22748 = \DFF_1531.D ;
  assign g22749 = \DFF_1549.D ;
  assign g22756 = \DFF_489.D ;
  assign g22757 = \DFF_491.D ;
  assign g22758 = \DFF_493.D ;
  assign g2276 = \DFF_1264.Q ;
  assign g22760 = \DFF_836.D ;
  assign g22761 = \DFF_838.D ;
  assign g22762 = \DFF_840.D ;
  assign g22763 = \DFF_854.D ;
  assign g22765 = \DFF_1183.D ;
  assign g22766 = \DFF_1185.D ;
  assign g22767 = \DFF_1187.D ;
  assign g22768 = \DFF_1201.D ;
  assign g22769 = \DFF_1203.D ;
  assign g22772 = \DFF_1530.D ;
  assign g22773 = \DFF_1532.D ;
  assign g22774 = \DFF_1534.D ;
  assign g22775 = \DFF_1550.D ;
  assign g22776 = \DFF_1552.D ;
  assign g22785 = \DFF_492.D ;
  assign g22786 = \DFF_494.D ;
  assign g2279 = \DFF_1268.Q ;
  assign g22790 = \DFF_839.D ;
  assign g22791 = \DFF_841.D ;
  assign g22792 = \DFF_843.D ;
  assign g22794 = \DFF_1186.D ;
  assign g22795 = \DFF_1188.D ;
  assign g22796 = \DFF_1190.D ;
  assign g22797 = \DFF_1204.D ;
  assign g22799 = \DFF_1533.D ;
  assign g228 = \DFF_232.Q ;
  assign g22800 = \DFF_1535.D ;
  assign g22801 = \DFF_1537.D ;
  assign g22802 = \DFF_1551.D ;
  assign g22803 = \DFF_1553.D ;
  assign g2282 = \DFF_1269.Q ;
  assign g22824 = \DFF_495.D ;
  assign g22827 = \DFF_842.D ;
  assign g22828 = \DFF_844.D ;
  assign g22832 = \DFF_1189.D ;
  assign g22833 = \DFF_1191.D ;
  assign g22834 = \DFF_1193.D ;
  assign g22836 = \DFF_1536.D ;
  assign g22837 = \DFF_1538.D ;
  assign g22838 = \DFF_1540.D ;
  assign g22839 = \DFF_1554.D ;
  assign g22840 = \DFF_4.D ;
  assign g2285 = \DFF_1270.Q ;
  assign g22864 = \DFF_845.D ;
  assign g22866 = \DFF_1192.D ;
  assign g22867 = \DFF_1194.D ;
  assign g22871 = \DFF_1539.D ;
  assign g22872 = \DFF_1541.D ;
  assign g22873 = \DFF_1543.D ;
  assign g2288 = \DFF_1274.Q ;
  assign g22899 = \DFF_1195.D ;
  assign g22901 = \DFF_1542.D ;
  assign g22902 = \DFF_1544.D ;
  assign g2291 = \DFF_1275.Q ;
  assign g22934 = \DFF_1545.D ;
  assign g2294 = \DFF_1276.Q ;
  assign g22945 = \DFF_400.D ;
  assign g22948 = \DFF_1561.D ;
  assign g2297 = \DFF_1280.Q ;
  assign g22970 = \DFF_1562.D ;
  assign g22979 = \DFF_317.D ;
  assign g23 = \DFF_1625.Q ;
  assign g2300 = \DFF_1281.Q ;
  assign g23000 = \DFF_390.D ;
  assign g23014 = \DFF_740.D ;
  assign g23022 = \DFF_391.D ;
  assign g2303 = \DFF_1282.Q ;
  assign g23030 = \DFF_1090.D ;
  assign g23039 = \DFF_741.D ;
  assign g23047 = \DFF_1440.D ;
  assign g23055 = \DFF_442.D ;
  assign g23058 = \DFF_1091.D ;
  assign g2306 = \DFF_1259.Q ;
  assign g23067 = \DFF_380.D ;
  assign g23076 = \DFF_1441.D ;
  assign g23081 = \DFF_730.D ;
  assign g2309 = \DFF_1260.Q ;
  assign g23092 = \DFF_389.D ;
  assign g23093 = \DFF_381.D ;
  assign g23097 = \DFF_1080.D ;
  assign g231 = \DFF_209.Q ;
  assign g23110 = \DFF_739.D ;
  assign g23111 = \DFF_731.D ;
  assign g23114 = \DFF_1430.D ;
  assign g23116 = \DFF_317.D ;
  assign g23117 = \DFF_382.D ;
  assign g2312 = \DFF_1261.Q ;
  assign g23123 = \DFF_1089.D ;
  assign g23124 = \DFF_1081.D ;
  assign g23126 = \DFF_732.D ;
  assign g23132 = \DFF_1439.D ;
  assign g23133 = \DFF_1431.D ;
  assign g23136 = \DFF_460.D ;
  assign g23137 = \DFF_1082.D ;
  assign g23148 = \DFF_317.D ;
  assign g2315 = \DFF_1265.Q ;
  assign g23154 = \DFF_442.D ;
  assign g23159 = \DFF_400.D ;
  assign g23160 = \DFF_359.D ;
  assign g23161 = \DFF_459.D ;
  assign g23162 = \DFF_469.D ;
  assign g23163 = \DFF_470.D ;
  assign g23164 = \DFF_471.D ;
  assign g23165 = \DFF_472.D ;
  assign g23166 = \DFF_473.D ;
  assign g23167 = \DFF_474.D ;
  assign g23168 = \DFF_475.D ;
  assign g23169 = \DFF_476.D ;
  assign g23170 = \DFF_477.D ;
  assign g23171 = \DFF_478.D ;
  assign g23172 = \DFF_479.D ;
  assign g23173 = \DFF_480.D ;
  assign g23174 = \DFF_481.D ;
  assign g23175 = \DFF_482.D ;
  assign g23176 = \DFF_483.D ;
  assign g23177 = \DFF_484.D ;
  assign g23178 = \DFF_485.D ;
  assign g23179 = \DFF_486.D ;
  assign g2318 = \DFF_1266.Q ;
  assign g23180 = \DFF_487.D ;
  assign g23181 = \DFF_488.D ;
  assign g23182 = \DFF_489.D ;
  assign g23183 = \DFF_490.D ;
  assign g23184 = \DFF_491.D ;
  assign g23185 = \DFF_492.D ;
  assign g23186 = \DFF_493.D ;
  assign g23187 = \DFF_494.D ;
  assign g23188 = \DFF_495.D ;
  assign g23189 = \DFF_496.D ;
  assign g23190 = \DFF_497.D ;
  assign g23191 = \DFF_498.D ;
  assign g23192 = \DFF_499.D ;
  assign g23193 = \DFF_500.D ;
  assign g23194 = \DFF_501.D ;
  assign g23195 = \DFF_502.D ;
  assign g23196 = \DFF_503.D ;
  assign g23197 = \DFF_504.D ;
  assign g23198 = \DFF_709.D ;
  assign g23199 = \DFF_809.D ;
  assign g23200 = \DFF_819.D ;
  assign g23201 = \DFF_820.D ;
  assign g23202 = \DFF_821.D ;
  assign g23203 = \DFF_822.D ;
  assign g23204 = \DFF_823.D ;
  assign g23205 = \DFF_824.D ;
  assign g23206 = \DFF_825.D ;
  assign g23207 = \DFF_826.D ;
  assign g23208 = \DFF_827.D ;
  assign g23209 = \DFF_828.D ;
  assign g2321 = \DFF_1267.Q ;
  assign g23210 = \DFF_829.D ;
  assign g23211 = \DFF_830.D ;
  assign g23212 = \DFF_831.D ;
  assign g23213 = \DFF_832.D ;
  assign g23214 = \DFF_833.D ;
  assign g23215 = \DFF_834.D ;
  assign g23216 = \DFF_835.D ;
  assign g23217 = \DFF_836.D ;
  assign g23218 = \DFF_837.D ;
  assign g23219 = \DFF_838.D ;
  assign g23220 = \DFF_839.D ;
  assign g23221 = \DFF_840.D ;
  assign g23222 = \DFF_841.D ;
  assign g23223 = \DFF_842.D ;
  assign g23224 = \DFF_843.D ;
  assign g23225 = \DFF_844.D ;
  assign g23226 = \DFF_845.D ;
  assign g23227 = \DFF_846.D ;
  assign g23228 = \DFF_847.D ;
  assign g23229 = \DFF_848.D ;
  assign g23230 = \DFF_849.D ;
  assign g23231 = \DFF_850.D ;
  assign g23232 = \DFF_851.D ;
  assign g23233 = \DFF_852.D ;
  assign g23234 = \DFF_853.D ;
  assign g23235 = \DFF_854.D ;
  assign g23236 = \DFF_1059.D ;
  assign g23237 = \DFF_1159.D ;
  assign g23238 = \DFF_1169.D ;
  assign g23239 = \DFF_1170.D ;
  assign g2324 = \DFF_1271.Q ;
  assign g23240 = \DFF_1171.D ;
  assign g23241 = \DFF_1172.D ;
  assign g23242 = \DFF_1173.D ;
  assign g23243 = \DFF_1174.D ;
  assign g23244 = \DFF_1175.D ;
  assign g23245 = \DFF_1176.D ;
  assign g23246 = \DFF_1177.D ;
  assign g23247 = \DFF_1178.D ;
  assign g23248 = \DFF_1179.D ;
  assign g23249 = \DFF_1180.D ;
  assign g23250 = \DFF_1181.D ;
  assign g23251 = \DFF_1182.D ;
  assign g23252 = \DFF_1183.D ;
  assign g23253 = \DFF_1184.D ;
  assign g23254 = \DFF_1185.D ;
  assign g23255 = \DFF_1186.D ;
  assign g23256 = \DFF_1187.D ;
  assign g23257 = \DFF_1188.D ;
  assign g23258 = \DFF_1189.D ;
  assign g23259 = \DFF_1190.D ;
  assign g23260 = \DFF_1191.D ;
  assign g23261 = \DFF_1192.D ;
  assign g23262 = \DFF_1193.D ;
  assign g23263 = \DFF_1194.D ;
  assign g23264 = \DFF_1195.D ;
  assign g23265 = \DFF_1196.D ;
  assign g23266 = \DFF_1197.D ;
  assign g23267 = \DFF_1198.D ;
  assign g23268 = \DFF_1199.D ;
  assign g23269 = \DFF_1200.D ;
  assign g2327 = \DFF_1272.Q ;
  assign g23270 = \DFF_1201.D ;
  assign g23271 = \DFF_1202.D ;
  assign g23272 = \DFF_1203.D ;
  assign g23273 = \DFF_1204.D ;
  assign g23274 = \DFF_1409.D ;
  assign g23275 = \DFF_1509.D ;
  assign g23276 = \DFF_1519.D ;
  assign g23277 = \DFF_1520.D ;
  assign g23278 = \DFF_1521.D ;
  assign g23279 = \DFF_1522.D ;
  assign g23280 = \DFF_1523.D ;
  assign g23281 = \DFF_1524.D ;
  assign g23282 = \DFF_1525.D ;
  assign g23283 = \DFF_1526.D ;
  assign g23284 = \DFF_1527.D ;
  assign g23285 = \DFF_1528.D ;
  assign g23286 = \DFF_1529.D ;
  assign g23287 = \DFF_1530.D ;
  assign g23288 = \DFF_1531.D ;
  assign g23289 = \DFF_1532.D ;
  assign g23290 = \DFF_1533.D ;
  assign g23291 = \DFF_1534.D ;
  assign g23292 = \DFF_1535.D ;
  assign g23293 = \DFF_1536.D ;
  assign g23294 = \DFF_1537.D ;
  assign g23295 = \DFF_1538.D ;
  assign g23296 = \DFF_1539.D ;
  assign g23297 = \DFF_1540.D ;
  assign g23298 = \DFF_1541.D ;
  assign g23299 = \DFF_1542.D ;
  assign g2330 = \DFF_1273.Q ;
  assign g23300 = \DFF_1543.D ;
  assign g23301 = \DFF_1544.D ;
  assign g23302 = \DFF_1545.D ;
  assign g23303 = \DFF_1546.D ;
  assign g23304 = \DFF_1547.D ;
  assign g23305 = \DFF_1548.D ;
  assign g23306 = \DFF_1549.D ;
  assign g23307 = \DFF_1550.D ;
  assign g23308 = \DFF_1551.D ;
  assign g23309 = \DFF_1552.D ;
  assign g23310 = \DFF_1553.D ;
  assign g23311 = \DFF_1554.D ;
  assign g23312 = \DFF_63.D ;
  assign g23313 = \DFF_46.D ;
  assign g23314 = \DFF_91.D ;
  assign g23315 = \DFF_4.D ;
  assign g23316 = \DFF_81.D ;
  assign g23317 = \DFF_1561.D ;
  assign g23318 = \DFF_1562.D ;
  assign g23324 = \DFF_461.D ;
  assign g23329 = \DFF_811.D ;
  assign g2333 = \DFF_1277.Q ;
  assign g23330 = \DFF_1602.D ;
  assign g23339 = \DFF_1161.D ;
  assign g23348 = \DFF_1511.D ;
  assign g23357 = \DFF_12.D ;
  assign g23358 = \DFF_6.D ;
  assign g23359 = \DFF_1608.D ;
  assign g2336 = \DFF_1278.Q ;
  assign g23385 = \DFF_383.D ;
  assign g2339 = \DFF_1279.Q ;
  assign g23392 = \DFF_733.D ;
  assign g23399 = \DFF_384.D ;
  assign g234 = \DFF_210.Q ;
  assign g23400 = \DFF_1083.D ;
  assign g23406 = \DFF_734.D ;
  assign g23407 = \DFF_1433.D ;
  assign g23413 = \DFF_1084.D ;
  assign g23418 = \DFF_1434.D ;
  assign g2342 = \DFF_1283.Q ;
  assign g23438 = \DFF_390.D ;
  assign g23439 = \DFF_382.D ;
  assign g2345 = \DFF_1284.Q ;
  assign g23452 = \DFF_740.D ;
  assign g23453 = \DFF_732.D ;
  assign g23454 = \DFF_391.D ;
  assign g23459 = \DFF_1090.D ;
  assign g23460 = \DFF_1082.D ;
  assign g23463 = \DFF_741.D ;
  assign g23468 = \DFF_1440.D ;
  assign g23469 = \DFF_1432.D ;
  assign g23472 = \DFF_1091.D ;
  assign g2348 = \DFF_1285.Q ;
  assign g23481 = \DFF_380.D ;
  assign g23485 = \DFF_1441.D ;
  assign g23492 = \DFF_730.D ;
  assign g23500 = \DFF_389.D ;
  assign g23501 = \DFF_381.D ;
  assign g23508 = \DFF_1080.D ;
  assign g2351 = \DFF_1427.Q ;
  assign g23516 = \DFF_739.D ;
  assign g23517 = \DFF_731.D ;
  assign g23524 = \DFF_1430.D ;
  assign g23531 = \DFF_1089.D ;
  assign g23532 = \DFF_1081.D ;
  assign g2354 = \DFF_1353.Q ;
  assign g23542 = \DFF_1439.D ;
  assign g23543 = \DFF_1431.D ;
  assign g23546 = \DFF_170.D ;
  assign g23548 = \DFF_171.D ;
  assign g23549 = \DFF_173.D ;
  assign g2355 = \DFF_1354.Q ;
  assign g23553 = \DFF_520.D ;
  assign g23555 = \DFF_172.D ;
  assign g23556 = \DFF_174.D ;
  assign g23557 = \DFF_176.D ;
  assign g2356 = \DFF_1355.Q ;
  assign g23561 = \DFF_521.D ;
  assign g23562 = \DFF_523.D ;
  assign g23566 = \DFF_870.D ;
  assign g23568 = \DFF_175.D ;
  assign g23569 = \DFF_177.D ;
  assign g2357 = \DFF_1356.Q ;
  assign g23570 = \DFF_179.D ;
  assign g23574 = \DFF_522.D ;
  assign g23575 = \DFF_524.D ;
  assign g23576 = \DFF_526.D ;
  assign g2358 = \DFF_1357.Q ;
  assign g23580 = \DFF_871.D ;
  assign g23581 = \DFF_873.D ;
  assign g23585 = \DFF_1220.D ;
  assign g23587 = \DFF_178.D ;
  assign g23588 = \DFF_180.D ;
  assign g23589 = \DFF_182.D ;
  assign g2359 = \DFF_1358.Q ;
  assign g23594 = \DFF_460.D ;
  assign g23595 = \DFF_525.D ;
  assign g23596 = \DFF_527.D ;
  assign g23597 = \DFF_529.D ;
  assign g2360 = \DFF_1359.Q ;
  assign g23601 = \DFF_872.D ;
  assign g23602 = \DFF_874.D ;
  assign g23603 = \DFF_876.D ;
  assign g23607 = \DFF_1221.D ;
  assign g23608 = \DFF_1223.D ;
  assign g2361 = \DFF_1360.Q ;
  assign g23612 = \DFF_181.D ;
  assign g23613 = \DFF_183.D ;
  assign g23614 = \DFF_185.D ;
  assign g23619 = \DFF_528.D ;
  assign g2362 = \DFF_1361.Q ;
  assign g23620 = \DFF_530.D ;
  assign g23621 = \DFF_532.D ;
  assign g23626 = \DFF_810.D ;
  assign g23627 = \DFF_875.D ;
  assign g23628 = \DFF_877.D ;
  assign g23629 = \DFF_879.D ;
  assign g2363 = \DFF_1362.Q ;
  assign g23633 = \DFF_1222.D ;
  assign g23634 = \DFF_1224.D ;
  assign g23635 = \DFF_1226.D ;
  assign g2364 = \DFF_1363.Q ;
  assign g23640 = \DFF_184.D ;
  assign g23641 = \DFF_186.D ;
  assign g23642 = \DFF_188.D ;
  assign g2365 = \DFF_1364.Q ;
  assign g2366 = \DFF_1365.Q ;
  assign g23661 = \DFF_531.D ;
  assign g23662 = \DFF_533.D ;
  assign g23663 = \DFF_535.D ;
  assign g23668 = \DFF_878.D ;
  assign g23669 = \DFF_880.D ;
  assign g23670 = \DFF_882.D ;
  assign g23675 = \DFF_1160.D ;
  assign g23676 = \DFF_1225.D ;
  assign g23677 = \DFF_1227.D ;
  assign g23678 = \DFF_1229.D ;
  assign g23682 = \DFF_164.D ;
  assign g23683 = \DFF_187.D ;
  assign g23684 = \DFF_189.D ;
  assign g23685 = \DFF_191.D ;
  assign g23690 = \DFF_534.D ;
  assign g23691 = \DFF_536.D ;
  assign g23692 = \DFF_538.D ;
  assign g237 = \DFF_211.Q ;
  assign g23711 = \DFF_881.D ;
  assign g23712 = \DFF_883.D ;
  assign g23713 = \DFF_885.D ;
  assign g23718 = \DFF_1228.D ;
  assign g23719 = \DFF_1230.D ;
  assign g23720 = \DFF_1232.D ;
  assign g23725 = \DFF_1510.D ;
  assign g23727 = \DFF_165.D ;
  assign g23728 = \DFF_167.D ;
  assign g23729 = \DFF_190.D ;
  assign g2373 = \DFF_1378.Q ;
  assign g23730 = \DFF_192.D ;
  assign g23736 = \DFF_514.D ;
  assign g23737 = \DFF_537.D ;
  assign g23738 = \DFF_539.D ;
  assign g23739 = \DFF_541.D ;
  assign g2374 = \DFF_1366.Q ;
  assign g23744 = \DFF_884.D ;
  assign g23745 = \DFF_886.D ;
  assign g23746 = \DFF_888.D ;
  assign g23765 = \DFF_1231.D ;
  assign g23766 = \DFF_1233.D ;
  assign g23767 = \DFF_1235.D ;
  assign g23773 = \DFF_166.D ;
  assign g23774 = \DFF_168.D ;
  assign g23775 = \DFF_193.D ;
  assign g23782 = \DFF_515.D ;
  assign g23783 = \DFF_517.D ;
  assign g23784 = \DFF_540.D ;
  assign g23785 = \DFF_542.D ;
  assign g23791 = \DFF_864.D ;
  assign g23792 = \DFF_887.D ;
  assign g23793 = \DFF_889.D ;
  assign g23794 = \DFF_891.D ;
  assign g23799 = \DFF_1234.D ;
  assign g2380 = \DFF_1367.Q ;
  assign g23800 = \DFF_1236.D ;
  assign g23801 = \DFF_1238.D ;
  assign g23821 = \DFF_169.D ;
  assign g23826 = \DFF_516.D ;
  assign g23827 = \DFF_518.D ;
  assign g23828 = \DFF_543.D ;
  assign g23835 = \DFF_865.D ;
  assign g23836 = \DFF_867.D ;
  assign g23837 = \DFF_890.D ;
  assign g23838 = \DFF_892.D ;
  assign g2384 = \DFF_1302.Q ;
  assign g23844 = \DFF_1214.D ;
  assign g23845 = \DFF_1237.D ;
  assign g23846 = \DFF_1239.D ;
  assign g23847 = \DFF_1241.D ;
  assign g23856 = \DFF_519.D ;
  assign g23861 = \DFF_866.D ;
  assign g23862 = \DFF_868.D ;
  assign g23863 = \DFF_893.D ;
  assign g2387 = \DFF_1333.Q ;
  assign g23870 = \DFF_1215.D ;
  assign g23871 = \DFF_1217.D ;
  assign g23872 = \DFF_1240.D ;
  assign g23873 = \DFF_1242.D ;
  assign g2388 = \DFF_1334.Q ;
  assign g2389 = \DFF_1335.Q ;
  assign g23890 = \DFF_869.D ;
  assign g23895 = \DFF_1216.D ;
  assign g23896 = \DFF_1218.D ;
  assign g23897 = \DFF_1243.D ;
  assign g2390 = \DFF_1336.Q ;
  assign g2391 = \DFF_1337.Q ;
  assign g23911 = \DFF_1219.D ;
  assign g23916 = \DFF_11.D ;
  assign g23919 = \DFF_131.D ;
  assign g2392 = \DFF_1338.Q ;
  assign g23923 = \DFF_433.D ;
  assign g2393 = \DFF_1339.Q ;
  assign g2394 = \DFF_1340.Q ;
  assign g23943 = \DFF_1607.D ;
  assign g2395 = \DFF_1341.Q ;
  assign g23955 = \DFF_783.D ;
  assign g2396 = \DFF_1344.Q ;
  assign g2397 = \DFF_1342.Q ;
  assign g2398 = \DFF_1343.Q ;
  assign g23984 = \DFF_1133.D ;
  assign g2399 = \DFF_1402.Q ;
  assign g240 = \DFF_215.Q ;
  assign g2400 = \DFF_1504.Q ;
  assign g24000 = \DFF_5.D ;
  assign g24001 = \DFF_508.D ;
  assign g24014 = \DFF_1483.D ;
  assign g24033 = \DFF_509.D ;
  assign g24035 = \DFF_858.D ;
  assign g24051 = \DFF_510.D ;
  assign g24053 = \DFF_859.D ;
  assign g24055 = \DFF_1208.D ;
  assign g24059 = \DFF_452.D ;
  assign g2406 = \DFF_1505.Q ;
  assign g24064 = \DFF_860.D ;
  assign g24066 = \DFF_1209.D ;
  assign g24068 = \DFF_1558.D ;
  assign g24072 = \DFF_802.D ;
  assign g24077 = \DFF_1210.D ;
  assign g24079 = \DFF_1559.D ;
  assign g24083 = \DFF_1152.D ;
  assign g24088 = \DFF_1560.D ;
  assign g24092 = \DFF_1502.D ;
  assign g2412 = \DFF_1506.Q ;
  assign g2417 = \DFF_1379.Q ;
  assign g24174 = \DFF_385.D ;
  assign g24178 = \DFF_386.D ;
  assign g24179 = \DFF_735.D ;
  assign g2418 = \DFF_1304.Q ;
  assign g24181 = \DFF_736.D ;
  assign g24182 = \DFF_1085.D ;
  assign g24206 = \DFF_392.D ;
  assign g24207 = \DFF_387.D ;
  assign g24208 = \DFF_1086.D ;
  assign g24209 = \DFF_1435.D ;
  assign g2421 = \DFF_1305.Q ;
  assign g24212 = \DFF_742.D ;
  assign g24213 = \DFF_737.D ;
  assign g24214 = \DFF_1436.D ;
  assign g24215 = \DFF_393.D ;
  assign g24216 = \DFF_388.D ;
  assign g24218 = \DFF_1092.D ;
  assign g24219 = \DFF_1087.D ;
  assign g24222 = \DFF_743.D ;
  assign g24223 = \DFF_738.D ;
  assign g24225 = \DFF_1442.D ;
  assign g24226 = \DFF_1437.D ;
  assign g24228 = \DFF_394.D ;
  assign g24230 = \DFF_1093.D ;
  assign g24231 = \DFF_1088.D ;
  assign g24233 = \DFF_433.D ;
  assign g24235 = \DFF_744.D ;
  assign g24237 = \DFF_1443.D ;
  assign g24238 = \DFF_1438.D ;
  assign g2424 = \DFF_1380.Q ;
  assign g24240 = \DFF_783.D ;
  assign g24243 = \DFF_1094.D ;
  assign g24248 = \DFF_1133.D ;
  assign g2425 = \DFF_1381.Q ;
  assign g24250 = \DFF_1444.D ;
  assign g24255 = \DFF_1483.D ;
  assign g24259 = \DFF_164.D ;
  assign g2426 = \DFF_1382.Q ;
  assign g24260 = \DFF_165.D ;
  assign g24261 = \DFF_166.D ;
  assign g24262 = \DFF_167.D ;
  assign g24263 = \DFF_168.D ;
  assign g24264 = \DFF_169.D ;
  assign g24265 = \DFF_170.D ;
  assign g24266 = \DFF_171.D ;
  assign g24267 = \DFF_172.D ;
  assign g24268 = \DFF_173.D ;
  assign g24269 = \DFF_174.D ;
  assign g2427 = \DFF_1383.Q ;
  assign g24270 = \DFF_175.D ;
  assign g24271 = \DFF_176.D ;
  assign g24272 = \DFF_177.D ;
  assign g24273 = \DFF_178.D ;
  assign g24274 = \DFF_179.D ;
  assign g24275 = \DFF_180.D ;
  assign g24276 = \DFF_181.D ;
  assign g24277 = \DFF_182.D ;
  assign g24278 = \DFF_183.D ;
  assign g24279 = \DFF_184.D ;
  assign g2428 = \DFF_1384.Q ;
  assign g24280 = \DFF_185.D ;
  assign g24281 = \DFF_186.D ;
  assign g24282 = \DFF_187.D ;
  assign g24283 = \DFF_188.D ;
  assign g24284 = \DFF_189.D ;
  assign g24285 = \DFF_190.D ;
  assign g24286 = \DFF_191.D ;
  assign g24287 = \DFF_192.D ;
  assign g24288 = \DFF_193.D ;
  assign g24289 = \DFF_389.D ;
  assign g2429 = \DFF_1303.Q ;
  assign g24290 = \DFF_390.D ;
  assign g24291 = \DFF_391.D ;
  assign g24292 = \DFF_380.D ;
  assign g24293 = \DFF_381.D ;
  assign g24294 = \DFF_382.D ;
  assign g24295 = \DFF_433.D ;
  assign g24296 = \DFF_460.D ;
  assign g24297 = \DFF_508.D ;
  assign g24298 = \DFF_509.D ;
  assign g24299 = \DFF_510.D ;
  assign g243 = \DFF_216.Q ;
  assign g24300 = \DFF_514.D ;
  assign g24301 = \DFF_515.D ;
  assign g24302 = \DFF_516.D ;
  assign g24303 = \DFF_517.D ;
  assign g24304 = \DFF_518.D ;
  assign g24305 = \DFF_519.D ;
  assign g24306 = \DFF_520.D ;
  assign g24307 = \DFF_521.D ;
  assign g24308 = \DFF_522.D ;
  assign g24309 = \DFF_523.D ;
  assign g24310 = \DFF_524.D ;
  assign g24311 = \DFF_525.D ;
  assign g24312 = \DFF_526.D ;
  assign g24313 = \DFF_527.D ;
  assign g24314 = \DFF_528.D ;
  assign g24315 = \DFF_529.D ;
  assign g24316 = \DFF_530.D ;
  assign g24317 = \DFF_531.D ;
  assign g24318 = \DFF_532.D ;
  assign g24319 = \DFF_533.D ;
  assign g2432 = \DFF_1385.Q ;
  assign g24320 = \DFF_534.D ;
  assign g24321 = \DFF_535.D ;
  assign g24322 = \DFF_536.D ;
  assign g24323 = \DFF_537.D ;
  assign g24324 = \DFF_538.D ;
  assign g24325 = \DFF_539.D ;
  assign g24326 = \DFF_540.D ;
  assign g24327 = \DFF_541.D ;
  assign g24328 = \DFF_542.D ;
  assign g24329 = \DFF_543.D ;
  assign g2433 = \DFF_1307.Q ;
  assign g24330 = \DFF_739.D ;
  assign g24331 = \DFF_740.D ;
  assign g24332 = \DFF_741.D ;
  assign g24333 = \DFF_730.D ;
  assign g24334 = \DFF_731.D ;
  assign g24335 = \DFF_732.D ;
  assign g24336 = \DFF_783.D ;
  assign g24337 = \DFF_810.D ;
  assign g24338 = \DFF_858.D ;
  assign g24339 = \DFF_859.D ;
  assign g24340 = \DFF_860.D ;
  assign g24341 = \DFF_864.D ;
  assign g24342 = \DFF_865.D ;
  assign g24343 = \DFF_866.D ;
  assign g24344 = \DFF_867.D ;
  assign g24345 = \DFF_868.D ;
  assign g24346 = \DFF_869.D ;
  assign g24347 = \DFF_870.D ;
  assign g24348 = \DFF_871.D ;
  assign g24349 = \DFF_872.D ;
  assign g24350 = \DFF_873.D ;
  assign g24351 = \DFF_874.D ;
  assign g24352 = \DFF_875.D ;
  assign g24353 = \DFF_876.D ;
  assign g24354 = \DFF_877.D ;
  assign g24355 = \DFF_878.D ;
  assign g24356 = \DFF_879.D ;
  assign g24357 = \DFF_880.D ;
  assign g24358 = \DFF_881.D ;
  assign g24359 = \DFF_882.D ;
  assign g2436 = \DFF_1308.Q ;
  assign g24360 = \DFF_883.D ;
  assign g24361 = \DFF_884.D ;
  assign g24362 = \DFF_885.D ;
  assign g24363 = \DFF_886.D ;
  assign g24364 = \DFF_887.D ;
  assign g24365 = \DFF_888.D ;
  assign g24366 = \DFF_889.D ;
  assign g24367 = \DFF_890.D ;
  assign g24368 = \DFF_891.D ;
  assign g24369 = \DFF_892.D ;
  assign g24370 = \DFF_893.D ;
  assign g24371 = \DFF_1089.D ;
  assign g24372 = \DFF_1090.D ;
  assign g24373 = \DFF_1091.D ;
  assign g24374 = \DFF_1080.D ;
  assign g24375 = \DFF_1081.D ;
  assign g24376 = \DFF_1082.D ;
  assign g24377 = \DFF_1133.D ;
  assign g24378 = \DFF_1160.D ;
  assign g24379 = \DFF_1208.D ;
  assign g24380 = \DFF_1209.D ;
  assign g24381 = \DFF_1210.D ;
  assign g24382 = \DFF_1214.D ;
  assign g24383 = \DFF_1215.D ;
  assign g24384 = \DFF_1216.D ;
  assign g24385 = \DFF_1217.D ;
  assign g24386 = \DFF_1218.D ;
  assign g24387 = \DFF_1219.D ;
  assign g24388 = \DFF_1220.D ;
  assign g24389 = \DFF_1221.D ;
  assign g2439 = \DFF_1386.Q ;
  assign g24390 = \DFF_1222.D ;
  assign g24391 = \DFF_1223.D ;
  assign g24392 = \DFF_1224.D ;
  assign g24393 = \DFF_1225.D ;
  assign g24394 = \DFF_1226.D ;
  assign g24395 = \DFF_1227.D ;
  assign g24396 = \DFF_1228.D ;
  assign g24397 = \DFF_1229.D ;
  assign g24398 = \DFF_1230.D ;
  assign g24399 = \DFF_1231.D ;
  assign g2440 = \DFF_1387.Q ;
  assign g24400 = \DFF_1232.D ;
  assign g24401 = \DFF_1233.D ;
  assign g24402 = \DFF_1234.D ;
  assign g24403 = \DFF_1235.D ;
  assign g24404 = \DFF_1236.D ;
  assign g24405 = \DFF_1237.D ;
  assign g24406 = \DFF_1238.D ;
  assign g24407 = \DFF_1239.D ;
  assign g24408 = \DFF_1240.D ;
  assign g24409 = \DFF_1241.D ;
  assign g2441 = \DFF_1388.Q ;
  assign g24410 = \DFF_1242.D ;
  assign g24411 = \DFF_1243.D ;
  assign g24412 = \DFF_1439.D ;
  assign g24413 = \DFF_1440.D ;
  assign g24414 = \DFF_1441.D ;
  assign g24415 = \DFF_1430.D ;
  assign g24416 = \DFF_1431.D ;
  assign g24417 = \DFF_1432.D ;
  assign g24418 = \DFF_1483.D ;
  assign g24419 = \DFF_1510.D ;
  assign g2442 = \DFF_1389.Q ;
  assign g24420 = \DFF_1558.D ;
  assign g24421 = \DFF_1559.D ;
  assign g24422 = \DFF_1560.D ;
  assign g24423 = \DFF_5.D ;
  assign g24424 = \DFF_11.D ;
  assign g24425 = \DFF_1607.D ;
  assign g24426 = \DFF_462.D ;
  assign g2443 = \DFF_1390.Q ;
  assign g24430 = \DFF_812.D ;
  assign g24434 = \DFF_1162.D ;
  assign g24438 = \DFF_1512.D ;
  assign g2444 = \DFF_1306.Q ;
  assign g24445 = \DFF_1603.D ;
  assign g24446 = \DFF_1609.D ;
  assign g2447 = \DFF_1391.Q ;
  assign g24473 = \DFF_7.D ;
  assign g24476 = \DFF_13.D ;
  assign g2448 = \DFF_1310.Q ;
  assign g24491 = \DFF_417.D ;
  assign g24498 = \DFF_418.D ;
  assign g24499 = \DFF_420.D ;
  assign g24501 = \DFF_767.D ;
  assign g24507 = \DFF_419.D ;
  assign g24508 = \DFF_421.D ;
  assign g2451 = \DFF_1311.Q ;
  assign g24510 = \DFF_768.D ;
  assign g24511 = \DFF_770.D ;
  assign g24513 = \DFF_1117.D ;
  assign g24518 = \DFF_384.D ;
  assign g24519 = \DFF_422.D ;
  assign g24521 = \DFF_769.D ;
  assign g24522 = \DFF_771.D ;
  assign g24524 = \DFF_1118.D ;
  assign g24525 = \DFF_1120.D ;
  assign g24527 = \DFF_1467.D ;
  assign g24531 = \DFF_734.D ;
  assign g24532 = \DFF_772.D ;
  assign g24534 = \DFF_1119.D ;
  assign g24535 = \DFF_1121.D ;
  assign g24537 = \DFF_1468.D ;
  assign g24538 = \DFF_1470.D ;
  assign g24539 = \DFF_385.D ;
  assign g2454 = \DFF_1392.Q ;
  assign g24544 = \DFF_1084.D ;
  assign g24545 = \DFF_1122.D ;
  assign g24547 = \DFF_1469.D ;
  assign g24548 = \DFF_1471.D ;
  assign g24549 = \DFF_386.D ;
  assign g2455 = \DFF_1393.Q ;
  assign g24551 = \DFF_735.D ;
  assign g24556 = \DFF_1434.D ;
  assign g24557 = \DFF_1472.D ;
  assign g2456 = \DFF_1394.Q ;
  assign g24560 = \DFF_736.D ;
  assign g24562 = \DFF_1085.D ;
  assign g24567 = \DFF_392.D ;
  assign g24568 = \DFF_387.D ;
  assign g2457 = \DFF_1395.Q ;
  assign g24570 = \DFF_1086.D ;
  assign g24572 = \DFF_1435.D ;
  assign g24576 = \DFF_742.D ;
  assign g24577 = \DFF_737.D ;
  assign g24579 = \DFF_1436.D ;
  assign g2458 = \DFF_1396.Q ;
  assign g24581 = \DFF_393.D ;
  assign g24582 = \DFF_388.D ;
  assign g24583 = \DFF_1092.D ;
  assign g24584 = \DFF_1087.D ;
  assign g24586 = \DFF_743.D ;
  assign g24587 = \DFF_738.D ;
  assign g24588 = \DFF_1442.D ;
  assign g24589 = \DFF_1437.D ;
  assign g2459 = \DFF_1309.Q ;
  assign g24592 = \DFF_394.D ;
  assign g24593 = \DFF_1093.D ;
  assign g24594 = \DFF_1088.D ;
  assign g24597 = \DFF_744.D ;
  assign g24598 = \DFF_1443.D ;
  assign g24599 = \DFF_1438.D ;
  assign g246 = \DFF_217.Q ;
  assign g24605 = \DFF_1094.D ;
  assign g24612 = \DFF_1444.D ;
  assign g2462 = \DFF_1397.Q ;
  assign g2463 = \DFF_1313.Q ;
  assign g2466 = \DFF_1314.Q ;
  assign g2469 = \DFF_1398.Q ;
  assign g2470 = \DFF_1399.Q ;
  assign g2471 = \DFF_1400.Q ;
  assign g2472 = \DFF_1401.Q ;
  assign g2473 = \DFF_1312.Q ;
  assign g24734 = \DFF_131.D ;
  assign g24735 = \DFF_131.D ;
  assign g2476 = \DFF_1429.Q ;
  assign g2477 = \DFF_1347.Q ;
  assign g2478 = \DFF_1345.Q ;
  assign g2479 = \DFF_1346.Q ;
  assign g2480 = \DFF_1428.Q ;
  assign g24816 = \DFF_383.D ;
  assign g2483 = \DFF_1315.Q ;
  assign g24835 = \DFF_733.D ;
  assign g24851 = \DFF_1083.D ;
  assign g24856 = \DFF_461.D ;
  assign g2486 = \DFF_1316.Q ;
  assign g24865 = \DFF_1433.D ;
  assign g24872 = \DFF_811.D ;
  assign g24879 = \DFF_1602.D ;
  assign g24886 = \DFF_1161.D ;
  assign g2489 = \DFF_1317.Q ;
  assign g24890 = \DFF_150.D ;
  assign g249 = \DFF_221.Q ;
  assign g24903 = \DFF_1511.D ;
  assign g24909 = \DFF_151.D ;
  assign g2492 = \DFF_1318.Q ;
  assign g24925 = \DFF_152.D ;
  assign g24949 = \DFF_12.D ;
  assign g2495 = \DFF_1319.Q ;
  assign g24956 = \DFF_6.D ;
  assign g24957 = \DFF_1608.D ;
  assign g2498 = \DFF_1320.Q ;
  assign g2501 = \DFF_1323.Q ;
  assign g2502 = \DFF_1321.Q ;
  assign g25027 = \DFF_236.D ;
  assign g2503 = \DFF_1322.Q ;
  assign g2504 = \DFF_1324.Q ;
  assign g25042 = \DFF_586.D ;
  assign g25056 = \DFF_936.D ;
  assign g25067 = \DFF_1286.D ;
  assign g2507 = \DFF_1325.Q ;
  assign g2510 = \DFF_1326.Q ;
  assign g25103 = \DFF_452.D ;
  assign g25109 = \DFF_802.D ;
  assign g25119 = \DFF_1152.D ;
  assign g25122 = \DFF_1502.D ;
  assign g2513 = \DFF_1327.Q ;
  assign g25131 = \DFF_384.D ;
  assign g25132 = \DFF_385.D ;
  assign g25133 = \DFF_392.D ;
  assign g25134 = \DFF_393.D ;
  assign g25135 = \DFF_394.D ;
  assign g25136 = \DFF_386.D ;
  assign g25137 = \DFF_387.D ;
  assign g25138 = \DFF_388.D ;
  assign g25139 = \DFF_383.D ;
  assign g25140 = \DFF_461.D ;
  assign g25142 = \DFF_734.D ;
  assign g25143 = \DFF_735.D ;
  assign g25144 = \DFF_742.D ;
  assign g25145 = \DFF_743.D ;
  assign g25146 = \DFF_744.D ;
  assign g25147 = \DFF_736.D ;
  assign g25148 = \DFF_737.D ;
  assign g25149 = \DFF_738.D ;
  assign g25150 = \DFF_733.D ;
  assign g25151 = \DFF_811.D ;
  assign g25153 = \DFF_1084.D ;
  assign g25154 = \DFF_1085.D ;
  assign g25155 = \DFF_1092.D ;
  assign g25156 = \DFF_1093.D ;
  assign g25157 = \DFF_1094.D ;
  assign g25158 = \DFF_1086.D ;
  assign g25159 = \DFF_1087.D ;
  assign g2516 = \DFF_1328.Q ;
  assign g25160 = \DFF_1088.D ;
  assign g25161 = \DFF_1083.D ;
  assign g25162 = \DFF_1161.D ;
  assign g25164 = \DFF_1434.D ;
  assign g25165 = \DFF_1435.D ;
  assign g25166 = \DFF_1442.D ;
  assign g25167 = \DFF_1443.D ;
  assign g25168 = \DFF_1444.D ;
  assign g25169 = \DFF_1436.D ;
  assign g25170 = \DFF_1437.D ;
  assign g25171 = \DFF_1438.D ;
  assign g25172 = \DFF_1433.D ;
  assign g25173 = \DFF_1511.D ;
  assign g25174 = \DFF_12.D ;
  assign g25175 = \DFF_6.D ;
  assign g25176 = \DFF_1608.D ;
  assign g25177 = \DFF_1602.D ;
  assign g25179 = \DFF_1152.D ;
  assign g25180 = \DFF_1502.D ;
  assign g25185 = \DFF_463.D ;
  assign g25189 = \DFF_813.D ;
  assign g2519 = \DFF_1329.Q ;
  assign g25191 = \DFF_1604.D ;
  assign g25194 = \DFF_1163.D ;
  assign g25197 = \DFF_1513.D ;
  assign g25199 = \DFF_14.D ;
  assign g252 = \DFF_222.Q ;
  assign g25201 = \DFF_8.D ;
  assign g25202 = \DFF_1610.D ;
  assign g25204 = \DFF_194.D ;
  assign g25206 = \DFF_195.D ;
  assign g25207 = \DFF_197.D ;
  assign g25209 = \DFF_544.D ;
  assign g25211 = \DFF_196.D ;
  assign g25212 = \DFF_198.D ;
  assign g25213 = \DFF_200.D ;
  assign g25214 = \DFF_545.D ;
  assign g25215 = \DFF_547.D ;
  assign g25217 = \DFF_894.D ;
  assign g25218 = \DFF_199.D ;
  assign g25219 = \DFF_201.D ;
  assign g2522 = \DFF_1332.Q ;
  assign g25220 = \DFF_203.D ;
  assign g25221 = \DFF_546.D ;
  assign g25222 = \DFF_548.D ;
  assign g25223 = \DFF_550.D ;
  assign g25224 = \DFF_895.D ;
  assign g25225 = \DFF_897.D ;
  assign g25227 = \DFF_1244.D ;
  assign g25228 = \DFF_202.D ;
  assign g25229 = \DFF_204.D ;
  assign g2523 = \DFF_1330.Q ;
  assign g25230 = \DFF_549.D ;
  assign g25231 = \DFF_551.D ;
  assign g25232 = \DFF_553.D ;
  assign g25233 = \DFF_896.D ;
  assign g25234 = \DFF_898.D ;
  assign g25235 = \DFF_900.D ;
  assign g25236 = \DFF_1245.D ;
  assign g25237 = \DFF_1247.D ;
  assign g25239 = \DFF_205.D ;
  assign g2524 = \DFF_1331.Q ;
  assign g25240 = \DFF_552.D ;
  assign g25241 = \DFF_554.D ;
  assign g25242 = \DFF_899.D ;
  assign g25243 = \DFF_901.D ;
  assign g25244 = \DFF_903.D ;
  assign g25245 = \DFF_1246.D ;
  assign g25246 = \DFF_1248.D ;
  assign g25247 = \DFF_1250.D ;
  assign g25248 = \DFF_555.D ;
  assign g25249 = \DFF_902.D ;
  assign g2525 = \DFF_1348.Q ;
  assign g25250 = \DFF_904.D ;
  assign g25251 = \DFF_1249.D ;
  assign g25252 = \DFF_1251.D ;
  assign g25253 = \DFF_1253.D ;
  assign g25255 = \DFF_905.D ;
  assign g25256 = \DFF_1252.D ;
  assign g25257 = \DFF_1254.D ;
  assign g25259 = \DFF_1255.D ;
  assign g2526 = \DFF_1349.Q ;
  assign g25260 = \DFF_505.D ;
  assign g25262 = \DFF_506.D ;
  assign g25263 = \DFF_855.D ;
  assign g25265 = \DFF_1600.D ;
  assign g25266 = \DFF_507.D ;
  assign g25267 = \DFF_856.D ;
  assign g25268 = \DFF_1205.D ;
  assign g2527 = \DFF_1350.Q ;
  assign g25270 = \DFF_857.D ;
  assign g25271 = \DFF_1206.D ;
  assign g25272 = \DFF_1555.D ;
  assign g25279 = \DFF_1207.D ;
  assign g2528 = \DFF_1351.Q ;
  assign g25280 = \DFF_1556.D ;
  assign g25288 = \DFF_1557.D ;
  assign g2529 = \DFF_1352.Q ;
  assign g2530 = \DFF_1433.Q ;
  assign g25327 = \DFF_236.D ;
  assign g2533 = \DFF_1434.Q ;
  assign g25336 = \DFF_586.D ;
  assign g25350 = \DFF_936.D ;
  assign g2536 = \DFF_1435.Q ;
  assign g25364 = \DFF_1286.D ;
  assign g2539 = \DFF_1441.Q ;
  assign g2540 = \DFF_1442.Q ;
  assign g25420 = \DFF_150.D ;
  assign g25421 = \DFF_150.D ;
  assign g2543 = \DFF_1443.Q ;
  assign g25435 = \DFF_151.D ;
  assign g25436 = \DFF_151.D ;
  assign g25442 = \DFF_152.D ;
  assign g25443 = \DFF_152.D ;
  assign g25450 = \DFF_107.D ;
  assign g25451 = \DFF_108.D ;
  assign g25452 = \DFF_109.D ;
  assign g2546 = \DFF_1444.Q ;
  assign g25462 = \DFF_462.D ;
  assign g25471 = \DFF_812.D ;
  assign g25488 = \DFF_1162.D ;
  assign g2549 = \DFF_1427.Q ;
  assign g25490 = \DFF_158.D ;
  assign g255 = \DFF_223.Q ;
  assign g25519 = \DFF_1512.D ;
  assign g2552 = \DFF_1436.Q ;
  assign g25520 = \DFF_159.D ;
  assign g2553 = \DFF_1437.Q ;
  assign g2554 = \DFF_1438.Q ;
  assign g2555 = \DFF_1439.Q ;
  assign g2556 = \DFF_1428.Q ;
  assign g25566 = \DFF_156.D ;
  assign g25588 = \DFF_417.D ;
  assign g2559 = \DFF_1440.Q ;
  assign g2560 = \DFF_1429.Q ;
  assign g2561 = \DFF_1430.Q ;
  assign g2562 = \DFF_1431.Q ;
  assign g2563 = \DFF_1432.Q ;
  assign g2564 = \DFF_1426.Q ;
  assign g25646 = \DFF_418.D ;
  assign g25647 = \DFF_420.D ;
  assign g2565 = \DFF_1479.Q ;
  assign g25667 = \DFF_767.D ;
  assign g2568 = \DFF_1480.Q ;
  assign g25706 = \DFF_419.D ;
  assign g25707 = \DFF_421.D ;
  assign g2571 = \DFF_1481.Q ;
  assign g25723 = \DFF_768.D ;
  assign g25724 = \DFF_770.D ;
  assign g2574 = \DFF_1452.Q ;
  assign g25744 = \DFF_1117.D ;
  assign g25762 = \DFF_1603.D ;
  assign g25763 = \DFF_1609.D ;
  assign g25770 = \DFF_422.D ;
  assign g25779 = \DFF_769.D ;
  assign g25780 = \DFF_771.D ;
  assign g25796 = \DFF_1118.D ;
  assign g25797 = \DFF_1120.D ;
  assign g258 = \DFF_227.Q ;
  assign g2580 = \DFF_1482.Q ;
  assign g2581 = \DFF_1483.Q ;
  assign g25817 = \DFF_1467.D ;
  assign g25824 = \DFF_772.D ;
  assign g25833 = \DFF_1119.D ;
  assign g25834 = \DFF_1121.D ;
  assign g2584 = \DFF_1411.Q ;
  assign g25850 = \DFF_1468.D ;
  assign g25851 = \DFF_1470.D ;
  assign g25859 = \DFF_1122.D ;
  assign g25868 = \DFF_1469.D ;
  assign g25869 = \DFF_1471.D ;
  assign g2587 = \DFF_1412.Q ;
  assign g25880 = \DFF_1472.D ;
  assign g25886 = \DFF_7.D ;
  assign g25891 = \DFF_13.D ;
  assign g25932 = \DFF_237.D ;
  assign g25935 = \DFF_587.D ;
  assign g25938 = \DFF_937.D ;
  assign g2594 = \DFF_1492.Q ;
  assign g25940 = \DFF_1287.D ;
  assign g25952 = \DFF_146.D ;
  assign g2597 = \DFF_1413.Q ;
  assign g25976 = \DFF_452.D ;
  assign g2598 = \DFF_1414.Q ;
  assign g25982 = \DFF_802.D ;
  assign g25983 = \DFF_236.D ;
  assign g25984 = \DFF_452.D ;
  assign g25985 = \DFF_417.D ;
  assign g25986 = \DFF_418.D ;
  assign g25987 = \DFF_419.D ;
  assign g25988 = \DFF_420.D ;
  assign g25989 = \DFF_421.D ;
  assign g2599 = \DFF_1493.Q ;
  assign g25990 = \DFF_422.D ;
  assign g25991 = \DFF_462.D ;
  assign g25992 = \DFF_586.D ;
  assign g25993 = \DFF_802.D ;
  assign g25994 = \DFF_767.D ;
  assign g25995 = \DFF_768.D ;
  assign g25996 = \DFF_769.D ;
  assign g25997 = \DFF_770.D ;
  assign g25998 = \DFF_771.D ;
  assign g25999 = \DFF_772.D ;
  assign g26 = \DFF_1623.Q ;
  assign g26000 = \DFF_812.D ;
  assign g26001 = \DFF_936.D ;
  assign g26002 = \DFF_1152.D ;
  assign g26003 = \DFF_1117.D ;
  assign g26004 = \DFF_1118.D ;
  assign g26005 = \DFF_1119.D ;
  assign g26006 = \DFF_1120.D ;
  assign g26007 = \DFF_1121.D ;
  assign g26008 = \DFF_1122.D ;
  assign g26009 = \DFF_1162.D ;
  assign g26010 = \DFF_1286.D ;
  assign g26011 = \DFF_1502.D ;
  assign g26012 = \DFF_1467.D ;
  assign g26013 = \DFF_1468.D ;
  assign g26014 = \DFF_1469.D ;
  assign g26015 = \DFF_1470.D ;
  assign g26016 = \DFF_1471.D ;
  assign g26017 = \DFF_1472.D ;
  assign g26018 = \DFF_1512.D ;
  assign g26019 = \DFF_7.D ;
  assign g2602 = \DFF_1445.Q ;
  assign g26020 = \DFF_13.D ;
  assign g26021 = \DFF_1603.D ;
  assign g26022 = \DFF_1609.D ;
  assign g26025 = \DFF_1347.D ;
  assign g2603 = \DFF_1494.Q ;
  assign g26031 = \DFF_1605.D ;
  assign g26037 = \DFF_9.D ;
  assign g2604 = \DFF_1495.Q ;
  assign g26048 = \DFF_1601.D ;
  assign g2605 = \DFF_1496.Q ;
  assign g2606 = \DFF_1497.Q ;
  assign g2607 = \DFF_1498.Q ;
  assign g2608 = \DFF_1499.Q ;
  assign g26086 = \DFF_237.D ;
  assign g2609 = \DFF_1446.Q ;
  assign g261 = \DFF_228.Q ;
  assign g2610 = \DFF_1500.Q ;
  assign g26102 = \DFF_587.D ;
  assign g26104 = \DFF_158.D ;
  assign g26105 = \DFF_158.D ;
  assign g26106 = \DFF_328.D ;
  assign g2611 = \DFF_1501.Q ;
  assign g26118 = \DFF_937.D ;
  assign g2612 = \DFF_1502.Q ;
  assign g26120 = \DFF_678.D ;
  assign g26125 = \DFF_1287.D ;
  assign g26130 = \DFF_1028.D ;
  assign g26135 = \DFF_159.D ;
  assign g26136 = \DFF_159.D ;
  assign g26144 = \DFF_1378.D ;
  assign g26149 = \DFF_156.D ;
  assign g2615 = \DFF_1503.Q ;
  assign g26150 = \DFF_156.D ;
  assign g26159 = \DFF_194.D ;
  assign g2616 = \DFF_1447.Q ;
  assign g26164 = \DFF_195.D ;
  assign g26165 = \DFF_197.D ;
  assign g26167 = \DFF_544.D ;
  assign g2617 = \DFF_1448.Q ;
  assign g26172 = \DFF_196.D ;
  assign g26173 = \DFF_198.D ;
  assign g26174 = \DFF_200.D ;
  assign g2618 = \DFF_1449.Q ;
  assign g26181 = \DFF_545.D ;
  assign g26182 = \DFF_547.D ;
  assign g26183 = \DFF_667.D ;
  assign g26187 = \DFF_894.D ;
  assign g26189 = \DFF_131.D ;
  assign g2619 = \DFF_1504.Q ;
  assign g26190 = \DFF_199.D ;
  assign g26191 = \DFF_201.D ;
  assign g26192 = \DFF_203.D ;
  assign g26193 = \DFF_546.D ;
  assign g26194 = \DFF_548.D ;
  assign g26195 = \DFF_550.D ;
  assign g26205 = \DFF_895.D ;
  assign g26206 = \DFF_897.D ;
  assign g26208 = \DFF_1244.D ;
  assign g26210 = \DFF_202.D ;
  assign g26211 = \DFF_204.D ;
  assign g26214 = \DFF_549.D ;
  assign g26215 = \DFF_551.D ;
  assign g26216 = \DFF_553.D ;
  assign g2622 = \DFF_1450.Q ;
  assign g26220 = \DFF_896.D ;
  assign g26221 = \DFF_898.D ;
  assign g26222 = \DFF_900.D ;
  assign g26229 = \DFF_1245.D ;
  assign g2623 = \DFF_1451.Q ;
  assign g26230 = \DFF_1247.D ;
  assign g26232 = \DFF_205.D ;
  assign g26238 = \DFF_552.D ;
  assign g26239 = \DFF_554.D ;
  assign g2624 = \DFF_1506.Q ;
  assign g26245 = \DFF_899.D ;
  assign g26246 = \DFF_901.D ;
  assign g26247 = \DFF_903.D ;
  assign g26248 = \DFF_1246.D ;
  assign g26249 = \DFF_1248.D ;
  assign g2625 = \DFF_1505.Q ;
  assign g26250 = \DFF_1250.D ;
  assign g26264 = \DFF_555.D ;
  assign g26272 = \DFF_792.D ;
  assign g26276 = \DFF_902.D ;
  assign g26277 = \DFF_904.D ;
  assign g2628 = \DFF_1409.Q ;
  assign g26280 = \DFF_1249.D ;
  assign g26281 = \DFF_1251.D ;
  assign g26282 = \DFF_1253.D ;
  assign g26294 = \DFF_463.D ;
  assign g26308 = \DFF_905.D ;
  assign g2631 = \DFF_1410.Q ;
  assign g26314 = \DFF_1252.D ;
  assign g26315 = \DFF_1254.D ;
  assign g2632 = \DFF_1453.Q ;
  assign g2633 = \DFF_1454.Q ;
  assign g26341 = \DFF_813.D ;
  assign g26349 = \DFF_1255.D ;
  assign g26354 = \DFF_1600.D ;
  assign g26355 = \DFF_1604.D ;
  assign g2636 = g2637;
  assign g26364 = \DFF_505.D ;
  assign g2638 = \DFF_1415.Q ;
  assign g26385 = \DFF_1163.D ;
  assign g2639 = \DFF_1422.Q ;
  assign g26398 = \DFF_506.D ;
  assign g264 = \DFF_229.Q ;
  assign g2640 = \DFF_1423.Q ;
  assign g26407 = \DFF_855.D ;
  assign g2641 = \DFF_1424.Q ;
  assign g2642 = \DFF_1425.Q ;
  assign g26428 = \DFF_1513.D ;
  assign g2643 = \DFF_1416.Q ;
  assign g26433 = \DFF_507.D ;
  assign g26439 = \DFF_856.D ;
  assign g2644 = \DFF_1417.Q ;
  assign g26448 = \DFF_1205.D ;
  assign g2645 = \DFF_1418.Q ;
  assign g2646 = \DFF_1419.Q ;
  assign g26465 = \DFF_857.D ;
  assign g2647 = \DFF_1420.Q ;
  assign g26471 = \DFF_1206.D ;
  assign g2648 = \DFF_1421.Q ;
  assign g26480 = \DFF_1555.D ;
  assign g26489 = \DFF_1207.D ;
  assign g2649 = \DFF_1457.Q ;
  assign g26495 = \DFF_1556.D ;
  assign g26496 = \DFF_14.D ;
  assign g2650 = \DFF_1455.Q ;
  assign g26505 = \DFF_1557.D ;
  assign g26506 = \DFF_8.D ;
  assign g26507 = \DFF_1610.D ;
  assign g2651 = \DFF_1456.Q ;
  assign g2652 = \DFF_1460.Q ;
  assign g26529 = \DFF_238.D ;
  assign g2653 = \DFF_1458.Q ;
  assign g26530 = \DFF_588.D ;
  assign g26531 = \DFF_938.D ;
  assign g26532 = \DFF_1288.D ;
  assign g26534 = \DFF_750.D ;
  assign g2654 = \DFF_1459.Q ;
  assign g26541 = \DFF_429.D ;
  assign g26545 = \DFF_430.D ;
  assign g26547 = \DFF_779.D ;
  assign g26548 = \DFF_107.D ;
  assign g2655 = \DFF_1463.Q ;
  assign g26553 = \DFF_431.D ;
  assign g26557 = \DFF_780.D ;
  assign g26559 = \DFF_1129.D ;
  assign g2656 = \DFF_1461.Q ;
  assign g26569 = \DFF_781.D ;
  assign g2657 = \DFF_1462.Q ;
  assign g26573 = \DFF_1130.D ;
  assign g26575 = \DFF_1479.D ;
  assign g26576 = \DFF_108.D ;
  assign g26577 = \DFF_144.D ;
  assign g2658 = \DFF_1466.Q ;
  assign g2659 = \DFF_1464.Q ;
  assign g26592 = \DFF_1131.D ;
  assign g26596 = \DFF_1480.D ;
  assign g2660 = \DFF_1465.Q ;
  assign g2661 = \DFF_1467.Q ;
  assign g26616 = \DFF_1481.D ;
  assign g26618 = \DFF_109.D ;
  assign g2664 = \DFF_1468.Q ;
  assign g26655 = \DFF_295.D ;
  assign g26659 = \DFF_296.D ;
  assign g26660 = \DFF_464.D ;
  assign g26661 = \DFF_645.D ;
  assign g26664 = \DFF_297.D ;
  assign g26665 = \DFF_646.D ;
  assign g26666 = \DFF_814.D ;
  assign g26667 = \DFF_995.D ;
  assign g26669 = \DFF_647.D ;
  assign g2667 = \DFF_1469.Q ;
  assign g26670 = \DFF_996.D ;
  assign g26671 = \DFF_1164.D ;
  assign g26672 = \DFF_1345.D ;
  assign g26675 = \DFF_997.D ;
  assign g26676 = \DFF_1346.D ;
  assign g26677 = \DFF_1514.D ;
  assign g26678 = \DFF_237.D ;
  assign g26679 = \DFF_194.D ;
  assign g26680 = \DFF_195.D ;
  assign g26681 = \DFF_196.D ;
  assign g26682 = \DFF_197.D ;
  assign g26683 = \DFF_198.D ;
  assign g26684 = \DFF_199.D ;
  assign g26685 = \DFF_200.D ;
  assign g26686 = \DFF_201.D ;
  assign g26687 = \DFF_202.D ;
  assign g26688 = \DFF_203.D ;
  assign g26689 = \DFF_204.D ;
  assign g26690 = \DFF_205.D ;
  assign g26691 = \DFF_463.D ;
  assign g26692 = \DFF_505.D ;
  assign g26693 = \DFF_506.D ;
  assign g26694 = \DFF_507.D ;
  assign g26695 = \DFF_587.D ;
  assign g26696 = \DFF_544.D ;
  assign g26697 = \DFF_545.D ;
  assign g26698 = \DFF_546.D ;
  assign g26699 = \DFF_547.D ;
  assign g267 = \DFF_233.Q ;
  assign g2670 = \DFF_1470.Q ;
  assign g26700 = \DFF_548.D ;
  assign g26701 = \DFF_549.D ;
  assign g26702 = \DFF_550.D ;
  assign g26703 = \DFF_551.D ;
  assign g26704 = \DFF_552.D ;
  assign g26705 = \DFF_553.D ;
  assign g26706 = \DFF_554.D ;
  assign g26707 = \DFF_555.D ;
  assign g26708 = \DFF_813.D ;
  assign g26709 = \DFF_855.D ;
  assign g26710 = \DFF_856.D ;
  assign g26711 = \DFF_857.D ;
  assign g26712 = \DFF_937.D ;
  assign g26713 = \DFF_894.D ;
  assign g26714 = \DFF_895.D ;
  assign g26715 = \DFF_896.D ;
  assign g26716 = \DFF_897.D ;
  assign g26717 = \DFF_898.D ;
  assign g26718 = \DFF_899.D ;
  assign g26719 = \DFF_900.D ;
  assign g26720 = \DFF_901.D ;
  assign g26721 = \DFF_902.D ;
  assign g26722 = \DFF_903.D ;
  assign g26723 = \DFF_904.D ;
  assign g26724 = \DFF_905.D ;
  assign g26725 = \DFF_1163.D ;
  assign g26726 = \DFF_1205.D ;
  assign g26727 = \DFF_1206.D ;
  assign g26728 = \DFF_1207.D ;
  assign g26729 = \DFF_1287.D ;
  assign g2673 = \DFF_1471.Q ;
  assign g26730 = \DFF_1244.D ;
  assign g26731 = \DFF_1245.D ;
  assign g26732 = \DFF_1246.D ;
  assign g26733 = \DFF_1247.D ;
  assign g26734 = \DFF_1248.D ;
  assign g26735 = \DFF_1249.D ;
  assign g26736 = \DFF_1250.D ;
  assign g26737 = \DFF_1251.D ;
  assign g26738 = \DFF_1252.D ;
  assign g26739 = \DFF_1253.D ;
  assign g26740 = \DFF_1254.D ;
  assign g26741 = \DFF_1255.D ;
  assign g26742 = \DFF_1513.D ;
  assign g26743 = \DFF_1555.D ;
  assign g26744 = \DFF_1556.D ;
  assign g26745 = \DFF_1557.D ;
  assign g26746 = \DFF_14.D ;
  assign g26747 = \DFF_8.D ;
  assign g26748 = \DFF_1600.D ;
  assign g26749 = \DFF_1610.D ;
  assign g26750 = \DFF_1604.D ;
  assign g26751 = \DFF_107.D ;
  assign g26752 = \DFF_108.D ;
  assign g26753 = \DFF_109.D ;
  assign g2676 = \DFF_1472.Q ;
  assign g26776 = \DFF_465.D ;
  assign g26781 = \DFF_815.D ;
  assign g26786 = \DFF_1606.D ;
  assign g26789 = \DFF_1165.D ;
  assign g2679 = \DFF_1476.Q ;
  assign g26795 = \DFF_1515.D ;
  assign g26798 = \DFF_10.D ;
  assign g26803 = \DFF_274.D ;
  assign g26804 = \DFF_275.D ;
  assign g26805 = \DFF_277.D ;
  assign g26806 = \DFF_624.D ;
  assign g26807 = \DFF_276.D ;
  assign g26808 = \DFF_278.D ;
  assign g26809 = \DFF_625.D ;
  assign g26810 = \DFF_627.D ;
  assign g26811 = \DFF_974.D ;
  assign g26812 = \DFF_279.D ;
  assign g26813 = \DFF_626.D ;
  assign g26814 = \DFF_628.D ;
  assign g26815 = \DFF_975.D ;
  assign g26816 = \DFF_977.D ;
  assign g26817 = \DFF_1324.D ;
  assign g26818 = \DFF_629.D ;
  assign g26819 = \DFF_750.D ;
  assign g2682 = \DFF_1477.Q ;
  assign g26820 = \DFF_976.D ;
  assign g26821 = \DFF_978.D ;
  assign g26822 = \DFF_1325.D ;
  assign g26823 = \DFF_1327.D ;
  assign g26824 = \DFF_979.D ;
  assign g26825 = \DFF_1326.D ;
  assign g26826 = \DFF_1328.D ;
  assign g26827 = \DFF_1329.D ;
  assign g26828 = \DFF_429.D ;
  assign g26830 = \DFF_430.D ;
  assign g26831 = \DFF_779.D ;
  assign g26832 = \DFF_431.D ;
  assign g26834 = \DFF_780.D ;
  assign g26836 = \DFF_1129.D ;
  assign g26840 = \DFF_781.D ;
  assign g26843 = \DFF_1130.D ;
  assign g26844 = \DFF_1479.D ;
  assign g2685 = \DFF_1478.Q ;
  assign g26850 = \DFF_1131.D ;
  assign g26852 = \DFF_1480.D ;
  assign g26858 = \DFF_1481.D ;
  assign g26864 = \DFF_238.D ;
  assign g26868 = \DFF_588.D ;
  assign g26872 = \DFF_295.D ;
  assign g26875 = \DFF_938.D ;
  assign g26876 = \DFF_296.D ;
  assign g2688 = \DFF_1473.Q ;
  assign g26881 = \DFF_645.D ;
  assign g26883 = \DFF_1288.D ;
  assign g26884 = \DFF_297.D ;
  assign g26886 = \DFF_646.D ;
  assign g26890 = \DFF_995.D ;
  assign g26895 = \DFF_647.D ;
  assign g26896 = \DFF_996.D ;
  assign g26900 = \DFF_1345.D ;
  assign g26909 = \DFF_997.D ;
  assign g2691 = \DFF_1474.Q ;
  assign g26910 = \DFF_1346.D ;
  assign g26921 = \DFF_1347.D ;
  assign g2694 = \DFF_1475.Q ;
  assign g26953 = \DFF_464.D ;
  assign g26954 = \DFF_150.D ;
  assign g26956 = \DFF_814.D ;
  assign g26957 = \DFF_151.D ;
  assign g26959 = \DFF_1164.D ;
  assign g26960 = \DFF_152.D ;
  assign g26964 = \DFF_1514.D ;
  assign g2697 = \DFF_1504.Q ;
  assign g26974 = \DFF_157.D ;
  assign g26983 = \DFF_792.D ;
  assign g27 = \DFF_1618.Q ;
  assign g270 = \DFF_234.Q ;
  assign g2700 = \DFF_1505.Q ;
  assign g2703 = \DFF_1506.Q ;
  assign g2704 = \DFF_1507.Q ;
  assign g2707 = \DFF_1510.Q ;
  assign g27075 = \DFF_1601.D ;
  assign g27102 = \DFF_1605.D ;
  assign g27116 = \DFF_9.D ;
  assign g27120 = \DFF_239.D ;
  assign g27123 = \DFF_589.D ;
  assign g27126 = \DFF_750.D ;
  assign g27129 = \DFF_939.D ;
  assign g27131 = \DFF_1289.D ;
  assign g27132 = \DFF_667.D ;
  assign g2714 = \DFF_1509.Q ;
  assign g27140 = \DFF_141.D ;
  assign g27145 = \DFF_328.D ;
  assign g27150 = \DFF_678.D ;
  assign g27156 = \DFF_792.D ;
  assign g27158 = \DFF_1028.D ;
  assign g27166 = \DFF_1378.D ;
  assign g27168 = \DFF_131.D ;
  assign g27183 = \DFF_667.D ;
  assign g27189 = \DFF_238.D ;
  assign g27190 = \DFF_328.D ;
  assign g27191 = \DFF_295.D ;
  assign g27192 = \DFF_296.D ;
  assign g27193 = \DFF_297.D ;
  assign g27194 = \DFF_429.D ;
  assign g27195 = \DFF_430.D ;
  assign g27196 = \DFF_431.D ;
  assign g27197 = \DFF_464.D ;
  assign g27198 = \DFF_588.D ;
  assign g27199 = \DFF_678.D ;
  assign g2720 = \DFF_1512.Q ;
  assign g27200 = \DFF_667.D ;
  assign g27206 = \DFF_645.D ;
  assign g27207 = \DFF_646.D ;
  assign g27208 = \DFF_647.D ;
  assign g27209 = \DFF_779.D ;
  assign g27210 = \DFF_780.D ;
  assign g27211 = \DFF_781.D ;
  assign g27212 = \DFF_792.D ;
  assign g27217 = \DFF_750.D ;
  assign g27218 = \DFF_814.D ;
  assign g27219 = \DFF_938.D ;
  assign g27220 = \DFF_1028.D ;
  assign g27221 = \DFF_995.D ;
  assign g27222 = \DFF_996.D ;
  assign g27223 = \DFF_997.D ;
  assign g27224 = \DFF_1129.D ;
  assign g27225 = \DFF_1130.D ;
  assign g27226 = \DFF_1131.D ;
  assign g27227 = \DFF_1164.D ;
  assign g27228 = \DFF_1288.D ;
  assign g27229 = \DFF_1378.D ;
  assign g27230 = \DFF_1345.D ;
  assign g27231 = \DFF_1346.D ;
  assign g27232 = \DFF_1347.D ;
  assign g27233 = \DFF_1479.D ;
  assign g27234 = \DFF_1480.D ;
  assign g27235 = \DFF_1481.D ;
  assign g27236 = \DFF_1514.D ;
  assign g27237 = \DFF_9.D ;
  assign g27238 = \DFF_1601.D ;
  assign g27239 = \DFF_1605.D ;
  assign g27243 = \DFF_1516.D ;
  assign g27253 = \DFF_253.D ;
  assign g27255 = \DFF_254.D ;
  assign g27256 = \DFF_256.D ;
  assign g27257 = \DFF_603.D ;
  assign g27258 = \DFF_255.D ;
  assign g27259 = \DFF_257.D ;
  assign g27260 = \DFF_259.D ;
  assign g27261 = \DFF_405.D ;
  assign g27262 = \DFF_604.D ;
  assign g27263 = \DFF_606.D ;
  assign g27264 = \DFF_953.D ;
  assign g27265 = \DFF_258.D ;
  assign g27266 = \DFF_260.D ;
  assign g27267 = \DFF_262.D ;
  assign g27268 = \DFF_406.D ;
  assign g27269 = \DFF_408.D ;
  assign g2727 = \DFF_1511.Q ;
  assign g27270 = \DFF_605.D ;
  assign g27271 = \DFF_607.D ;
  assign g27272 = \DFF_609.D ;
  assign g27273 = \DFF_755.D ;
  assign g27274 = \DFF_954.D ;
  assign g27275 = \DFF_956.D ;
  assign g27276 = \DFF_1303.D ;
  assign g27277 = \DFF_261.D ;
  assign g27278 = \DFF_263.D ;
  assign g27279 = \DFF_407.D ;
  assign g27280 = \DFF_409.D ;
  assign g27281 = \DFF_411.D ;
  assign g27282 = \DFF_608.D ;
  assign g27283 = \DFF_610.D ;
  assign g27284 = \DFF_612.D ;
  assign g27285 = \DFF_756.D ;
  assign g27286 = \DFF_758.D ;
  assign g27287 = \DFF_955.D ;
  assign g27288 = \DFF_957.D ;
  assign g27289 = \DFF_959.D ;
  assign g27290 = \DFF_1105.D ;
  assign g27291 = \DFF_1304.D ;
  assign g27292 = \DFF_1306.D ;
  assign g27293 = \DFF_264.D ;
  assign g27294 = \DFF_410.D ;
  assign g27295 = \DFF_412.D ;
  assign g27296 = \DFF_414.D ;
  assign g27297 = \DFF_611.D ;
  assign g27298 = \DFF_613.D ;
  assign g27299 = \DFF_757.D ;
  assign g273 = \DFF_235.Q ;
  assign g27300 = \DFF_759.D ;
  assign g27301 = \DFF_761.D ;
  assign g27302 = \DFF_958.D ;
  assign g27303 = \DFF_960.D ;
  assign g27304 = \DFF_962.D ;
  assign g27305 = \DFF_1106.D ;
  assign g27306 = \DFF_1108.D ;
  assign g27307 = \DFF_1305.D ;
  assign g27308 = \DFF_1307.D ;
  assign g27309 = \DFF_1309.D ;
  assign g27310 = \DFF_1455.D ;
  assign g27311 = \DFF_413.D ;
  assign g27312 = \DFF_415.D ;
  assign g27313 = \DFF_614.D ;
  assign g27314 = \DFF_760.D ;
  assign g27315 = \DFF_762.D ;
  assign g27316 = \DFF_764.D ;
  assign g27317 = \DFF_961.D ;
  assign g27318 = \DFF_963.D ;
  assign g27319 = \DFF_1107.D ;
  assign g27320 = \DFF_1109.D ;
  assign g27321 = \DFF_1111.D ;
  assign g27322 = \DFF_1308.D ;
  assign g27323 = \DFF_1310.D ;
  assign g27324 = \DFF_1312.D ;
  assign g27325 = \DFF_1456.D ;
  assign g27326 = \DFF_1458.D ;
  assign g27327 = \DFF_416.D ;
  assign g27328 = \DFF_763.D ;
  assign g27329 = \DFF_765.D ;
  assign g2733 = \DFF_1508.Q ;
  assign g27330 = \DFF_964.D ;
  assign g27331 = \DFF_1110.D ;
  assign g27332 = \DFF_1112.D ;
  assign g27333 = \DFF_1114.D ;
  assign g27334 = \DFF_1311.D ;
  assign g27335 = \DFF_1313.D ;
  assign g27336 = \DFF_1457.D ;
  assign g27337 = \DFF_1459.D ;
  assign g27338 = \DFF_1461.D ;
  assign g27339 = \DFF_766.D ;
  assign g2734 = \DFF_1513.Q ;
  assign g27340 = \DFF_1113.D ;
  assign g27341 = \DFF_1115.D ;
  assign g27342 = \DFF_1314.D ;
  assign g27343 = \DFF_1460.D ;
  assign g27344 = \DFF_1462.D ;
  assign g27345 = \DFF_1464.D ;
  assign g27346 = \DFF_1116.D ;
  assign g27347 = \DFF_1463.D ;
  assign g27348 = \DFF_1465.D ;
  assign g27353 = \DFF_239.D ;
  assign g27354 = \DFF_1466.D ;
  assign g27357 = \DFF_589.D ;
  assign g27360 = \DFF_939.D ;
  assign g27366 = \DFF_1289.D ;
  assign g27380 = \DFF_157.D ;
  assign g27381 = \DFF_157.D ;
  assign g27383 = \DFF_158.D ;
  assign g27384 = \DFF_159.D ;
  assign g27385 = \DFF_131.D ;
  assign g27386 = \DFF_156.D ;
  assign g2740 = \DFF_1515.Q ;
  assign g2746 = \DFF_1514.Q ;
  assign g27463 = \DFF_274.D ;
  assign g27479 = \DFF_275.D ;
  assign g27480 = \DFF_277.D ;
  assign g27483 = \DFF_624.D ;
  assign g27493 = \DFF_276.D ;
  assign g27494 = \DFF_278.D ;
  assign g27497 = \DFF_465.D ;
  assign g27502 = \DFF_625.D ;
  assign g27503 = \DFF_627.D ;
  assign g27505 = \DFF_974.D ;
  assign g27508 = \DFF_279.D ;
  assign g27514 = \DFF_626.D ;
  assign g27515 = \DFF_628.D ;
  assign g27517 = \DFF_815.D ;
  assign g27522 = \DFF_975.D ;
  assign g27523 = \DFF_977.D ;
  assign g27525 = \DFF_1324.D ;
  assign g27526 = \DFF_1606.D ;
  assign g2753 = \DFF_1516.Q ;
  assign g27533 = \DFF_629.D ;
  assign g27539 = \DFF_976.D ;
  assign g27540 = \DFF_978.D ;
  assign g27542 = \DFF_1165.D ;
  assign g27547 = \DFF_1325.D ;
  assign g27548 = \DFF_1327.D ;
  assign g27553 = \DFF_979.D ;
  assign g27559 = \DFF_1326.D ;
  assign g27560 = \DFF_1328.D ;
  assign g27562 = \DFF_1515.D ;
  assign g27569 = \DFF_1329.D ;
  assign g27586 = \DFF_10.D ;
  assign g27589 = \DFF_146.D ;
  assign g27594 = \DFF_240.D ;
  assign g276 = \DFF_1427.Q ;
  assign g2760 = \DFF_1517.Q ;
  assign g27603 = \DFF_590.D ;
  assign g27612 = \DFF_940.D ;
  assign g27621 = \DFF_1290.D ;
  assign g2766 = \DFF_1518.Q ;
  assign g27662 = \DFF_152.D ;
  assign g27667 = \DFF_151.D ;
  assign g27672 = \DFF_466.D ;
  assign g27674 = \DFF_150.D ;
  assign g27678 = \DFF_816.D ;
  assign g27682 = \DFF_1166.D ;
  assign g27683 = \DFF_239.D ;
  assign g27684 = \DFF_274.D ;
  assign g27685 = \DFF_275.D ;
  assign g27686 = \DFF_276.D ;
  assign g27687 = \DFF_277.D ;
  assign g27688 = \DFF_278.D ;
  assign g27689 = \DFF_279.D ;
  assign g27690 = \DFF_465.D ;
  assign g27691 = \DFF_589.D ;
  assign g27692 = \DFF_624.D ;
  assign g27693 = \DFF_625.D ;
  assign g27694 = \DFF_626.D ;
  assign g27695 = \DFF_627.D ;
  assign g27696 = \DFF_628.D ;
  assign g27697 = \DFF_629.D ;
  assign g27698 = \DFF_815.D ;
  assign g27699 = \DFF_939.D ;
  assign g27700 = \DFF_974.D ;
  assign g27701 = \DFF_975.D ;
  assign g27702 = \DFF_976.D ;
  assign g27703 = \DFF_977.D ;
  assign g27704 = \DFF_978.D ;
  assign g27705 = \DFF_979.D ;
  assign g27706 = \DFF_1165.D ;
  assign g27707 = \DFF_1289.D ;
  assign g27708 = \DFF_1324.D ;
  assign g27709 = \DFF_1325.D ;
  assign g27710 = \DFF_1326.D ;
  assign g27711 = \DFF_1327.D ;
  assign g27712 = \DFF_1328.D ;
  assign g27713 = \DFF_1329.D ;
  assign g27714 = \DFF_1515.D ;
  assign g27715 = \DFF_10.D ;
  assign g27716 = \DFF_1606.D ;
  assign g27717 = \DFF_131.D ;
  assign g27718 = \DFF_817.D ;
  assign g2772 = \DFF_1521.Q ;
  assign g27722 = \DFF_1167.D ;
  assign g27724 = \DFF_1517.D ;
  assign g2773 = \DFF_1519.Q ;
  assign g2774 = \DFF_1520.Q ;
  assign g2775 = \DFF_1524.Q ;
  assign g27759 = \DFF_280.D ;
  assign g2776 = \DFF_1522.Q ;
  assign g27760 = \DFF_281.D ;
  assign g27761 = \DFF_630.D ;
  assign g27762 = \DFF_282.D ;
  assign g27763 = \DFF_631.D ;
  assign g27764 = \DFF_980.D ;
  assign g27765 = \DFF_632.D ;
  assign g27766 = \DFF_981.D ;
  assign g27767 = \DFF_1330.D ;
  assign g27768 = \DFF_982.D ;
  assign g27769 = \DFF_1331.D ;
  assign g2777 = \DFF_1523.Q ;
  assign g27771 = \DFF_1332.D ;
  assign g2778 = \DFF_1527.Q ;
  assign g27784 = \DFF_152.D ;
  assign g27785 = \DFF_146.D ;
  assign g27786 = \DFF_240.D ;
  assign g2779 = \DFF_1525.Q ;
  assign g27791 = \DFF_151.D ;
  assign g27792 = \DFF_152.D ;
  assign g27793 = \DFF_590.D ;
  assign g27797 = \DFF_150.D ;
  assign g27799 = \DFF_940.D ;
  assign g2780 = \DFF_1526.Q ;
  assign g27800 = \DFF_150.D ;
  assign g27805 = \DFF_1290.D ;
  assign g2781 = \DFF_1530.Q ;
  assign g2782 = \DFF_1528.Q ;
  assign g2783 = \DFF_1529.Q ;
  assign g2784 = \DFF_1533.Q ;
  assign g2785 = \DFF_1531.Q ;
  assign g2786 = \DFF_1532.Q ;
  assign g2787 = \DFF_1536.Q ;
  assign g2788 = \DFF_1534.Q ;
  assign g2789 = \DFF_1535.Q ;
  assign g279 = \DFF_303.Q ;
  assign g2790 = \DFF_1539.Q ;
  assign g27903 = \DFF_152.D ;
  assign g27905 = \DFF_466.D ;
  assign g27907 = \DFF_151.D ;
  assign g2791 = \DFF_1537.Q ;
  assign g27910 = \DFF_816.D ;
  assign g27912 = \DFF_150.D ;
  assign g27918 = \DFF_1166.D ;
  assign g2792 = \DFF_1538.Q ;
  assign g27927 = \DFF_1516.D ;
  assign g2793 = \DFF_1542.Q ;
  assign g2794 = \DFF_1540.Q ;
  assign g2795 = \DFF_1541.Q ;
  assign g27955 = \DFF_253.D ;
  assign g2796 = \DFF_1545.Q ;
  assign g2797 = \DFF_1543.Q ;
  assign g27971 = \DFF_254.D ;
  assign g27972 = \DFF_256.D ;
  assign g27976 = \DFF_603.D ;
  assign g2798 = \DFF_1544.Q ;
  assign g27986 = \DFF_255.D ;
  assign g27987 = \DFF_257.D ;
  assign g27988 = \DFF_259.D ;
  assign g27989 = \DFF_405.D ;
  assign g2799 = \DFF_1548.Q ;
  assign g27992 = \DFF_604.D ;
  assign g27993 = \DFF_606.D ;
  assign g27998 = \DFF_953.D ;
  assign g280 = \DFF_304.Q ;
  assign g2800 = \DFF_1546.Q ;
  assign g28003 = \DFF_258.D ;
  assign g28004 = \DFF_260.D ;
  assign g28005 = \DFF_262.D ;
  assign g28006 = \DFF_406.D ;
  assign g28007 = \DFF_408.D ;
  assign g2801 = \DFF_1547.Q ;
  assign g28010 = \DFF_605.D ;
  assign g28011 = \DFF_607.D ;
  assign g28012 = \DFF_609.D ;
  assign g28013 = \DFF_755.D ;
  assign g28016 = \DFF_954.D ;
  assign g28017 = \DFF_956.D ;
  assign g2802 = \DFF_1551.Q ;
  assign g28021 = \DFF_1303.D ;
  assign g28022 = \DFF_261.D ;
  assign g28023 = \DFF_263.D ;
  assign g28024 = \DFF_407.D ;
  assign g28025 = \DFF_409.D ;
  assign g28026 = \DFF_411.D ;
  assign g2803 = \DFF_1549.Q ;
  assign g28030 = \DFF_608.D ;
  assign g28031 = \DFF_610.D ;
  assign g28032 = \DFF_612.D ;
  assign g28033 = \DFF_756.D ;
  assign g28034 = \DFF_758.D ;
  assign g28037 = \DFF_955.D ;
  assign g28038 = \DFF_957.D ;
  assign g28039 = \DFF_959.D ;
  assign g2804 = \DFF_1550.Q ;
  assign g28040 = \DFF_1105.D ;
  assign g28043 = \DFF_1304.D ;
  assign g28044 = \DFF_1306.D ;
  assign g28045 = \DFF_264.D ;
  assign g28047 = \DFF_410.D ;
  assign g28048 = \DFF_412.D ;
  assign g28049 = \DFF_414.D ;
  assign g2805 = \DFF_1554.Q ;
  assign g28052 = \DFF_611.D ;
  assign g28053 = \DFF_613.D ;
  assign g28054 = \DFF_757.D ;
  assign g28055 = \DFF_759.D ;
  assign g28056 = \DFF_761.D ;
  assign g2806 = \DFF_1552.Q ;
  assign g28060 = \DFF_958.D ;
  assign g28061 = \DFF_960.D ;
  assign g28062 = \DFF_962.D ;
  assign g28063 = \DFF_1106.D ;
  assign g28064 = \DFF_1108.D ;
  assign g28067 = \DFF_1305.D ;
  assign g28068 = \DFF_1307.D ;
  assign g28069 = \DFF_1309.D ;
  assign g2807 = \DFF_1553.Q ;
  assign g28070 = \DFF_1455.D ;
  assign g28071 = \DFF_413.D ;
  assign g28072 = \DFF_415.D ;
  assign g28074 = \DFF_614.D ;
  assign g28076 = \DFF_760.D ;
  assign g28077 = \DFF_762.D ;
  assign g28078 = \DFF_764.D ;
  assign g2808 = \DFF_1557.Q ;
  assign g28081 = \DFF_961.D ;
  assign g28082 = \DFF_963.D ;
  assign g28083 = \DFF_1107.D ;
  assign g28084 = \DFF_1109.D ;
  assign g28085 = \DFF_1111.D ;
  assign g28089 = \DFF_1308.D ;
  assign g2809 = \DFF_1555.Q ;
  assign g28090 = \DFF_1310.D ;
  assign g28091 = \DFF_1312.D ;
  assign g28092 = \DFF_1456.D ;
  assign g28093 = \DFF_1458.D ;
  assign g28095 = \DFF_416.D ;
  assign g28096 = \DFF_763.D ;
  assign g28097 = \DFF_765.D ;
  assign g28099 = \DFF_964.D ;
  assign g281 = \DFF_305.Q ;
  assign g2810 = \DFF_1556.Q ;
  assign g28101 = \DFF_1110.D ;
  assign g28102 = \DFF_1112.D ;
  assign g28103 = \DFF_1114.D ;
  assign g28106 = \DFF_1311.D ;
  assign g28107 = \DFF_1313.D ;
  assign g28108 = \DFF_1457.D ;
  assign g28109 = \DFF_1459.D ;
  assign g2811 = \DFF_1560.Q ;
  assign g28110 = \DFF_1461.D ;
  assign g28113 = \DFF_766.D ;
  assign g28114 = \DFF_1113.D ;
  assign g28115 = \DFF_1115.D ;
  assign g28117 = \DFF_1314.D ;
  assign g28119 = \DFF_1460.D ;
  assign g2812 = \DFF_1558.Q ;
  assign g28120 = \DFF_1462.D ;
  assign g28121 = \DFF_1464.D ;
  assign g28124 = \DFF_1116.D ;
  assign g28125 = \DFF_1463.D ;
  assign g28126 = \DFF_1465.D ;
  assign g2813 = \DFF_1559.Q ;
  assign g28132 = \DFF_1466.D ;
  assign g2814 = \DFF_17.Q ;
  assign g28145 = \DFF_241.D ;
  assign g28146 = \DFF_591.D ;
  assign g28147 = \DFF_941.D ;
  assign g28148 = \DFF_1291.D ;
  assign g28149 = \DFF_144.D ;
  assign g28151 = \DFF_160.D ;
  assign g2817 = \DFF_1.Q ;
  assign g28179 = \DFF_158.D ;
  assign g2818 = \DFF_55.Q ;
  assign g28194 = \DFF_156.D ;
  assign g28199 = \DFF_467.D ;
  assign g282 = \DFF_306.Q ;
  assign g28200 = \DFF_159.D ;
  assign g28206 = \DFF_240.D ;
  assign g28207 = \DFF_253.D ;
  assign g28208 = \DFF_254.D ;
  assign g28209 = \DFF_255.D ;
  assign g2821 = \DFF_57.Q ;
  assign g28210 = \DFF_256.D ;
  assign g28211 = \DFF_257.D ;
  assign g28212 = \DFF_258.D ;
  assign g28213 = \DFF_259.D ;
  assign g28214 = \DFF_260.D ;
  assign g28215 = \DFF_261.D ;
  assign g28216 = \DFF_262.D ;
  assign g28217 = \DFF_263.D ;
  assign g28218 = \DFF_264.D ;
  assign g28219 = \DFF_405.D ;
  assign g28220 = \DFF_406.D ;
  assign g28221 = \DFF_407.D ;
  assign g28222 = \DFF_408.D ;
  assign g28223 = \DFF_409.D ;
  assign g28224 = \DFF_410.D ;
  assign g28225 = \DFF_411.D ;
  assign g28226 = \DFF_412.D ;
  assign g28227 = \DFF_413.D ;
  assign g28228 = \DFF_414.D ;
  assign g28229 = \DFF_415.D ;
  assign g28230 = \DFF_416.D ;
  assign g28231 = \DFF_466.D ;
  assign g28232 = \DFF_590.D ;
  assign g28233 = \DFF_603.D ;
  assign g28234 = \DFF_604.D ;
  assign g28235 = \DFF_605.D ;
  assign g28236 = \DFF_606.D ;
  assign g28237 = \DFF_607.D ;
  assign g28238 = \DFF_608.D ;
  assign g28239 = \DFF_609.D ;
  assign g2824 = \DFF_59.Q ;
  assign g28240 = \DFF_610.D ;
  assign g28241 = \DFF_611.D ;
  assign g28242 = \DFF_612.D ;
  assign g28243 = \DFF_613.D ;
  assign g28244 = \DFF_614.D ;
  assign g28245 = \DFF_755.D ;
  assign g28246 = \DFF_756.D ;
  assign g28247 = \DFF_757.D ;
  assign g28248 = \DFF_758.D ;
  assign g28249 = \DFF_759.D ;
  assign g28250 = \DFF_760.D ;
  assign g28251 = \DFF_761.D ;
  assign g28252 = \DFF_762.D ;
  assign g28253 = \DFF_763.D ;
  assign g28254 = \DFF_764.D ;
  assign g28255 = \DFF_765.D ;
  assign g28256 = \DFF_766.D ;
  assign g28257 = \DFF_816.D ;
  assign g28258 = \DFF_940.D ;
  assign g28259 = \DFF_953.D ;
  assign g28260 = \DFF_954.D ;
  assign g28261 = \DFF_955.D ;
  assign g28262 = \DFF_956.D ;
  assign g28263 = \DFF_957.D ;
  assign g28264 = \DFF_958.D ;
  assign g28265 = \DFF_959.D ;
  assign g28266 = \DFF_960.D ;
  assign g28267 = \DFF_961.D ;
  assign g28268 = \DFF_962.D ;
  assign g28269 = \DFF_963.D ;
  assign g2827 = \DFF_61.Q ;
  assign g28270 = \DFF_964.D ;
  assign g28271 = \DFF_1105.D ;
  assign g28272 = \DFF_1106.D ;
  assign g28273 = \DFF_1107.D ;
  assign g28274 = \DFF_1108.D ;
  assign g28275 = \DFF_1109.D ;
  assign g28276 = \DFF_1110.D ;
  assign g28277 = \DFF_1111.D ;
  assign g28278 = \DFF_1112.D ;
  assign g28279 = \DFF_1113.D ;
  assign g28280 = \DFF_1114.D ;
  assign g28281 = \DFF_1115.D ;
  assign g28282 = \DFF_1116.D ;
  assign g28283 = \DFF_1166.D ;
  assign g28284 = \DFF_1290.D ;
  assign g28285 = \DFF_1303.D ;
  assign g28286 = \DFF_1304.D ;
  assign g28287 = \DFF_1305.D ;
  assign g28288 = \DFF_1306.D ;
  assign g28289 = \DFF_1307.D ;
  assign g28290 = \DFF_1308.D ;
  assign g28291 = \DFF_1309.D ;
  assign g28292 = \DFF_1310.D ;
  assign g28293 = \DFF_1311.D ;
  assign g28294 = \DFF_1312.D ;
  assign g28295 = \DFF_1313.D ;
  assign g28296 = \DFF_1314.D ;
  assign g28297 = \DFF_1455.D ;
  assign g28298 = \DFF_1456.D ;
  assign g28299 = \DFF_1457.D ;
  assign g283 = \DFF_307.Q ;
  assign g2830 = \DFF_63.Q ;
  assign g28300 = \DFF_1458.D ;
  assign g28301 = \DFF_1459.D ;
  assign g28302 = \DFF_1460.D ;
  assign g28303 = \DFF_1461.D ;
  assign g28304 = \DFF_1462.D ;
  assign g28305 = \DFF_1463.D ;
  assign g28306 = \DFF_1464.D ;
  assign g28307 = \DFF_1465.D ;
  assign g28308 = \DFF_1466.D ;
  assign g28309 = \DFF_1516.D ;
  assign g28310 = \DFF_152.D ;
  assign g28311 = \DFF_151.D ;
  assign g28312 = \DFF_150.D ;
  assign g28313 = \DFF_146.D ;
  assign g28314 = \DFF_152.D ;
  assign g28315 = \DFF_150.D ;
  assign g28316 = \DFF_152.D ;
  assign g28317 = \DFF_151.D ;
  assign g28318 = \DFF_150.D ;
  assign g28321 = \DFF_818.D ;
  assign g28325 = \DFF_1168.D ;
  assign g28328 = \DFF_1518.D ;
  assign g2833 = \DFF_65.Q ;
  assign g28341 = \DFF_156.D ;
  assign g28342 = \DFF_426.D ;
  assign g28343 = \DFF_159.D ;
  assign g28344 = \DFF_427.D ;
  assign g28345 = \DFF_423.D ;
  assign g28346 = \DFF_776.D ;
  assign g28347 = \DFF_158.D ;
  assign g28348 = \DFF_428.D ;
  assign g28349 = \DFF_424.D ;
  assign g28350 = \DFF_777.D ;
  assign g28351 = \DFF_773.D ;
  assign g28352 = \DFF_1126.D ;
  assign g28353 = \DFF_425.D ;
  assign g28354 = \DFF_778.D ;
  assign g28355 = \DFF_774.D ;
  assign g28356 = \DFF_1127.D ;
  assign g28357 = \DFF_1123.D ;
  assign g28358 = \DFF_1476.D ;
  assign g28359 = \DFF_159.D ;
  assign g2836 = \DFF_67.Q ;
  assign g28360 = \DFF_775.D ;
  assign g28361 = \DFF_1128.D ;
  assign g28362 = \DFF_1124.D ;
  assign g28363 = \DFF_1477.D ;
  assign g28364 = \DFF_1473.D ;
  assign g28365 = \DFF_158.D ;
  assign g28366 = \DFF_1125.D ;
  assign g28367 = \DFF_1478.D ;
  assign g28368 = \DFF_1474.D ;
  assign g28369 = \DFF_159.D ;
  assign g28370 = \DFF_241.D ;
  assign g28371 = \DFF_1475.D ;
  assign g28372 = \DFF_158.D ;
  assign g28374 = \DFF_591.D ;
  assign g28375 = \DFF_158.D ;
  assign g28377 = \DFF_941.D ;
  assign g28382 = \DFF_1291.D ;
  assign g2839 = \DFF_69.Q ;
  assign g28390 = \DFF_144.D ;
  assign g28393 = \DFF_156.D ;
  assign g28395 = \DFF_156.D ;
  assign g284 = \DFF_308.Q ;
  assign g28419 = \DFF_157.D ;
  assign g2842 = \DFF_71.Q ;
  assign g28420 = \DFF_110.D ;
  assign g28421 = \DFF_111.D ;
  assign g28425 = \DFF_112.D ;
  assign g28432 = \DFF_467.D ;
  assign g28437 = \DFF_156.D ;
  assign g28443 = \DFF_817.D ;
  assign g28447 = \DFF_159.D ;
  assign g2845 = \DFF_73.Q ;
  assign g28455 = \DFF_1167.D ;
  assign g28458 = \DFF_158.D ;
  assign g28467 = \DFF_1517.D ;
  assign g2848 = \DFF_75.Q ;
  assign g28498 = \DFF_280.D ;
  assign g285 = \DFF_309.Q ;
  assign g2851 = \DFF_77.Q ;
  assign g28524 = \DFF_281.D ;
  assign g28526 = \DFF_630.D ;
  assign g28527 = \DFF_282.D ;
  assign g2854 = \DFF_79.Q ;
  assign g28552 = \DFF_631.D ;
  assign g28553 = \DFF_980.D ;
  assign g28555 = \DFF_632.D ;
  assign g2857 = \DFF_82.Q ;
  assign g28579 = \DFF_981.D ;
  assign g2858 = \DFF_81.Q ;
  assign g28580 = \DFF_1330.D ;
  assign g28583 = \DFF_982.D ;
  assign g286 = \DFF_310.Q ;
  assign g28607 = \DFF_1331.D ;
  assign g2861 = \DFF_47.Q ;
  assign g28611 = \DFF_1332.D ;
  assign g28634 = \DFF_242.D ;
  assign g28635 = \DFF_592.D ;
  assign g28636 = \DFF_942.D ;
  assign g28637 = \DFF_1292.D ;
  assign g28638 = \DFF_141.D ;
  assign g2864 = \DFF_49.Q ;
  assign g28668 = \DFF_468.D ;
  assign g2867 = \DFF_51.Q ;
  assign g28673 = \DFF_241.D ;
  assign g28674 = \DFF_280.D ;
  assign g28675 = \DFF_281.D ;
  assign g28676 = \DFF_282.D ;
  assign g28677 = \DFF_467.D ;
  assign g28678 = \DFF_591.D ;
  assign g28679 = \DFF_630.D ;
  assign g28680 = \DFF_631.D ;
  assign g28681 = \DFF_632.D ;
  assign g28682 = \DFF_817.D ;
  assign g28683 = \DFF_941.D ;
  assign g28684 = \DFF_980.D ;
  assign g28685 = \DFF_981.D ;
  assign g28686 = \DFF_982.D ;
  assign g28687 = \DFF_1167.D ;
  assign g28688 = \DFF_1291.D ;
  assign g28689 = \DFF_1330.D ;
  assign g28690 = \DFF_1331.D ;
  assign g28691 = \DFF_1332.D ;
  assign g28692 = \DFF_1517.D ;
  assign g28693 = \DFF_156.D ;
  assign g28694 = \DFF_159.D ;
  assign g28695 = \DFF_158.D ;
  assign g28696 = \DFF_144.D ;
  assign g28697 = \DFF_156.D ;
  assign g28698 = \DFF_158.D ;
  assign g28699 = \DFF_156.D ;
  assign g287 = \DFF_311.Q ;
  assign g2870 = \DFF_53.Q ;
  assign g28700 = \DFF_159.D ;
  assign g28701 = \DFF_158.D ;
  assign g28702 = \DFF_159.D ;
  assign g28703 = \DFF_158.D ;
  assign g28704 = \DFF_156.D ;
  assign g28705 = \DFF_159.D ;
  assign g28706 = \DFF_158.D ;
  assign g28720 = \DFF_1571.D ;
  assign g28721 = \DFF_1570.D ;
  assign g28723 = \DFF_1569.D ;
  assign g28725 = \DFF_1568.D ;
  assign g28727 = \DFF_1567.D ;
  assign g2873 = \DFF_64.Q ;
  assign g28730 = \DFF_1566.D ;
  assign g28732 = \DFF_265.D ;
  assign g28734 = \DFF_1565.D ;
  assign g28735 = \DFF_266.D ;
  assign g28736 = \DFF_271.D ;
  assign g28738 = \DFF_615.D ;
  assign g2874 = \DFF_37.Q ;
  assign g28740 = \DFF_1564.D ;
  assign g28744 = \DFF_267.D ;
  assign g28745 = \DFF_272.D ;
  assign g28746 = \DFF_616.D ;
  assign g28747 = \DFF_621.D ;
  assign g28749 = \DFF_965.D ;
  assign g28754 = \DFF_273.D ;
  assign g28758 = \DFF_617.D ;
  assign g28759 = \DFF_622.D ;
  assign g28760 = \DFF_966.D ;
  assign g28761 = \DFF_971.D ;
  assign g28763 = \DFF_1315.D ;
  assign g28767 = \DFF_623.D ;
  assign g2877 = \DFF_46.Q ;
  assign g28771 = \DFF_967.D ;
  assign g28772 = \DFF_972.D ;
  assign g28773 = \DFF_1316.D ;
  assign g28774 = \DFF_1321.D ;
  assign g28778 = \DFF_973.D ;
  assign g2878 = \DFF_91.Q ;
  assign g28782 = \DFF_1317.D ;
  assign g28783 = \DFF_1322.D ;
  assign g28788 = \DFF_1323.D ;
  assign g2879 = \DFF_19.Q ;
  assign g288 = \DFF_312.Q ;
  assign g2883 = \DFF_4.Q ;
  assign g28832 = \DFF_141.D ;
  assign g28833 = \DFF_242.D ;
  assign g28835 = \DFF_592.D ;
  assign g28837 = \DFF_942.D ;
  assign g28839 = \DFF_1292.D ;
  assign g2888 = \DFF_5.Q ;
  assign g28882 = \DFF_468.D ;
  assign g28899 = \DFF_818.D ;
  assign g289 = \DFF_313.Q ;
  assign g28903 = \DFF_1017.D ;
  assign g2892 = \DFF_7.Q ;
  assign g28924 = \DFF_1168.D ;
  assign g28950 = \DFF_1518.D ;
  assign g2896 = \DFF_6.Q ;
  assign g28990 = \DFF_1142.D ;
  assign g290 = \DFF_314.Q ;
  assign g2900 = \DFF_9.Q ;
  assign g2903 = \DFF_8.Q ;
  assign g29061 = \DFF_426.D ;
  assign g29073 = \DFF_427.D ;
  assign g29074 = \DFF_423.D ;
  assign g29075 = \DFF_776.D ;
  assign g2908 = \DFF_10.Q ;
  assign g29081 = \DFF_428.D ;
  assign g29082 = \DFF_424.D ;
  assign g29084 = \DFF_777.D ;
  assign g29085 = \DFF_773.D ;
  assign g29086 = \DFF_1126.D ;
  assign g29089 = \DFF_425.D ;
  assign g29091 = \DFF_778.D ;
  assign g29092 = \DFF_774.D ;
  assign g29093 = \DFF_1127.D ;
  assign g29094 = \DFF_1123.D ;
  assign g29095 = \DFF_1476.D ;
  assign g29098 = \DFF_775.D ;
  assign g29099 = \DFF_1128.D ;
  assign g291 = \DFF_315.Q ;
  assign g29100 = \DFF_1124.D ;
  assign g29101 = \DFF_1477.D ;
  assign g29102 = \DFF_1473.D ;
  assign g29104 = \DFF_1125.D ;
  assign g29105 = \DFF_1478.D ;
  assign g29106 = \DFF_1474.D ;
  assign g29108 = \DFF_1475.D ;
  assign g29109 = \DFF_243.D ;
  assign g29110 = \DFF_593.D ;
  assign g29111 = \DFF_943.D ;
  assign g29112 = \DFF_1293.D ;
  assign g29113 = \DFF_1100.D ;
  assign g29117 = \DFF_110.D ;
  assign g29118 = \DFF_111.D ;
  assign g29119 = \DFF_112.D ;
  assign g2912 = \DFF_11.Q ;
  assign g29120 = \DFF_157.D ;
  assign g29131 = \DFF_242.D ;
  assign g29132 = \DFF_426.D ;
  assign g29133 = \DFF_427.D ;
  assign g29134 = \DFF_428.D ;
  assign g29135 = \DFF_423.D ;
  assign g29136 = \DFF_424.D ;
  assign g29137 = \DFF_425.D ;
  assign g29138 = \DFF_468.D ;
  assign g29139 = \DFF_592.D ;
  assign g29140 = \DFF_776.D ;
  assign g29141 = \DFF_777.D ;
  assign g29142 = \DFF_778.D ;
  assign g29143 = \DFF_773.D ;
  assign g29144 = \DFF_774.D ;
  assign g29145 = \DFF_775.D ;
  assign g29146 = \DFF_818.D ;
  assign g29147 = \DFF_942.D ;
  assign g29148 = \DFF_1126.D ;
  assign g29149 = \DFF_1127.D ;
  assign g29150 = \DFF_1128.D ;
  assign g29151 = \DFF_1123.D ;
  assign g29152 = \DFF_1124.D ;
  assign g29153 = \DFF_1125.D ;
  assign g29154 = \DFF_1168.D ;
  assign g29155 = \DFF_1292.D ;
  assign g29156 = \DFF_1476.D ;
  assign g29157 = \DFF_1477.D ;
  assign g29158 = \DFF_1478.D ;
  assign g29159 = \DFF_1473.D ;
  assign g29160 = \DFF_1474.D ;
  assign g29161 = \DFF_1475.D ;
  assign g29162 = \DFF_1518.D ;
  assign g29163 = \DFF_110.D ;
  assign g29164 = \DFF_111.D ;
  assign g29165 = \DFF_112.D ;
  assign g29166 = \DFF_141.D ;
  assign g29167 = \DFF_292.D ;
  assign g29169 = \DFF_293.D ;
  assign g2917 = \DFF_12.Q ;
  assign g29170 = \DFF_642.D ;
  assign g29172 = \DFF_294.D ;
  assign g29173 = \DFF_643.D ;
  assign g29178 = \DFF_992.D ;
  assign g29179 = \DFF_644.D ;
  assign g29181 = \DFF_993.D ;
  assign g29182 = \DFF_1342.D ;
  assign g29184 = \DFF_994.D ;
  assign g29185 = \DFF_1343.D ;
  assign g29187 = \DFF_1344.D ;
  assign g29192 = \DFF_1572.D ;
  assign g29194 = \DFF_268.D ;
  assign g29197 = \DFF_269.D ;
  assign g29198 = \DFF_618.D ;
  assign g2920 = \DFF_14.Q ;
  assign g29201 = \DFF_270.D ;
  assign g29204 = \DFF_619.D ;
  assign g29205 = \DFF_968.D ;
  assign g29209 = \DFF_620.D ;
  assign g29212 = \DFF_969.D ;
  assign g29213 = \DFF_1318.D ;
  assign g29218 = \DFF_970.D ;
  assign g29221 = \DFF_1319.D ;
  assign g29226 = \DFF_1320.D ;
  assign g29230 = \DFF_1100.D ;
  assign g29237 = \DFF_157.D ;
  assign g2924 = \DFF_13.Q ;
  assign g29244 = \DFF_157.D ;
  assign g29246 = \DFF_243.D ;
  assign g29249 = \DFF_593.D ;
  assign g29253 = \DFF_943.D ;
  assign g29258 = \DFF_1293.D ;
  assign g29267 = \DFF_1565.D ;
  assign g29270 = \DFF_1566.D ;
  assign g29273 = \DFF_1567.D ;
  assign g29276 = \DFF_1568.D ;
  assign g29278 = \DFF_1569.D ;
  assign g29279 = \DFF_1570.D ;
  assign g29281 = \DFF_1571.D ;
  assign g29288 = \DFF_1564.D ;
  assign g2929 = \DFF_18.Q ;
  assign g29293 = \DFF_265.D ;
  assign g29297 = \DFF_266.D ;
  assign g29298 = \DFF_271.D ;
  assign g29299 = \DFF_615.D ;
  assign g2930 = \DFF_17.Q ;
  assign g29304 = \DFF_267.D ;
  assign g29305 = \DFF_272.D ;
  assign g29306 = \DFF_616.D ;
  assign g29307 = \DFF_621.D ;
  assign g29308 = \DFF_965.D ;
  assign g29309 = \DFF_157.D ;
  assign g29311 = \DFF_273.D ;
  assign g29314 = \DFF_617.D ;
  assign g29315 = \DFF_622.D ;
  assign g29316 = \DFF_966.D ;
  assign g29317 = \DFF_971.D ;
  assign g29318 = \DFF_1142.D ;
  assign g29319 = \DFF_1315.D ;
  assign g29322 = \DFF_623.D ;
  assign g29325 = \DFF_967.D ;
  assign g29326 = \DFF_972.D ;
  assign g29327 = \DFF_1316.D ;
  assign g29328 = \DFF_1321.D ;
  assign g2933 = \DFF_2.Q ;
  assign g29331 = \DFF_973.D ;
  assign g29334 = \DFF_1317.D ;
  assign g29335 = \DFF_1322.D ;
  assign g29339 = \DFF_1323.D ;
  assign g2934 = \DFF_20.Q ;
  assign g2935 = \DFF_21.Q ;
  assign g29350 = \DFF_1100.D ;
  assign g29353 = \DFF_244.D ;
  assign g29354 = \DFF_594.D ;
  assign g29355 = \DFF_944.D ;
  assign g29356 = \DFF_160.D ;
  assign g29357 = \DFF_1294.D ;
  assign g29358 = \DFF_160.D ;
  assign g29359 = \DFF_1017.D ;
  assign g2938 = \DFF_22.Q ;
  assign g29401 = \DFF_1142.D ;
  assign g2941 = \DFF_23.Q ;
  assign g29412 = \DFF_1017.D ;
  assign g29413 = \DFF_243.D ;
  assign g29414 = \DFF_265.D ;
  assign g29415 = \DFF_266.D ;
  assign g29416 = \DFF_267.D ;
  assign g29417 = \DFF_271.D ;
  assign g29418 = \DFF_272.D ;
  assign g29419 = \DFF_273.D ;
  assign g29420 = \DFF_593.D ;
  assign g29421 = \DFF_615.D ;
  assign g29422 = \DFF_616.D ;
  assign g29423 = \DFF_617.D ;
  assign g29424 = \DFF_621.D ;
  assign g29425 = \DFF_622.D ;
  assign g29426 = \DFF_623.D ;
  assign g29427 = \DFF_943.D ;
  assign g29428 = \DFF_1017.D ;
  assign g29434 = \DFF_965.D ;
  assign g29435 = \DFF_966.D ;
  assign g29436 = \DFF_967.D ;
  assign g29437 = \DFF_971.D ;
  assign g29438 = \DFF_972.D ;
  assign g29439 = \DFF_973.D ;
  assign g2944 = \DFF_24.Q ;
  assign g29440 = \DFF_1142.D ;
  assign g29445 = \DFF_1100.D ;
  assign g29446 = \DFF_1293.D ;
  assign g29447 = \DFF_1315.D ;
  assign g29448 = \DFF_1316.D ;
  assign g29449 = \DFF_1317.D ;
  assign g29450 = \DFF_1321.D ;
  assign g29451 = \DFF_1322.D ;
  assign g29452 = \DFF_1323.D ;
  assign g29453 = \DFF_1564.D ;
  assign g29454 = \DFF_1565.D ;
  assign g29455 = \DFF_1566.D ;
  assign g29456 = \DFF_1567.D ;
  assign g29457 = \DFF_1568.D ;
  assign g29458 = \DFF_1569.D ;
  assign g29459 = \DFF_1570.D ;
  assign g29460 = \DFF_1571.D ;
  assign g29461 = \DFF_157.D ;
  assign g29462 = \DFF_157.D ;
  assign g29463 = \DFF_157.D ;
  assign g2947 = \DFF_25.Q ;
  assign g29495 = \DFF_160.D ;
  assign g29496 = \DFF_244.D ;
  assign g29497 = \DFF_160.D ;
  assign g29499 = \DFF_594.D ;
  assign g2950 = \DFF_3.Q ;
  assign g29501 = \DFF_944.D ;
  assign g29504 = \DFF_1294.D ;
  assign g29506 = \DFF_292.D ;
  assign g29507 = \DFF_293.D ;
  assign g29508 = \DFF_642.D ;
  assign g29509 = \DFF_294.D ;
  assign g29510 = \DFF_643.D ;
  assign g29511 = \DFF_992.D ;
  assign g29512 = \DFF_644.D ;
  assign g29513 = \DFF_993.D ;
  assign g29514 = \DFF_1342.D ;
  assign g29515 = \DFF_994.D ;
  assign g29516 = \DFF_1343.D ;
  assign g29517 = \DFF_1344.D ;
  assign g29519 = \DFF_1572.D ;
  assign g2953 = \DFF_26.Q ;
  assign g29530 = \DFF_268.D ;
  assign g29535 = \DFF_269.D ;
  assign g29537 = \DFF_618.D ;
  assign g29542 = \DFF_270.D ;
  assign g29544 = \DFF_619.D ;
  assign g29546 = \DFF_968.D ;
  assign g29551 = \DFF_620.D ;
  assign g29554 = \DFF_969.D ;
  assign g29556 = \DFF_1318.D ;
  assign g2956 = \DFF_27.Q ;
  assign g29561 = \DFF_970.D ;
  assign g29563 = \DFF_1319.D ;
  assign g29568 = \DFF_1320.D ;
  assign g29579 = \DFF_245.D ;
  assign g29580 = \DFF_595.D ;
  assign g29581 = \DFF_945.D ;
  assign g29582 = \DFF_1295.D ;
  assign g2959 = \DFF_28.Q ;
  assign g29606 = \DFF_283.D ;
  assign g29608 = \DFF_284.D ;
  assign g29609 = \DFF_633.D ;
  assign g29611 = \DFF_285.D ;
  assign g29612 = \DFF_634.D ;
  assign g29613 = \DFF_983.D ;
  assign g29616 = \DFF_635.D ;
  assign g29617 = \DFF_984.D ;
  assign g29618 = \DFF_1333.D ;
  assign g2962 = \DFF_29.Q ;
  assign g29620 = \DFF_985.D ;
  assign g29621 = \DFF_1334.D ;
  assign g29623 = \DFF_1335.D ;
  assign g29627 = \DFF_244.D ;
  assign g29628 = \DFF_292.D ;
  assign g29629 = \DFF_293.D ;
  assign g2963 = \DFF_30.Q ;
  assign g29630 = \DFF_294.D ;
  assign g29631 = \DFF_268.D ;
  assign g29632 = \DFF_269.D ;
  assign g29633 = \DFF_270.D ;
  assign g29634 = \DFF_594.D ;
  assign g29635 = \DFF_642.D ;
  assign g29636 = \DFF_643.D ;
  assign g29637 = \DFF_644.D ;
  assign g29638 = \DFF_618.D ;
  assign g29639 = \DFF_619.D ;
  assign g29640 = \DFF_620.D ;
  assign g29641 = \DFF_944.D ;
  assign g29642 = \DFF_992.D ;
  assign g29643 = \DFF_993.D ;
  assign g29644 = \DFF_994.D ;
  assign g29645 = \DFF_968.D ;
  assign g29646 = \DFF_969.D ;
  assign g29647 = \DFF_970.D ;
  assign g29648 = \DFF_1294.D ;
  assign g29649 = \DFF_1342.D ;
  assign g29650 = \DFF_1343.D ;
  assign g29651 = \DFF_1344.D ;
  assign g29652 = \DFF_1318.D ;
  assign g29653 = \DFF_1319.D ;
  assign g29654 = \DFF_1320.D ;
  assign g29655 = \DFF_1572.D ;
  assign g29656 = \DFF_160.D ;
  assign g29657 = \DFF_160.D ;
  assign g29658 = \DFF_1580.D ;
  assign g29659 = \DFF_1579.D ;
  assign g2966 = \DFF_31.Q ;
  assign g29660 = \DFF_1578.D ;
  assign g29661 = \DFF_1577.D ;
  assign g29662 = \DFF_1576.D ;
  assign g29664 = \DFF_1575.D ;
  assign g29666 = \DFF_1574.D ;
  assign g29668 = \DFF_1573.D ;
  assign g29689 = \DFF_245.D ;
  assign g2969 = \DFF_32.Q ;
  assign g29690 = \DFF_283.D ;
  assign g29691 = \DFF_284.D ;
  assign g29692 = \DFF_595.D ;
  assign g29693 = \DFF_633.D ;
  assign g29694 = \DFF_285.D ;
  assign g29695 = \DFF_634.D ;
  assign g29696 = \DFF_945.D ;
  assign g29697 = \DFF_983.D ;
  assign g29698 = \DFF_635.D ;
  assign g29699 = \DFF_984.D ;
  assign g29700 = \DFF_1295.D ;
  assign g29701 = \DFF_1333.D ;
  assign g29702 = \DFF_985.D ;
  assign g29704 = \DFF_1334.D ;
  assign g29708 = \DFF_1335.D ;
  assign g2972 = \DFF_33.Q ;
  assign g2975 = \DFF_34.Q ;
  assign g2978 = \DFF_35.Q ;
  assign g29794 = \DFF_245.D ;
  assign g29795 = \DFF_283.D ;
  assign g29796 = \DFF_284.D ;
  assign g29797 = \DFF_285.D ;
  assign g29798 = \DFF_595.D ;
  assign g29799 = \DFF_633.D ;
  assign g298 = \DFF_328.Q ;
  assign g29800 = \DFF_634.D ;
  assign g29801 = \DFF_635.D ;
  assign g29802 = \DFF_945.D ;
  assign g29803 = \DFF_983.D ;
  assign g29804 = \DFF_984.D ;
  assign g29805 = \DFF_985.D ;
  assign g29806 = \DFF_1295.D ;
  assign g29807 = \DFF_1333.D ;
  assign g29808 = \DFF_1334.D ;
  assign g29809 = \DFF_1335.D ;
  assign g2981 = \DFF_36.Q ;
  assign g2984 = \DFF_15.Q ;
  assign g29848 = \DFF_1581.D ;
  assign g2985 = \DFF_16.Q ;
  assign g2986 = \DFF_1612.Q ;
  assign g2987 = \DFF_1613.Q ;
  assign g299 = \DFF_316.Q ;
  assign g2990 = \DFF_1633.Q ;
  assign g2991 = \DFF_1634.Q ;
  assign g2992 = \DFF_1624.Q ;
  assign g2993 = \DFF_1600.Q ;
  assign g29932 = \DFF_1575.D ;
  assign g29933 = \DFF_1576.D ;
  assign g29934 = \DFF_1577.D ;
  assign g29935 = \DFF_1578.D ;
  assign g29936 = \DFF_113.D ;
  assign g29937 = \DFF_1579.D ;
  assign g29938 = \DFF_1580.D ;
  assign g29939 = \DFF_114.D ;
  assign g29940 = \DFF_1573.D ;
  assign g29941 = \DFF_115.D ;
  assign g29943 = \DFF_1574.D ;
  assign g2997 = \DFF_1599.Q ;
  assign g29972 = \DFF_1573.D ;
  assign g29973 = \DFF_1574.D ;
  assign g29974 = \DFF_1575.D ;
  assign g29975 = \DFF_1576.D ;
  assign g29976 = \DFF_1577.D ;
  assign g29977 = \DFF_1578.D ;
  assign g29978 = \DFF_1579.D ;
  assign g29979 = \DFF_1580.D ;
  assign g2998 = \DFF_1601.Q ;
  assign g30 = \DFF_1619.Q ;
  assign g3002 = \DFF_1603.Q ;
  assign g30052 = \DFF_1581.D ;
  assign g30055 = \DFF_1367.D ;
  assign g3006 = \DFF_1602.Q ;
  assign g30061 = \DFF_1492.D ;
  assign g30072 = \DFF_1450.D ;
  assign g30076 = \DFF_113.D ;
  assign g30078 = \DFF_114.D ;
  assign g30084 = \DFF_115.D ;
  assign g3010 = \DFF_1605.Q ;
  assign g30119 = \DFF_1581.D ;
  assign g30120 = \DFF_113.D ;
  assign g30121 = \DFF_114.D ;
  assign g30122 = \DFF_115.D ;
  assign g30124 = \DFF_1367.D ;
  assign g3013 = \DFF_1604.Q ;
  assign g3018 = \DFF_1607.Q ;
  assign g30215 = \DFF_1450.D ;
  assign g3024 = \DFF_1606.Q ;
  assign g30245 = \DFF_224.D ;
  assign g30246 = \DFF_225.D ;
  assign g30247 = \DFF_574.D ;
  assign g30248 = \DFF_226.D ;
  assign g30249 = \DFF_575.D ;
  assign g30250 = \DFF_924.D ;
  assign g30251 = \DFF_576.D ;
  assign g30252 = \DFF_925.D ;
  assign g30253 = \DFF_1274.D ;
  assign g30254 = \DFF_221.D ;
  assign g30255 = \DFF_926.D ;
  assign g30256 = \DFF_1275.D ;
  assign g30257 = \DFF_222.D ;
  assign g30258 = \DFF_227.D ;
  assign g30259 = \DFF_571.D ;
  assign g30260 = \DFF_1276.D ;
  assign g30261 = \DFF_206.D ;
  assign g30262 = \DFF_223.D ;
  assign g30263 = \DFF_228.D ;
  assign g30264 = \DFF_572.D ;
  assign g30265 = \DFF_577.D ;
  assign g30266 = \DFF_921.D ;
  assign g30267 = \DFF_207.D ;
  assign g30268 = \DFF_229.D ;
  assign g30269 = \DFF_556.D ;
  assign g30270 = \DFF_573.D ;
  assign g30271 = \DFF_578.D ;
  assign g30272 = \DFF_922.D ;
  assign g30273 = \DFF_927.D ;
  assign g30274 = \DFF_1271.D ;
  assign g30275 = \DFF_208.D ;
  assign g30276 = \DFF_218.D ;
  assign g30277 = \DFF_557.D ;
  assign g30278 = \DFF_579.D ;
  assign g30279 = \DFF_906.D ;
  assign g3028 = \DFF_1608.Q ;
  assign g30280 = \DFF_923.D ;
  assign g30281 = \DFF_928.D ;
  assign g30282 = \DFF_1272.D ;
  assign g30283 = \DFF_1277.D ;
  assign g30284 = \DFF_219.D ;
  assign g30285 = \DFF_558.D ;
  assign g30286 = \DFF_568.D ;
  assign g30287 = \DFF_907.D ;
  assign g30288 = \DFF_929.D ;
  assign g30289 = \DFF_1256.D ;
  assign g30290 = \DFF_1273.D ;
  assign g30291 = \DFF_1278.D ;
  assign g30292 = \DFF_220.D ;
  assign g30293 = \DFF_569.D ;
  assign g30294 = \DFF_908.D ;
  assign g30295 = \DFF_918.D ;
  assign g30296 = \DFF_1257.D ;
  assign g30297 = \DFF_1279.D ;
  assign g30298 = \DFF_570.D ;
  assign g30299 = \DFF_919.D ;
  assign g30300 = \DFF_1258.D ;
  assign g30301 = \DFF_1268.D ;
  assign g30302 = \DFF_920.D ;
  assign g30303 = \DFF_1269.D ;
  assign g30304 = \DFF_1270.D ;
  assign g30306 = \DFF_1450.D ;
  assign g30308 = \DFF_1492.D ;
  assign g30314 = \DFF_1367.D ;
  assign g3032 = \DFF_1610.Q ;
  assign g30320 = \DFF_1492.D ;
  assign g30325 = \DFF_1450.D ;
  assign g30326 = \DFF_207.D ;
  assign g30328 = \DFF_229.D ;
  assign g30329 = \DFF_556.D ;
  assign g30331 = \DFF_573.D ;
  assign g30332 = \DFF_578.D ;
  assign g30335 = \DFF_922.D ;
  assign g30336 = \DFF_927.D ;
  assign g30338 = \DFF_991.D ;
  assign g30339 = \DFF_1271.D ;
  assign g30341 = \DFF_1340.D ;
  assign g30342 = \DFF_208.D ;
  assign g30343 = \DFF_218.D ;
  assign g30344 = \DFF_557.D ;
  assign g30346 = \DFF_579.D ;
  assign g30347 = \DFF_906.D ;
  assign g30349 = \DFF_923.D ;
  assign g30350 = \DFF_928.D ;
  assign g30353 = \DFF_1272.D ;
  assign g30354 = \DFF_1277.D ;
  assign g30356 = \DFF_1341.D ;
  assign g30357 = \DFF_219.D ;
  assign g30358 = \DFF_558.D ;
  assign g30359 = \DFF_568.D ;
  assign g3036 = \DFF_1609.Q ;
  assign g30360 = \DFF_907.D ;
  assign g30362 = \DFF_929.D ;
  assign g30363 = \DFF_1256.D ;
  assign g30365 = \DFF_1273.D ;
  assign g30366 = \DFF_1278.D ;
  assign g30368 = \DFF_220.D ;
  assign g30369 = \DFF_569.D ;
  assign g30370 = \DFF_908.D ;
  assign g30371 = \DFF_918.D ;
  assign g30373 = \DFF_1257.D ;
  assign g30375 = \DFF_1279.D ;
  assign g30376 = \DFF_570.D ;
  assign g30377 = \DFF_919.D ;
  assign g30378 = \DFF_1258.D ;
  assign g30379 = \DFF_1268.D ;
  assign g30380 = \DFF_920.D ;
  assign g30381 = \DFF_1269.D ;
  assign g30382 = \DFF_1270.D ;
  assign g3040 = \DFF_1611.Q ;
  assign g30408 = \DFF_224.D ;
  assign g3043 = \DFF_1564.Q ;
  assign g30435 = \DFF_225.D ;
  assign g30439 = \DFF_574.D ;
  assign g3044 = \DFF_1565.Q ;
  assign g30443 = \DFF_226.D ;
  assign g30446 = \DFF_575.D ;
  assign g3045 = \DFF_1566.Q ;
  assign g30450 = \DFF_924.D ;
  assign g30455 = \DFF_289.D ;
  assign g30456 = \DFF_576.D ;
  assign g30459 = \DFF_925.D ;
  assign g3046 = \DFF_1567.Q ;
  assign g30463 = \DFF_1274.D ;
  assign g30466 = \DFF_221.D ;
  assign g30468 = \DFF_290.D ;
  assign g3047 = \DFF_1568.Q ;
  assign g30470 = \DFF_639.D ;
  assign g30471 = \DFF_926.D ;
  assign g30474 = \DFF_1275.D ;
  assign g30479 = \DFF_222.D ;
  assign g3048 = \DFF_1569.Q ;
  assign g30480 = \DFF_227.D ;
  assign g30482 = \DFF_291.D ;
  assign g30483 = \DFF_571.D ;
  assign g30485 = \DFF_640.D ;
  assign g30487 = \DFF_989.D ;
  assign g30488 = \DFF_1276.D ;
  assign g3049 = \DFF_1570.Q ;
  assign g30491 = \DFF_206.D ;
  assign g30493 = \DFF_223.D ;
  assign g30494 = \DFF_228.D ;
  assign g30497 = \DFF_572.D ;
  assign g30498 = \DFF_577.D ;
  assign g305 = \DFF_317.Q ;
  assign g3050 = \DFF_1571.Q ;
  assign g30500 = \DFF_641.D ;
  assign g30501 = \DFF_921.D ;
  assign g30503 = \DFF_990.D ;
  assign g30505 = \DFF_1339.D ;
  assign g30506 = \DFF_206.D ;
  assign g30507 = \DFF_207.D ;
  assign g30508 = \DFF_208.D ;
  assign g30509 = \DFF_218.D ;
  assign g3051 = \DFF_1572.Q ;
  assign g30510 = \DFF_219.D ;
  assign g30511 = \DFF_220.D ;
  assign g30512 = \DFF_224.D ;
  assign g30513 = \DFF_225.D ;
  assign g30514 = \DFF_226.D ;
  assign g30515 = \DFF_221.D ;
  assign g30516 = \DFF_222.D ;
  assign g30517 = \DFF_223.D ;
  assign g30518 = \DFF_227.D ;
  assign g30519 = \DFF_228.D ;
  assign g3052 = \DFF_1573.Q ;
  assign g30520 = \DFF_229.D ;
  assign g30521 = \DFF_556.D ;
  assign g30522 = \DFF_557.D ;
  assign g30523 = \DFF_558.D ;
  assign g30524 = \DFF_568.D ;
  assign g30525 = \DFF_569.D ;
  assign g30526 = \DFF_570.D ;
  assign g30527 = \DFF_574.D ;
  assign g30528 = \DFF_575.D ;
  assign g30529 = \DFF_576.D ;
  assign g3053 = \DFF_1574.Q ;
  assign g30530 = \DFF_571.D ;
  assign g30531 = \DFF_572.D ;
  assign g30532 = \DFF_573.D ;
  assign g30533 = \DFF_577.D ;
  assign g30534 = \DFF_578.D ;
  assign g30535 = \DFF_579.D ;
  assign g30536 = \DFF_906.D ;
  assign g30537 = \DFF_907.D ;
  assign g30538 = \DFF_908.D ;
  assign g30539 = \DFF_918.D ;
  assign g3054 = \DFF_1561.Q ;
  assign g30540 = \DFF_919.D ;
  assign g30541 = \DFF_920.D ;
  assign g30542 = \DFF_924.D ;
  assign g30543 = \DFF_925.D ;
  assign g30544 = \DFF_926.D ;
  assign g30545 = \DFF_921.D ;
  assign g30546 = \DFF_922.D ;
  assign g30547 = \DFF_923.D ;
  assign g30548 = \DFF_927.D ;
  assign g30549 = \DFF_928.D ;
  assign g3055 = \DFF_1575.Q ;
  assign g30550 = \DFF_929.D ;
  assign g30551 = \DFF_1256.D ;
  assign g30552 = \DFF_1257.D ;
  assign g30553 = \DFF_1258.D ;
  assign g30554 = \DFF_1268.D ;
  assign g30555 = \DFF_1269.D ;
  assign g30556 = \DFF_1270.D ;
  assign g30557 = \DFF_1274.D ;
  assign g30558 = \DFF_1275.D ;
  assign g30559 = \DFF_1276.D ;
  assign g3056 = \DFF_1576.Q ;
  assign g30560 = \DFF_1271.D ;
  assign g30561 = \DFF_1272.D ;
  assign g30562 = \DFF_1273.D ;
  assign g30563 = \DFF_1277.D ;
  assign g30564 = \DFF_1278.D ;
  assign g30565 = \DFF_1279.D ;
  assign g30566 = \DFF_1338.D ;
  assign g30567 = \DFF_1589.D ;
  assign g30568 = \DFF_1588.D ;
  assign g30569 = \DFF_1587.D ;
  assign g3057 = \DFF_1577.Q ;
  assign g30570 = \DFF_1586.D ;
  assign g30571 = \DFF_1585.D ;
  assign g30572 = \DFF_1584.D ;
  assign g30573 = \DFF_1583.D ;
  assign g30574 = \DFF_1582.D ;
  assign g30578 = \DFF_289.D ;
  assign g30579 = \DFF_290.D ;
  assign g3058 = \DFF_1578.Q ;
  assign g30580 = \DFF_639.D ;
  assign g30581 = \DFF_291.D ;
  assign g30582 = \DFF_640.D ;
  assign g30583 = \DFF_989.D ;
  assign g30585 = \DFF_641.D ;
  assign g30586 = \DFF_990.D ;
  assign g30587 = \DFF_1339.D ;
  assign g3059 = \DFF_1579.Q ;
  assign g30591 = \DFF_991.D ;
  assign g30592 = \DFF_1340.D ;
  assign g3060 = \DFF_1580.Q ;
  assign g30600 = \DFF_1341.D ;
  assign g3061 = \DFF_1581.Q ;
  assign g3062 = \DFF_1582.Q ;
  assign g3063 = \DFF_1583.Q ;
  assign g30635 = \DFF_230.D ;
  assign g30636 = \DFF_231.D ;
  assign g30637 = \DFF_209.D ;
  assign g30638 = \DFF_580.D ;
  assign g30639 = \DFF_232.D ;
  assign g3064 = \DFF_1584.Q ;
  assign g30640 = \DFF_210.D ;
  assign g30641 = \DFF_215.D ;
  assign g30642 = \DFF_581.D ;
  assign g30643 = \DFF_559.D ;
  assign g30644 = \DFF_930.D ;
  assign g30645 = \DFF_211.D ;
  assign g30646 = \DFF_216.D ;
  assign g30647 = \DFF_582.D ;
  assign g30648 = \DFF_560.D ;
  assign g30649 = \DFF_565.D ;
  assign g3065 = \DFF_1585.Q ;
  assign g30650 = \DFF_931.D ;
  assign g30651 = \DFF_909.D ;
  assign g30652 = \DFF_1280.D ;
  assign g30653 = \DFF_217.D ;
  assign g30654 = \DFF_561.D ;
  assign g30655 = \DFF_566.D ;
  assign g30656 = \DFF_932.D ;
  assign g30657 = \DFF_910.D ;
  assign g30658 = \DFF_915.D ;
  assign g30659 = \DFF_1281.D ;
  assign g3066 = \DFF_1586.Q ;
  assign g30660 = \DFF_1259.D ;
  assign g30661 = \DFF_233.D ;
  assign g30662 = \DFF_567.D ;
  assign g30663 = \DFF_911.D ;
  assign g30664 = \DFF_916.D ;
  assign g30665 = \DFF_1282.D ;
  assign g30666 = \DFF_1260.D ;
  assign g30667 = \DFF_1265.D ;
  assign g30668 = \DFF_212.D ;
  assign g30669 = \DFF_234.D ;
  assign g3067 = \DFF_1587.Q ;
  assign g30670 = \DFF_583.D ;
  assign g30671 = \DFF_917.D ;
  assign g30672 = \DFF_1261.D ;
  assign g30673 = \DFF_1266.D ;
  assign g30674 = \DFF_213.D ;
  assign g30675 = \DFF_235.D ;
  assign g30676 = \DFF_562.D ;
  assign g30677 = \DFF_584.D ;
  assign g30678 = \DFF_933.D ;
  assign g30679 = \DFF_1267.D ;
  assign g3068 = \DFF_1588.Q ;
  assign g30680 = \DFF_214.D ;
  assign g30681 = \DFF_563.D ;
  assign g30682 = \DFF_585.D ;
  assign g30683 = \DFF_912.D ;
  assign g30684 = \DFF_934.D ;
  assign g30686 = \DFF_1283.D ;
  assign g30687 = \DFF_564.D ;
  assign g30688 = \DFF_913.D ;
  assign g30689 = \DFF_935.D ;
  assign g3069 = \DFF_1589.Q ;
  assign g30690 = \DFF_1262.D ;
  assign g30691 = \DFF_1284.D ;
  assign g30692 = \DFF_914.D ;
  assign g30693 = \DFF_1263.D ;
  assign g30694 = \DFF_1285.D ;
  assign g30695 = \DFF_1264.D ;
  assign g30699 = \DFF_286.D ;
  assign g3070 = \DFF_1590.Q ;
  assign g30700 = \DFF_287.D ;
  assign g30701 = \DFF_636.D ;
  assign g30702 = \DFF_288.D ;
  assign g30703 = \DFF_637.D ;
  assign g30704 = \DFF_986.D ;
  assign g30705 = \DFF_638.D ;
  assign g30706 = \DFF_987.D ;
  assign g30707 = \DFF_1336.D ;
  assign g30708 = \DFF_988.D ;
  assign g30709 = \DFF_1337.D ;
  assign g3071 = \DFF_1591.Q ;
  assign g30710 = \DFF_289.D ;
  assign g30711 = \DFF_290.D ;
  assign g30712 = \DFF_291.D ;
  assign g30713 = \DFF_639.D ;
  assign g30714 = \DFF_640.D ;
  assign g30715 = \DFF_641.D ;
  assign g30716 = \DFF_989.D ;
  assign g30717 = \DFF_990.D ;
  assign g30718 = \DFF_991.D ;
  assign g30719 = \DFF_1339.D ;
  assign g3072 = \DFF_1592.Q ;
  assign g30720 = \DFF_1340.D ;
  assign g30721 = \DFF_1341.D ;
  assign g30722 = \DFF_212.D ;
  assign g30723 = \DFF_234.D ;
  assign g30724 = \DFF_583.D ;
  assign g30725 = \DFF_917.D ;
  assign g30726 = \DFF_1261.D ;
  assign g30727 = \DFF_1266.D ;
  assign g30729 = \DFF_213.D ;
  assign g3073 = \DFF_1593.Q ;
  assign g30730 = \DFF_235.D ;
  assign g30731 = \DFF_562.D ;
  assign g30732 = \DFF_584.D ;
  assign g30733 = \DFF_933.D ;
  assign g30734 = \DFF_1267.D ;
  assign g30737 = \DFF_214.D ;
  assign g30738 = \DFF_563.D ;
  assign g30739 = \DFF_585.D ;
  assign g3074 = \DFF_1594.Q ;
  assign g30740 = \DFF_912.D ;
  assign g30741 = \DFF_934.D ;
  assign g30742 = \DFF_1283.D ;
  assign g30745 = \DFF_564.D ;
  assign g30746 = \DFF_913.D ;
  assign g30747 = \DFF_935.D ;
  assign g30748 = \DFF_1262.D ;
  assign g30749 = \DFF_1284.D ;
  assign g3075 = \DFF_1595.Q ;
  assign g30751 = \DFF_914.D ;
  assign g30752 = \DFF_1263.D ;
  assign g30753 = \DFF_1285.D ;
  assign g30756 = \DFF_1264.D ;
  assign g3076 = \DFF_1596.Q ;
  assign g30765 = \DFF_1590.D ;
  assign g30767 = \DFF_286.D ;
  assign g30769 = \DFF_287.D ;
  assign g3077 = \DFF_1597.Q ;
  assign g30770 = \DFF_636.D ;
  assign g30772 = \DFF_288.D ;
  assign g30773 = \DFF_637.D ;
  assign g30774 = \DFF_986.D ;
  assign g30776 = \DFF_638.D ;
  assign g30777 = \DFF_987.D ;
  assign g30778 = \DFF_1336.D ;
  assign g3078 = \DFF_1598.Q ;
  assign g30781 = \DFF_988.D ;
  assign g30782 = \DFF_1337.D ;
  assign g30784 = \DFF_1338.D ;
  assign g3079 = \DFF_1562.Q ;
  assign g30792 = \DFF_1585.D ;
  assign g30793 = \DFF_1586.D ;
  assign g30794 = \DFF_1587.D ;
  assign g30795 = \DFF_1588.D ;
  assign g30796 = \DFF_116.D ;
  assign g30797 = \DFF_1589.D ;
  assign g30798 = \DFF_117.D ;
  assign g30799 = \DFF_1582.D ;
  assign g3080 = \DFF_1563.Q ;
  assign g30800 = \DFF_1583.D ;
  assign g30801 = \DFF_118.D ;
  assign g30802 = \DFF_1584.D ;
  assign g30803 = \DFF_230.D ;
  assign g30804 = \DFF_231.D ;
  assign g30805 = \DFF_209.D ;
  assign g30806 = \DFF_580.D ;
  assign g30807 = \DFF_232.D ;
  assign g30808 = \DFF_210.D ;
  assign g30809 = \DFF_215.D ;
  assign g30810 = \DFF_581.D ;
  assign g30811 = \DFF_559.D ;
  assign g30812 = \DFF_930.D ;
  assign g30813 = \DFF_211.D ;
  assign g30814 = \DFF_216.D ;
  assign g30815 = \DFF_582.D ;
  assign g30816 = \DFF_560.D ;
  assign g30817 = \DFF_565.D ;
  assign g30818 = \DFF_931.D ;
  assign g30819 = \DFF_909.D ;
  assign g30820 = \DFF_1280.D ;
  assign g30821 = \DFF_217.D ;
  assign g30822 = \DFF_561.D ;
  assign g30823 = \DFF_566.D ;
  assign g30824 = \DFF_932.D ;
  assign g30825 = \DFF_910.D ;
  assign g30826 = \DFF_915.D ;
  assign g30827 = \DFF_1281.D ;
  assign g30828 = \DFF_1259.D ;
  assign g30829 = \DFF_233.D ;
  assign g3083 = \DFF_1622.Q ;
  assign g30830 = \DFF_567.D ;
  assign g30831 = \DFF_911.D ;
  assign g30832 = \DFF_916.D ;
  assign g30833 = \DFF_1282.D ;
  assign g30834 = \DFF_1260.D ;
  assign g30835 = \DFF_1265.D ;
  assign g30836 = \DFF_212.D ;
  assign g30837 = \DFF_213.D ;
  assign g30838 = \DFF_214.D ;
  assign g30839 = \DFF_230.D ;
  assign g3084 = \DFF_97.Q ;
  assign g30840 = \DFF_231.D ;
  assign g30841 = \DFF_232.D ;
  assign g30842 = \DFF_209.D ;
  assign g30843 = \DFF_210.D ;
  assign g30844 = \DFF_211.D ;
  assign g30845 = \DFF_215.D ;
  assign g30846 = \DFF_216.D ;
  assign g30847 = \DFF_217.D ;
  assign g30848 = \DFF_233.D ;
  assign g30849 = \DFF_234.D ;
  assign g3085 = \DFF_98.Q ;
  assign g30850 = \DFF_235.D ;
  assign g30851 = \DFF_286.D ;
  assign g30852 = \DFF_287.D ;
  assign g30853 = \DFF_288.D ;
  assign g30854 = \DFF_562.D ;
  assign g30855 = \DFF_563.D ;
  assign g30856 = \DFF_564.D ;
  assign g30857 = \DFF_580.D ;
  assign g30858 = \DFF_581.D ;
  assign g30859 = \DFF_582.D ;
  assign g3086 = \DFF_99.Q ;
  assign g30860 = \DFF_559.D ;
  assign g30861 = \DFF_560.D ;
  assign g30862 = \DFF_561.D ;
  assign g30863 = \DFF_565.D ;
  assign g30864 = \DFF_566.D ;
  assign g30865 = \DFF_567.D ;
  assign g30866 = \DFF_583.D ;
  assign g30867 = \DFF_584.D ;
  assign g30868 = \DFF_585.D ;
  assign g30869 = \DFF_636.D ;
  assign g3087 = \DFF_100.Q ;
  assign g30870 = \DFF_637.D ;
  assign g30871 = \DFF_638.D ;
  assign g30872 = \DFF_912.D ;
  assign g30873 = \DFF_913.D ;
  assign g30874 = \DFF_914.D ;
  assign g30875 = \DFF_930.D ;
  assign g30876 = \DFF_931.D ;
  assign g30877 = \DFF_932.D ;
  assign g30878 = \DFF_909.D ;
  assign g30879 = \DFF_910.D ;
  assign g3088 = \DFF_130.Q ;
  assign g30880 = \DFF_911.D ;
  assign g30881 = \DFF_915.D ;
  assign g30882 = \DFF_916.D ;
  assign g30883 = \DFF_917.D ;
  assign g30884 = \DFF_933.D ;
  assign g30885 = \DFF_934.D ;
  assign g30886 = \DFF_935.D ;
  assign g30887 = \DFF_986.D ;
  assign g30888 = \DFF_987.D ;
  assign g30889 = \DFF_988.D ;
  assign g30890 = \DFF_1262.D ;
  assign g30891 = \DFF_1263.D ;
  assign g30892 = \DFF_1264.D ;
  assign g30893 = \DFF_1280.D ;
  assign g30894 = \DFF_1281.D ;
  assign g30895 = \DFF_1282.D ;
  assign g30896 = \DFF_1259.D ;
  assign g30897 = \DFF_1260.D ;
  assign g30898 = \DFF_1261.D ;
  assign g30899 = \DFF_1265.D ;
  assign g309 = \DFF_1302.Q ;
  assign g30900 = \DFF_1266.D ;
  assign g30901 = \DFF_1267.D ;
  assign g30902 = \DFF_1283.D ;
  assign g30903 = \DFF_1284.D ;
  assign g30904 = \DFF_1285.D ;
  assign g30905 = \DFF_1336.D ;
  assign g30906 = \DFF_1337.D ;
  assign g30907 = \DFF_1338.D ;
  assign g30908 = \DFF_1582.D ;
  assign g30909 = \DFF_1583.D ;
  assign g3091 = \DFF_101.Q ;
  assign g30910 = \DFF_1584.D ;
  assign g30911 = \DFF_1585.D ;
  assign g30912 = \DFF_1586.D ;
  assign g30913 = \DFF_1587.D ;
  assign g30914 = \DFF_1588.D ;
  assign g30915 = \DFF_1589.D ;
  assign g3092 = \DFF_102.Q ;
  assign g30928 = \DFF_1590.D ;
  assign g3093 = \DFF_103.Q ;
  assign g30937 = \DFF_116.D ;
  assign g30938 = \DFF_117.D ;
  assign g30939 = \DFF_118.D ;
  assign g3094 = \DFF_104.Q ;
  assign g30940 = \DFF_1590.D ;
  assign g30941 = \DFF_116.D ;
  assign g30942 = \DFF_117.D ;
  assign g30943 = \DFF_118.D ;
  assign g3095 = \DFF_105.Q ;
  assign g3096 = \DFF_106.Q ;
  assign g30962 = \DFF_1598.D ;
  assign g30963 = \DFF_1597.D ;
  assign g30964 = \DFF_1596.D ;
  assign g30965 = \DFF_1595.D ;
  assign g30966 = \DFF_1594.D ;
  assign g30967 = \DFF_1593.D ;
  assign g30968 = \DFF_1592.D ;
  assign g30969 = \DFF_1591.D ;
  assign g3097 = \DFF_107.Q ;
  assign g30971 = \DFF_1599.D ;
  assign g30972 = \DFF_1595.D ;
  assign g30973 = \DFF_1596.D ;
  assign g30974 = \DFF_1597.D ;
  assign g30975 = \DFF_1598.D ;
  assign g30976 = \DFF_1591.D ;
  assign g30977 = \DFF_1592.D ;
  assign g30978 = \DFF_1593.D ;
  assign g30979 = \DFF_1594.D ;
  assign g3098 = \DFF_108.Q ;
  assign g30980 = \DFF_1591.D ;
  assign g30981 = \DFF_1592.D ;
  assign g30982 = \DFF_1593.D ;
  assign g30983 = \DFF_1594.D ;
  assign g30984 = \DFF_1595.D ;
  assign g30985 = \DFF_1596.D ;
  assign g30986 = \DFF_1597.D ;
  assign g30987 = \DFF_1598.D ;
  assign g30988 = \DFF_1599.D ;
  assign g30989 = \DFF_1599.D ;
  assign g3099 = \DFF_109.Q ;
  assign g3100 = \DFF_110.Q ;
  assign g3101 = \DFF_111.Q ;
  assign g3102 = \DFF_112.Q ;
  assign g3103 = \DFF_113.Q ;
  assign g3104 = \DFF_114.Q ;
  assign g3105 = \DFF_115.Q ;
  assign g3106 = \DFF_116.Q ;
  assign g3107 = \DFF_117.Q ;
  assign g3108 = \DFF_118.Q ;
  assign g3109 = \DFF_1506.Q ;
  assign g3110 = \DFF_151.Q ;
  assign g3111 = \DFF_152.Q ;
  assign g3112 = \DFF_150.Q ;
  assign g3113 = \DFF_156.Q ;
  assign g3114 = \DFF_159.Q ;
  assign g3117 = \DFF_1505.Q ;
  assign g312 = \DFF_283.Q ;
  assign g3120 = \DFF_158.Q ;
  assign g3123 = \DFF_146.Q ;
  assign g3124 = \DFF_152.Q ;
  assign g3125 = \DFF_144.Q ;
  assign g3126 = \DFF_150.Q ;
  assign g3127 = \DFF_156.Q ;
  assign g3128 = \DFF_141.Q ;
  assign g3129 = \DFF_1504.Q ;
  assign g313 = \DFF_284.Q ;
  assign g3132 = \DFF_158.Q ;
  assign g3133 = \DFF_160.Q ;
  assign g3134 = \DFF_159.Q ;
  assign g3135 = \DFF_156.Q ;
  assign g3136 = \DFF_158.Q ;
  assign g3139 = \DFF_157.Q ;
  assign g314 = \DFF_285.Q ;
  assign g3142 = \DFF_158.Q ;
  assign g3147 = \DFF_159.Q ;
  assign g315 = \DFF_286.Q ;
  assign g3151 = \DFF_157.Q ;
  assign g3155 = \DFF_119.Q ;
  assign g3158 = \DFF_120.Q ;
  assign g316 = \DFF_287.Q ;
  assign g3161 = \DFF_121.Q ;
  assign g3164 = \DFF_122.Q ;
  assign g3167 = \DFF_123.Q ;
  assign g317 = \DFF_288.Q ;
  assign g3170 = \DFF_124.Q ;
  assign g3173 = \DFF_125.Q ;
  assign g3176 = \DFF_126.Q ;
  assign g3179 = \DFF_127.Q ;
  assign g318 = \DFF_289.Q ;
  assign g3182 = \DFF_128.Q ;
  assign g3185 = \DFF_129.Q ;
  assign g3188 = \DFF_157.Q ;
  assign g319 = \DFF_290.Q ;
  assign g3191 = \DFF_131.Q ;
  assign g3194 = \DFF_152.Q ;
  assign g3197 = \DFF_151.Q ;
  assign g3198 = \DFF_150.Q ;
  assign g320 = \DFF_291.Q ;
  assign g3201 = \DFF_156.Q ;
  assign g3204 = \DFF_159.Q ;
  assign g3207 = \DFF_158.Q ;
  assign g321 = \DFF_294.Q ;
  assign g3210 = \DFF_95.Q ;
  assign g3211 = \DFF_96.Q ;
  assign g322 = \DFF_292.Q ;
  assign g323 = \DFF_293.Q ;
  assign g3235 = \DFF_1635.Q ;
  assign g3236 = \DFF_1632.Q ;
  assign g3237 = \DFF_1630.Q ;
  assign g3238 = \DFF_1631.Q ;
  assign g3239 = \DFF_1628.Q ;
  assign g324 = \DFF_352.Q ;
  assign g3240 = \DFF_1629.Q ;
  assign g3241 = \DFF_1627.Q ;
  assign g3242 = \DFF_1626.Q ;
  assign g3243 = \DFF_1625.Q ;
  assign g3244 = \DFF_1623.Q ;
  assign g3245 = \DFF_1618.Q ;
  assign g3246 = \DFF_1619.Q ;
  assign g3247 = \DFF_1620.Q ;
  assign g3248 = \DFF_1621.Q ;
  assign g3249 = \DFF_1617.Q ;
  assign g325 = \DFF_1504.Q ;
  assign g3250 = \DFF_1616.Q ;
  assign g3251 = \DFF_1615.Q ;
  assign g3252 = \DFF_1614.Q ;
  assign g3253 = g51;
  assign g3254 = \DFF_1429.Q ;
  assign g33 = \DFF_1620.Q ;
  assign g3306 = \DFF_1429.Q ;
  assign g331 = \DFF_1505.Q ;
  assign g3338 = \DFF_1506.Q ;
  assign g3366 = \DFF_1506.Q ;
  assign g337 = \DFF_1506.Q ;
  assign g3398 = \DFF_457.Q ;
  assign g3410 = \DFF_1429.Q ;
  assign g342 = \DFF_329.Q ;
  assign g343 = \DFF_254.Q ;
  assign g346 = \DFF_255.Q ;
  assign g3462 = \DFF_1429.Q ;
  assign g349 = \DFF_330.Q ;
  assign g3494 = \DFF_1506.Q ;
  assign g350 = \DFF_331.Q ;
  assign g351 = \DFF_332.Q ;
  assign g352 = \DFF_333.Q ;
  assign g3522 = \DFF_1506.Q ;
  assign g353 = \DFF_334.Q ;
  assign g354 = \DFF_253.Q ;
  assign g3554 = \DFF_807.Q ;
  assign g3566 = \DFF_1429.Q ;
  assign g357 = \DFF_335.Q ;
  assign g358 = \DFF_257.Q ;
  assign g36 = \DFF_1621.Q ;
  assign g361 = \DFF_258.Q ;
  assign g3618 = \DFF_1429.Q ;
  assign g364 = \DFF_336.Q ;
  assign g365 = \DFF_337.Q ;
  assign g3650 = \DFF_1506.Q ;
  assign g366 = \DFF_338.Q ;
  assign g367 = \DFF_339.Q ;
  assign g3678 = \DFF_1506.Q ;
  assign g368 = \DFF_340.Q ;
  assign g369 = \DFF_256.Q ;
  assign g3710 = \DFF_1157.Q ;
  assign g372 = \DFF_341.Q ;
  assign g3722 = \DFF_1429.Q ;
  assign g373 = \DFF_260.Q ;
  assign g376 = \DFF_261.Q ;
  assign g3774 = \DFF_1429.Q ;
  assign g379 = \DFF_342.Q ;
  assign g380 = \DFF_343.Q ;
  assign g3806 = \DFF_1506.Q ;
  assign g381 = \DFF_344.Q ;
  assign g382 = \DFF_345.Q ;
  assign g383 = \DFF_346.Q ;
  assign g3834 = \DFF_1506.Q ;
  assign g384 = \DFF_259.Q ;
  assign g3866 = \DFF_1507.Q ;
  assign g387 = \DFF_347.Q ;
  assign g3878 = \DFF_19.Q ;
  assign g388 = \DFF_263.Q ;
  assign g39 = \DFF_1617.Q ;
  assign g3900 = \DFF_1613.Q ;
  assign g391 = \DFF_264.Q ;
  assign g394 = \DFF_348.Q ;
  assign g395 = \DFF_349.Q ;
  assign g396 = \DFF_350.Q ;
  assign g397 = \DFF_351.Q ;
  assign g398 = \DFF_262.Q ;
  assign g3993 = \DFF_75.Q ;
  assign g401 = \DFF_1429.Q ;
  assign g402 = \DFF_297.Q ;
  assign g403 = \DFF_295.Q ;
  assign g404 = \DFF_296.Q ;
  assign g405 = \DFF_1428.Q ;
  assign g408 = \DFF_265.Q ;
  assign g4088 = \DFF_67.Q ;
  assign g4090 = \DFF_49.Q ;
  assign g411 = \DFF_266.Q ;
  assign g414 = \DFF_267.Q ;
  assign g417 = \DFF_268.Q ;
  assign g42 = \DFF_1616.Q ;
  assign g420 = \DFF_269.Q ;
  assign g4200 = \DFF_77.Q ;
  assign g423 = \DFF_270.Q ;
  assign g426 = \DFF_273.Q ;
  assign g427 = \DFF_271.Q ;
  assign g428 = \DFF_272.Q ;
  assign g429 = \DFF_274.Q ;
  assign g432 = \DFF_275.Q ;
  assign g4321 = \DFF_69.Q ;
  assign g4323 = \DFF_51.Q ;
  assign g4338 = \DFF_78.Q ;
  assign g4339 = \DFF_76.Q ;
  assign g435 = \DFF_276.Q ;
  assign g438 = \DFF_277.Q ;
  assign g441 = \DFF_278.Q ;
  assign g444 = \DFF_279.Q ;
  assign g4450 = \DFF_79.Q ;
  assign g447 = \DFF_282.Q ;
  assign g448 = \DFF_280.Q ;
  assign g449 = \DFF_281.Q ;
  assign g45 = \DFF_1615.Q ;
  assign g450 = \DFF_298.Q ;
  assign g4507 = \DFF_60.Q ;
  assign g4508 = \DFF_58.Q ;
  assign g451 = \DFF_299.Q ;
  assign g452 = \DFF_300.Q ;
  assign g453 = \DFF_301.Q ;
  assign g454 = \DFF_302.Q ;
  assign g455 = \DFF_383.Q ;
  assign g458 = \DFF_384.Q ;
  assign g4590 = \DFF_53.Q ;
  assign g461 = \DFF_385.Q ;
  assign g464 = \DFF_391.Q ;
  assign g465 = \DFF_392.Q ;
  assign g468 = \DFF_393.Q ;
  assign g4683 = \DFF_44.Q ;
  assign g4684 = \DFF_43.Q ;
  assign g471 = \DFF_394.Q ;
  assign g4735 = \DFF_68.Q ;
  assign g4736 = \DFF_66.Q ;
  assign g474 = \DFF_1427.Q ;
  assign g477 = \DFF_386.Q ;
  assign g478 = \DFF_387.Q ;
  assign g479 = \DFF_388.Q ;
  assign g48 = \DFF_1614.Q ;
  assign g480 = \DFF_389.Q ;
  assign g481 = \DFF_1428.Q ;
  assign g484 = \DFF_390.Q ;
  assign g485 = \DFF_1429.Q ;
  assign g486 = \DFF_380.Q ;
  assign g4860 = \DFF_89.Q ;
  assign g4861 = \DFF_88.Q ;
  assign g487 = \DFF_381.Q ;
  assign g488 = \DFF_382.Q ;
  assign g489 = \DFF_376.Q ;
  assign g490 = \DFF_429.Q ;
  assign g4911 = \DFF_50.Q ;
  assign g4912 = \DFF_48.Q ;
  assign g493 = \DFF_430.Q ;
  assign g496 = \DFF_431.Q ;
  assign g499 = \DFF_402.Q ;
  assign g5 = \DFF_1630.Q ;
  assign g506 = \DFF_432.Q ;
  assign g507 = \DFF_433.Q ;
  assign g5070 = \DFF_39.Q ;
  assign g5071 = \DFF_38.Q ;
  assign g510 = \DFF_361.Q ;
  assign g513 = \DFF_362.Q ;
  assign g5141 = \DFF_74.Q ;
  assign g5199 = \DFF_84.Q ;
  assign g52 = \DFF_245.Q ;
  assign g520 = \DFF_442.Q ;
  assign g5200 = \DFF_83.Q ;
  assign g523 = \DFF_363.Q ;
  assign g5234 = \DFF_56.Q ;
  assign g524 = \DFF_364.Q ;
  assign g525 = \DFF_443.Q ;
  assign g528 = \DFF_395.Q ;
  assign g529 = \DFF_444.Q ;
  assign g5297 = \DFF_42.Q ;
  assign g530 = \DFF_445.Q ;
  assign g531 = \DFF_446.Q ;
  assign g532 = \DFF_447.Q ;
  assign g533 = \DFF_448.Q ;
  assign g5334 = \DFF_87.Q ;
  assign g534 = \DFF_449.Q ;
  assign g535 = \DFF_396.Q ;
  assign g536 = \DFF_450.Q ;
  assign g537 = \DFF_451.Q ;
  assign g538 = \DFF_452.Q ;
  assign g5388 = \DFF_1611.Q ;
  assign g5390 = \DFF_254.Q ;
  assign g5395 = \DFF_255.Q ;
  assign g5396 = \DFF_257.Q ;
  assign g5397 = \DFF_604.Q ;
  assign g5398 = \DFF_258.Q ;
  assign g5399 = \DFF_260.Q ;
  assign g5400 = \DFF_605.Q ;
  assign g5401 = \DFF_607.Q ;
  assign g5402 = \DFF_954.Q ;
  assign g5403 = \DFF_261.Q ;
  assign g5404 = \DFF_263.Q ;
  assign g5405 = \DFF_608.Q ;
  assign g5406 = \DFF_610.Q ;
  assign g5407 = \DFF_955.Q ;
  assign g5408 = \DFF_957.Q ;
  assign g5409 = \DFF_1304.Q ;
  assign g541 = \DFF_453.Q ;
  assign g5411 = \DFF_264.Q ;
  assign g5412 = \DFF_611.Q ;
  assign g5413 = \DFF_613.Q ;
  assign g5414 = \DFF_958.Q ;
  assign g5415 = \DFF_960.Q ;
  assign g5416 = \DFF_1305.Q ;
  assign g5417 = \DFF_1307.Q ;
  assign g5418 = \DFF_614.Q ;
  assign g5419 = \DFF_961.Q ;
  assign g542 = \DFF_397.Q ;
  assign g5420 = \DFF_963.Q ;
  assign g5421 = \DFF_1308.Q ;
  assign g5422 = \DFF_1310.Q ;
  assign g5424 = \DFF_964.Q ;
  assign g5425 = \DFF_1311.Q ;
  assign g5426 = \DFF_1313.Q ;
  assign g5427 = \DFF_1314.Q ;
  assign g543 = \DFF_398.Q ;
  assign g5437 = \DFF_1427.Q ;
  assign g5438 = \DFF_1427.Q ;
  assign g544 = \DFF_399.Q ;
  assign g545 = \DFF_1504.Q ;
  assign g5472 = \DFF_1427.Q ;
  assign g5473 = \DFF_1427.Q ;
  assign g548 = \DFF_400.Q ;
  assign g549 = \DFF_401.Q ;
  assign g550 = \DFF_1506.Q ;
  assign g5508 = \DFF_402.Q ;
  assign g551 = \DFF_1505.Q ;
  assign g5511 = \DFF_1427.Q ;
  assign g5512 = \DFF_1427.Q ;
  assign g554 = \DFF_359.Q ;
  assign g5547 = \DFF_310.D ;
  assign g5548 = \DFF_308.D ;
  assign g5549 = \DFF_1297.Q ;
  assign g5550 = \DFF_1297.Q ;
  assign g5552 = \DFF_752.Q ;
  assign g5555 = \DFF_1427.Q ;
  assign g5556 = \DFF_1427.Q ;
  assign g557 = \DFF_360.Q ;
  assign g558 = \DFF_403.Q ;
  assign g559 = \DFF_404.Q ;
  assign g5593 = \DFF_660.D ;
  assign g5594 = \DFF_658.D ;
  assign g5595 = \DFF_1297.Q ;
  assign g5596 = \DFF_1297.Q ;
  assign g5598 = \DFF_1102.Q ;
  assign g56 = \DFF_244.Q ;
  assign g5610 = \DFF_1010.D ;
  assign g5611 = \DFF_1008.D ;
  assign g5612 = \DFF_1297.Q ;
  assign g5613 = \DFF_1297.Q ;
  assign g5615 = \DFF_1452.Q ;
  assign g562 = g563;
  assign g5626 = \DFF_300.D ;
  assign g5627 = \DFF_298.D ;
  assign g5629 = \DFF_1504.Q ;
  assign g5635 = \DFF_1360.D ;
  assign g5636 = \DFF_1358.D ;
  assign g5637 = \DFF_1297.Q ;
  assign g5638 = \DFF_1297.Q ;
  assign g564 = \DFF_365.Q ;
  assign g5645 = \DFF_310.D ;
  assign g5648 = \DFF_1505.Q ;
  assign g565 = \DFF_372.Q ;
  assign g5654 = \DFF_650.D ;
  assign g5655 = \DFF_648.D ;
  assign g5657 = \DFF_1504.Q ;
  assign g566 = \DFF_373.Q ;
  assign g5665 = \DFF_308.D ;
  assign g567 = \DFF_374.Q ;
  assign g568 = \DFF_375.Q ;
  assign g5683 = \DFF_660.D ;
  assign g5686 = \DFF_1505.Q ;
  assign g569 = \DFF_366.Q ;
  assign g5692 = \DFF_1000.D ;
  assign g5693 = \DFF_998.D ;
  assign g5695 = \DFF_1504.Q ;
  assign g570 = \DFF_367.Q ;
  assign g5701 = g3231;
  assign g5703 = \DFF_306.D ;
  assign g5707 = \DFF_306.D ;
  assign g571 = \DFF_368.Q ;
  assign g5713 = \DFF_72.Q ;
  assign g5717 = \DFF_658.D ;
  assign g572 = \DFF_369.Q ;
  assign g573 = \DFF_370.Q ;
  assign g5735 = \DFF_1010.D ;
  assign g5738 = \DFF_1505.Q ;
  assign g574 = \DFF_371.Q ;
  assign g5744 = \DFF_1350.D ;
  assign g5745 = \DFF_1348.D ;
  assign g5747 = \DFF_1504.Q ;
  assign g5749 = g3212;
  assign g575 = \DFF_407.Q ;
  assign g5752 = \DFF_304.D ;
  assign g576 = \DFF_405.Q ;
  assign g5761 = \DFF_656.D ;
  assign g5765 = \DFF_656.D ;
  assign g577 = \DFF_406.Q ;
  assign g5771 = \DFF_54.Q ;
  assign g5775 = \DFF_1008.D ;
  assign g578 = \DFF_410.Q ;
  assign g579 = \DFF_408.Q ;
  assign g5793 = \DFF_1360.D ;
  assign g5796 = \DFF_1505.Q ;
  assign g5799 = g3221;
  assign g580 = \DFF_409.Q ;
  assign g5800 = g3227;
  assign g5801 = g3216;
  assign g5803 = \DFF_302.D ;
  assign g581 = \DFF_413.Q ;
  assign g5811 = \DFF_654.D ;
  assign g582 = \DFF_411.Q ;
  assign g5820 = \DFF_1006.D ;
  assign g5824 = \DFF_1006.D ;
  assign g583 = \DFF_412.Q ;
  assign g5830 = \DFF_41.Q ;
  assign g5834 = \DFF_1358.D ;
  assign g584 = \DFF_416.Q ;
  assign g5849 = g3228;
  assign g585 = \DFF_414.Q ;
  assign g5850 = g3217;
  assign g5852 = \DFF_300.D ;
  assign g5856 = \DFF_80.Q ;
  assign g5859 = \DFF_652.D ;
  assign g586 = \DFF_415.Q ;
  assign g5867 = \DFF_1004.D ;
  assign g587 = \DFF_417.Q ;
  assign g5876 = \DFF_1356.D ;
  assign g5880 = \DFF_1356.D ;
  assign g5886 = \DFF_86.Q ;
  assign g5889 = g3219;
  assign g5893 = \DFF_298.D ;
  assign g5899 = \DFF_650.D ;
  assign g590 = \DFF_418.Q ;
  assign g5903 = \DFF_62.Q ;
  assign g5906 = \DFF_1002.D ;
  assign g5914 = \DFF_1354.D ;
  assign g5922 = g3234;
  assign g5923 = g3223;
  assign g5924 = g3218;
  assign g593 = \DFF_419.Q ;
  assign g5932 = \DFF_648.D ;
  assign g5938 = \DFF_1000.D ;
  assign g5942 = \DFF_45.Q ;
  assign g5945 = \DFF_1352.D ;
  assign g5951 = g3233;
  assign g5952 = g3222;
  assign g5953 = \DFF_312.D ;
  assign g5958 = \DFF_70.Q ;
  assign g596 = \DFF_420.Q ;
  assign g5966 = \DFF_998.D ;
  assign g5972 = \DFF_1350.D ;
  assign g5976 = \DFF_90.Q ;
  assign g5978 = g3230;
  assign g5979 = g3224;
  assign g5982 = \DFF_662.D ;
  assign g5987 = \DFF_52.Q ;
  assign g599 = \DFF_421.Q ;
  assign g5995 = \DFF_1348.D ;
  assign g6000 = \DFF_1563.Q ;
  assign g6014 = g3225;
  assign g6015 = g3213;
  assign g6019 = \DFF_1012.D ;
  assign g602 = \DFF_422.Q ;
  assign g6024 = \DFF_40.Q ;
  assign g6029 = g3226;
  assign g6030 = g3214;
  assign g6031 = \DFF_394.Q ;
  assign g6035 = \DFF_1362.D ;
  assign g6040 = \DFF_85.Q ;
  assign g6041 = g3215;
  assign g6042 = \DFF_744.Q ;
  assign g6046 = \DFF_1094.Q ;
  assign g6048 = \DFF_158.Q ;
  assign g605 = \DFF_426.Q ;
  assign g6051 = \DFF_253.Q ;
  assign g6052 = \DFF_1444.Q ;
  assign g6053 = \DFF_256.Q ;
  assign g6054 = \DFF_383.Q ;
  assign g6055 = \DFF_603.Q ;
  assign g6056 = \DFF_259.Q ;
  assign g6057 = \DFF_384.Q ;
  assign g6058 = \DFF_606.Q ;
  assign g6059 = \DFF_733.Q ;
  assign g6060 = \DFF_953.Q ;
  assign g6061 = \DFF_262.Q ;
  assign g6062 = \DFF_385.Q ;
  assign g6063 = \DFF_609.Q ;
  assign g6064 = \DFF_734.Q ;
  assign g6065 = \DFF_956.Q ;
  assign g6066 = \DFF_1083.Q ;
  assign g6067 = \DFF_1303.Q ;
  assign g6079 = \DFF_392.Q ;
  assign g608 = \DFF_427.Q ;
  assign g6080 = \DFF_612.Q ;
  assign g6081 = \DFF_735.Q ;
  assign g6082 = \DFF_959.Q ;
  assign g6083 = \DFF_1084.Q ;
  assign g6084 = \DFF_1306.Q ;
  assign g6085 = \DFF_1433.Q ;
  assign g6086 = \DFF_393.Q ;
  assign g6098 = \DFF_742.Q ;
  assign g6099 = \DFF_962.Q ;
  assign g61 = \DFF_243.Q ;
  assign g6100 = \DFF_1085.Q ;
  assign g6101 = \DFF_1309.Q ;
  assign g6102 = \DFF_1434.Q ;
  assign g6103 = \DFF_743.Q ;
  assign g611 = \DFF_428.Q ;
  assign g6115 = \DFF_1092.Q ;
  assign g6116 = \DFF_1312.Q ;
  assign g6117 = \DFF_1435.Q ;
  assign g6118 = \DFF_1093.Q ;
  assign g6130 = \DFF_1442.Q ;
  assign g6131 = \DFF_158.Q ;
  assign g6134 = \DFF_1443.Q ;
  assign g6135 = \DFF_443.Q ;
  assign g6139 = g3220;
  assign g614 = \DFF_423.Q ;
  assign g6145 = \DFF_793.Q ;
  assign g6153 = \DFF_159.Q ;
  assign g6156 = g3232;
  assign g6166 = \DFF_1143.Q ;
  assign g617 = \DFF_424.Q ;
  assign g6183 = \DFF_453.D ;
  assign g6193 = \DFF_1493.Q ;
  assign g620 = \DFF_425.Q ;
  assign g6204 = \DFF_451.D ;
  assign g6215 = \DFF_803.D ;
  assign g6225 = \DFF_55.Q ;
  assign g623 = \DFF_1504.Q ;
  assign g6230 = g3229;
  assign g6231 = \DFF_1427.Q ;
  assign g6232 = \DFF_1427.Q ;
  assign g626 = \DFF_1505.Q ;
  assign g6288 = \DFF_450.D ;
  assign g629 = \DFF_1506.Q ;
  assign g6293 = \DFF_801.D ;
  assign g630 = \DFF_457.Q ;
  assign g6304 = \DFF_1153.D ;
  assign g6313 = \DFF_1428.Q ;
  assign g6314 = \DFF_1428.Q ;
  assign g633 = \DFF_460.Q ;
  assign g6367 = \DFF_449.D ;
  assign g6368 = \DFF_1427.Q ;
  assign g6369 = \DFF_1427.Q ;
  assign g640 = \DFF_459.Q ;
  assign g6425 = \DFF_800.D ;
  assign g6430 = \DFF_1151.D ;
  assign g6441 = \DFF_1503.D ;
  assign g6442 = \DFF_57.Q ;
  assign g6447 = \DFF_1428.Q ;
  assign g6448 = \DFF_1428.Q ;
  assign g646 = \DFF_462.Q ;
  assign g6485 = \DFF_1504.Q ;
  assign g6486 = \DFF_1504.Q ;
  assign g65 = \DFF_242.Q ;
  assign g6517 = \DFF_448.D ;
  assign g6518 = \DFF_1428.Q ;
  assign g6519 = \DFF_1428.Q ;
  assign g653 = \DFF_461.Q ;
  assign g6572 = \DFF_799.D ;
  assign g6573 = \DFF_1427.Q ;
  assign g6574 = \DFF_1427.Q ;
  assign g659 = \DFF_458.Q ;
  assign g660 = \DFF_463.Q ;
  assign g6630 = \DFF_1150.D ;
  assign g6635 = \DFF_1501.D ;
  assign g6636 = \DFF_1004.D ;
  assign g6641 = \DFF_304.D ;
  assign g6642 = \DFF_1505.Q ;
  assign g6643 = \DFF_1505.Q ;
  assign g666 = \DFF_465.Q ;
  assign g6677 = \DFF_1504.Q ;
  assign g6678 = \DFF_1504.Q ;
  assign g6711 = \DFF_447.D ;
  assign g6712 = \DFF_1428.Q ;
  assign g6713 = \DFF_1428.Q ;
  assign g672 = \DFF_464.Q ;
  assign g6750 = \DFF_1504.Q ;
  assign g6751 = \DFF_1504.Q ;
  assign g6781 = \DFF_798.D ;
  assign g6782 = \DFF_1428.Q ;
  assign g6783 = \DFF_1428.Q ;
  assign g679 = \DFF_466.Q ;
  assign g6836 = \DFF_1149.D ;
  assign g6837 = \DFF_1427.Q ;
  assign g6838 = \DFF_1427.Q ;
  assign g686 = \DFF_467.Q ;
  assign g6894 = \DFF_1500.D ;
  assign g6895 = \DFF_59.Q ;
  assign g6897 = \DFF_1006.D ;
  assign g6911 = \DFF_1505.Q ;
  assign g6912 = \DFF_1505.Q ;
  assign g692 = \DFF_468.Q ;
  assign g6942 = \DFF_446.D ;
  assign g6943 = \DFF_654.D ;
  assign g6944 = \DFF_1505.Q ;
  assign g6945 = \DFF_1505.Q ;
  assign g6979 = \DFF_1504.Q ;
  assign g698 = \DFF_471.Q ;
  assign g6980 = \DFF_1504.Q ;
  assign g699 = \DFF_469.Q ;
  assign g70 = \DFF_241.Q ;
  assign g700 = \DFF_470.Q ;
  assign g701 = \DFF_474.Q ;
  assign g7013 = \DFF_797.D ;
  assign g7014 = \DFF_1428.Q ;
  assign g7015 = \DFF_1428.Q ;
  assign g702 = \DFF_472.Q ;
  assign g703 = \DFF_473.Q ;
  assign g704 = \DFF_477.Q ;
  assign g705 = \DFF_475.Q ;
  assign g7052 = \DFF_1504.Q ;
  assign g7053 = \DFF_1504.Q ;
  assign g706 = \DFF_476.Q ;
  assign g707 = \DFF_480.Q ;
  assign g708 = \DFF_478.Q ;
  assign g7083 = \DFF_1148.D ;
  assign g7084 = \DFF_1428.Q ;
  assign g7085 = \DFF_1428.Q ;
  assign g709 = \DFF_479.Q ;
  assign g710 = \DFF_483.Q ;
  assign g711 = \DFF_481.Q ;
  assign g712 = \DFF_482.Q ;
  assign g713 = \DFF_486.Q ;
  assign g7138 = \DFF_1499.D ;
  assign g7139 = \DFF_1008.D ;
  assign g714 = \DFF_484.Q ;
  assign g7140 = \DFF_1360.D ;
  assign g7141 = \DFF_1350.D ;
  assign g715 = \DFF_485.Q ;
  assign g7157 = \DFF_445.D ;
  assign g716 = \DFF_489.Q ;
  assign g7161 = \DFF_1505.Q ;
  assign g7162 = \DFF_1505.Q ;
  assign g717 = \DFF_487.Q ;
  assign g718 = \DFF_488.Q ;
  assign g719 = \DFF_492.Q ;
  assign g7192 = \DFF_796.D ;
  assign g7193 = \DFF_1004.D ;
  assign g7194 = \DFF_1505.Q ;
  assign g7195 = \DFF_1505.Q ;
  assign g720 = \DFF_490.Q ;
  assign g721 = \DFF_491.Q ;
  assign g722 = \DFF_495.Q ;
  assign g7229 = \DFF_1504.Q ;
  assign g723 = \DFF_493.Q ;
  assign g7230 = \DFF_1504.Q ;
  assign g724 = \DFF_494.Q ;
  assign g725 = \DFF_498.Q ;
  assign g726 = \DFF_496.Q ;
  assign g7263 = \DFF_1147.D ;
  assign g7264 = \DFF_1428.Q ;
  assign g7265 = \DFF_1428.Q ;
  assign g727 = \DFF_497.Q ;
  assign g728 = \DFF_501.Q ;
  assign g729 = \DFF_499.Q ;
  assign g730 = \DFF_500.Q ;
  assign g7302 = \DFF_1504.Q ;
  assign g7303 = \DFF_1504.Q ;
  assign g731 = \DFF_504.Q ;
  assign g732 = \DFF_502.Q ;
  assign g733 = \DFF_503.Q ;
  assign g7333 = \DFF_1498.D ;
  assign g7334 = \DFF_61.Q ;
  assign g7336 = \DFF_1010.D ;
  assign g7337 = \DFF_1352.D ;
  assign g734 = \DFF_507.Q ;
  assign g7346 = \DFF_312.D ;
  assign g7348 = \DFF_444.D ;
  assign g735 = \DFF_505.Q ;
  assign g7353 = \DFF_795.D ;
  assign g7357 = \DFF_1505.Q ;
  assign g7358 = \DFF_1505.Q ;
  assign g736 = \DFF_506.Q ;
  assign g737 = \DFF_510.Q ;
  assign g738 = \DFF_508.Q ;
  assign g7388 = \DFF_1146.D ;
  assign g7389 = \DFF_1354.D ;
  assign g739 = \DFF_509.Q ;
  assign g7390 = \DFF_1505.Q ;
  assign g7391 = \DFF_1505.Q ;
  assign g74 = \DFF_240.Q ;
  assign g740 = \DFF_595.Q ;
  assign g7425 = \DFF_1504.Q ;
  assign g7426 = \DFF_1504.Q ;
  assign g744 = \DFF_594.Q ;
  assign g7459 = \DFF_1497.D ;
  assign g7460 = \DFF_1012.D ;
  assign g7461 = \DFF_1358.D ;
  assign g7476 = \DFF_662.D ;
  assign g7478 = \DFF_794.D ;
  assign g7483 = \DFF_1145.D ;
  assign g7487 = \DFF_1505.Q ;
  assign g7488 = \DFF_1505.Q ;
  assign g749 = \DFF_593.Q ;
  assign g7518 = \DFF_1496.D ;
  assign g7519 = \DFF_63.Q ;
  assign g7521 = \DFF_1348.D ;
  assign g753 = \DFF_592.Q ;
  assign g7532 = \DFF_1012.D ;
  assign g7534 = \DFF_1144.D ;
  assign g7539 = \DFF_1495.D ;
  assign g7540 = \DFF_998.D ;
  assign g7541 = \DFF_1356.D ;
  assign g7554 = \DFF_302.D ;
  assign g7558 = \DFF_1362.D ;
  assign g7560 = \DFF_1494.D ;
  assign g7561 = \DFF_1000.D ;
  assign g7577 = \DFF_652.D ;
  assign g758 = \DFF_591.Q ;
  assign g7581 = \DFF_1002.D ;
  assign g7582 = \DFF_1354.D ;
  assign g7591 = \DFF_1002.D ;
  assign g7594 = \DFF_1362.D ;
  assign g7606 = \DFF_1352.D ;
  assign g762 = \DFF_590.Q ;
  assign g767 = \DFF_589.Q ;
  assign g771 = \DFF_588.Q ;
  assign g776 = \DFF_587.Q ;
  assign g780 = \DFF_586.Q ;
  assign g785 = \DFF_62.Q ;
  assign g789 = \DFF_60.Q ;
  assign g79 = \DFF_239.Q ;
  assign g7901 = \DFF_157.Q ;
  assign g7909 = \DFF_1427.Q ;
  assign g7911 = \DFF_402.Q ;
  assign g793 = \DFF_58.Q ;
  assign g7936 = \DFF_3.Q ;
  assign g7956 = \DFF_1428.Q ;
  assign g7961 = \DFF_1427.Q ;
  assign g7963 = \DFF_752.Q ;
  assign g797 = \DFF_56.Q ;
  assign g7976 = \DFF_1506.Q ;
  assign g8 = \DFF_1631.Q ;
  assign g8007 = \DFF_1428.Q ;
  assign g801 = \DFF_54.Q ;
  assign g8012 = \DFF_1427.Q ;
  assign g8014 = \DFF_1102.Q ;
  assign g8021 = \DFF_17.Q ;
  assign g8023 = \DFF_71.Q ;
  assign g8030 = \DFF_1505.Q ;
  assign g8031 = \DFF_1505.Q ;
  assign g805 = \DFF_52.Q ;
  assign g8082 = \DFF_1428.Q ;
  assign g8087 = \DFF_1427.Q ;
  assign g8089 = \DFF_1452.Q ;
  assign g809 = \DFF_50.Q ;
  assign g8096 = \DFF_81.Q ;
  assign g8106 = \DFF_1504.Q ;
  assign g8107 = \DFF_1504.Q ;
  assign g813 = \DFF_48.Q ;
  assign g8167 = \DFF_1428.Q ;
  assign g817 = \DFF_516.Q ;
  assign g8175 = \DFF_73.Q ;
  assign g818 = \DFF_514.Q ;
  assign g819 = \DFF_515.Q ;
  assign g820 = \DFF_519.Q ;
  assign g821 = \DFF_517.Q ;
  assign g822 = \DFF_518.Q ;
  assign g823 = \DFF_1428.Q ;
  assign g8249 = \DFF_65.Q ;
  assign g8251 = \DFF_47.Q ;
  assign g8258 = \DFF_1635.Q ;
  assign g8259 = \DFF_1632.Q ;
  assign g826 = \DFF_1427.Q ;
  assign g8260 = \DFF_1630.Q ;
  assign g8261 = \DFF_1631.Q ;
  assign g8262 = \DFF_1628.Q ;
  assign g8263 = \DFF_1629.Q ;
  assign g8264 = \DFF_1627.Q ;
  assign g8265 = \DFF_1626.Q ;
  assign g8266 = \DFF_1625.Q ;
  assign g8267 = \DFF_1623.Q ;
  assign g8268 = \DFF_1618.Q ;
  assign g8269 = \DFF_1619.Q ;
  assign g8270 = \DFF_1620.Q ;
  assign g8271 = \DFF_1621.Q ;
  assign g8272 = \DFF_1617.Q ;
  assign g8273 = \DFF_1616.Q ;
  assign g8274 = \DFF_1615.Q ;
  assign g8275 = \DFF_1614.Q ;
  assign g8277 = \DFF_317.Q ;
  assign g8278 = \DFF_1302.Q ;
  assign g8284 = \DFF_402.Q ;
  assign g8285 = \DFF_402.Q ;
  assign g8286 = \DFF_667.Q ;
  assign g8287 = \DFF_1302.Q ;
  assign g829 = \DFF_522.Q ;
  assign g8293 = \DFF_752.Q ;
  assign g8294 = \DFF_752.Q ;
  assign g8295 = \DFF_1017.Q ;
  assign g8296 = \DFF_1302.Q ;
  assign g83 = \DFF_238.Q ;
  assign g830 = \DFF_520.Q ;
  assign g8302 = \DFF_1102.Q ;
  assign g8303 = \DFF_1102.Q ;
  assign g8304 = \DFF_1367.Q ;
  assign g8305 = \DFF_1302.Q ;
  assign g831 = \DFF_521.Q ;
  assign g8311 = \DFF_1452.Q ;
  assign g8312 = \DFF_1452.Q ;
  assign g8313 = \DFF_3.Q ;
  assign g8317 = \DFF_1563.Q ;
  assign g832 = \DFF_525.Q ;
  assign g8321 = \DFF_1429.Q ;
  assign g8324 = \DFF_1428.Q ;
  assign g833 = \DFF_523.Q ;
  assign g8330 = \DFF_1429.Q ;
  assign g8333 = \DFF_1428.Q ;
  assign g8336 = \DFF_1427.Q ;
  assign g834 = \DFF_524.Q ;
  assign g8341 = \DFF_1429.Q ;
  assign g8344 = \DFF_1428.Q ;
  assign g8347 = \DFF_1427.Q ;
  assign g835 = \DFF_528.Q ;
  assign g8351 = \DFF_1429.Q ;
  assign g8354 = \DFF_1428.Q ;
  assign g8357 = \DFF_1428.Q ;
  assign g836 = \DFF_526.Q ;
  assign g8363 = \DFF_1427.Q ;
  assign g8366 = \DFF_1429.Q ;
  assign g8369 = \DFF_1428.Q ;
  assign g837 = \DFF_527.Q ;
  assign g8372 = \DFF_1427.Q ;
  assign g8375 = \DFF_1428.Q ;
  assign g838 = \DFF_531.Q ;
  assign g8382 = \DFF_1429.Q ;
  assign g8388 = \DFF_1429.Q ;
  assign g839 = \DFF_529.Q ;
  assign g8391 = \DFF_1428.Q ;
  assign g8397 = \DFF_1429.Q ;
  assign g840 = \DFF_530.Q ;
  assign g8400 = \DFF_1428.Q ;
  assign g8403 = \DFF_1427.Q ;
  assign g8408 = \DFF_1429.Q ;
  assign g841 = \DFF_534.Q ;
  assign g8411 = \DFF_1428.Q ;
  assign g8414 = \DFF_1427.Q ;
  assign g8418 = \DFF_1429.Q ;
  assign g842 = \DFF_532.Q ;
  assign g8421 = \DFF_1428.Q ;
  assign g8424 = \DFF_1428.Q ;
  assign g843 = \DFF_533.Q ;
  assign g8434 = \DFF_1429.Q ;
  assign g844 = \DFF_537.Q ;
  assign g8440 = \DFF_1429.Q ;
  assign g8443 = \DFF_1428.Q ;
  assign g8449 = \DFF_1429.Q ;
  assign g845 = \DFF_535.Q ;
  assign g8452 = \DFF_1428.Q ;
  assign g8455 = \DFF_1427.Q ;
  assign g846 = \DFF_536.Q ;
  assign g8460 = \DFF_1429.Q ;
  assign g8469 = \DFF_1429.Q ;
  assign g847 = \DFF_540.Q ;
  assign g8475 = \DFF_1429.Q ;
  assign g8478 = \DFF_1428.Q ;
  assign g848 = \DFF_538.Q ;
  assign g849 = \DFF_539.Q ;
  assign g8494 = \DFF_1429.Q ;
  assign g850 = \DFF_543.Q ;
  assign g851 = \DFF_541.Q ;
  assign g852 = \DFF_542.Q ;
  assign g853 = \DFF_1429.Q ;
  assign g856 = \DFF_546.Q ;
  assign g8569 = \DFF_1563.Q ;
  assign g857 = \DFF_544.Q ;
  assign g8575 = \DFF_1563.Q ;
  assign g8578 = \DFF_1563.Q ;
  assign g8579 = \DFF_1563.Q ;
  assign g858 = \DFF_545.Q ;
  assign g8580 = \DFF_361.Q ;
  assign g8587 = \DFF_711.Q ;
  assign g859 = \DFF_549.Q ;
  assign g8594 = \DFF_1061.Q ;
  assign g860 = \DFF_547.Q ;
  assign g8602 = \DFF_1506.Q ;
  assign g8605 = \DFF_1411.Q ;
  assign g861 = \DFF_548.Q ;
  assign g8614 = \DFF_1506.Q ;
  assign g8617 = \DFF_1504.Q ;
  assign g862 = \DFF_552.Q ;
  assign g8620 = \DFF_1297.Q ;
  assign g8622 = \DFF_1506.Q ;
  assign g8627 = \DFF_1506.Q ;
  assign g863 = \DFF_550.Q ;
  assign g8630 = \DFF_1297.Q ;
  assign g8632 = \DFF_1506.Q ;
  assign g8637 = \DFF_1506.Q ;
  assign g864 = \DFF_551.Q ;
  assign g8640 = \DFF_1505.Q ;
  assign g8643 = \DFF_1506.Q ;
  assign g8646 = \DFF_1506.Q ;
  assign g8649 = \DFF_1297.Q ;
  assign g865 = \DFF_555.Q ;
  assign g8651 = \DFF_1506.Q ;
  assign g8655 = \DFF_19.Q ;
  assign g8658 = \DFF_298.D ;
  assign g8659 = \DFF_1506.Q ;
  assign g866 = \DFF_553.Q ;
  assign g8662 = \DFF_1506.Q ;
  assign g8665 = \DFF_1297.Q ;
  assign g8667 = \DFF_1506.Q ;
  assign g867 = \DFF_554.Q ;
  assign g8670 = \DFF_19.Q ;
  assign g8673 = \DFF_1506.Q ;
  assign g8677 = \DFF_648.D ;
  assign g8678 = \DFF_1506.Q ;
  assign g868 = \DFF_1296.Q ;
  assign g8681 = \DFF_1506.Q ;
  assign g8684 = \DFF_19.Q ;
  assign g8689 = \DFF_998.D ;
  assign g869 = \DFF_1302.Q ;
  assign g8690 = \DFF_1506.Q ;
  assign g8693 = \DFF_1506.Q ;
  assign g8696 = \DFF_19.Q ;
  assign g8699 = \DFF_300.D ;
  assign g870 = \DFF_1297.Q ;
  assign g8700 = \DFF_1504.Q ;
  assign g8707 = \DFF_1348.D ;
  assign g8708 = \DFF_19.Q ;
  assign g8711 = \DFF_19.Q ;
  assign g8714 = \DFF_1505.Q ;
  assign g8718 = \DFF_650.D ;
  assign g8719 = \DFF_1504.Q ;
  assign g873 = \DFF_556.Q ;
  assign g8745 = \DFF_19.Q ;
  assign g8748 = \DFF_1506.Q ;
  assign g8752 = \DFF_1505.Q ;
  assign g8756 = \DFF_1000.D ;
  assign g8757 = \DFF_1504.Q ;
  assign g876 = \DFF_557.Q ;
  assign g8763 = \DFF_19.Q ;
  assign g8766 = \DFF_19.Q ;
  assign g8769 = \DFF_253.Q ;
  assign g8770 = \DFF_302.D ;
  assign g8771 = \DFF_1506.Q ;
  assign g8775 = \DFF_1505.Q ;
  assign g8779 = \DFF_1350.D ;
  assign g8780 = \DFF_1504.Q ;
  assign g8785 = \DFF_19.Q ;
  assign g8788 = \DFF_19.Q ;
  assign g879 = \DFF_558.Q ;
  assign g8791 = \DFF_256.Q ;
  assign g8792 = \DFF_603.Q ;
  assign g8793 = \DFF_652.D ;
  assign g8794 = \DFF_1506.Q ;
  assign g8798 = \DFF_1505.Q ;
  assign g88 = \DFF_237.Q ;
  assign g8802 = \DFF_19.Q ;
  assign g8805 = \DFF_19.Q ;
  assign g8808 = \DFF_254.Q ;
  assign g8809 = \DFF_259.Q ;
  assign g8810 = \DFF_606.Q ;
  assign g8811 = \DFF_953.Q ;
  assign g8812 = \DFF_1002.D ;
  assign g8813 = \DFF_1506.Q ;
  assign g8817 = \DFF_19.Q ;
  assign g882 = \DFF_562.Q ;
  assign g8820 = \DFF_257.Q ;
  assign g8821 = \DFF_262.Q ;
  assign g8822 = \DFF_443.Q ;
  assign g8823 = \DFF_1504.Q ;
  assign g8824 = \DFF_604.Q ;
  assign g8825 = \DFF_609.Q ;
  assign g8826 = \DFF_956.Q ;
  assign g8827 = \DFF_1303.Q ;
  assign g8828 = \DFF_1352.D ;
  assign g8829 = \DFF_19.Q ;
  assign g8832 = \DFF_1613.Q ;
  assign g8835 = \DFF_3.Q ;
  assign g8836 = \DFF_1427.Q ;
  assign g8839 = \DFF_255.Q ;
  assign g8840 = \DFF_260.Q ;
  assign g8843 = \DFF_393.Q ;
  assign g8844 = \DFF_607.Q ;
  assign g8845 = \DFF_612.Q ;
  assign g8846 = \DFF_793.Q ;
  assign g8847 = \DFF_1504.Q ;
  assign g885 = \DFF_563.Q ;
  assign g8850 = \DFF_954.Q ;
  assign g8851 = \DFF_959.Q ;
  assign g8852 = \DFF_1306.Q ;
  assign g8853 = \DFF_19.Q ;
  assign g8856 = \DFF_1428.Q ;
  assign g8859 = \DFF_258.Q ;
  assign g8860 = \DFF_263.Q ;
  assign g8862 = \DFF_3.Q ;
  assign g8863 = \DFF_1427.Q ;
  assign g8866 = \DFF_605.Q ;
  assign g8867 = \DFF_610.Q ;
  assign g8870 = \DFF_743.Q ;
  assign g8871 = \DFF_957.Q ;
  assign g8872 = \DFF_962.Q ;
  assign g8873 = \DFF_1143.Q ;
  assign g8874 = \DFF_1504.Q ;
  assign g8877 = \DFF_1304.Q ;
  assign g8878 = \DFF_1309.Q ;
  assign g8879 = \DFF_19.Q ;
  assign g888 = \DFF_564.Q ;
  assign g8882 = \DFF_1613.Q ;
  assign g8885 = \DFF_1429.Q ;
  assign g8888 = \DFF_1427.Q ;
  assign g8891 = \DFF_261.Q ;
  assign g8893 = \DFF_394.Q ;
  assign g8894 = \DFF_1428.Q ;
  assign g8897 = \DFF_608.Q ;
  assign g8898 = \DFF_613.Q ;
  assign g8900 = \DFF_3.Q ;
  assign g8901 = \DFF_1427.Q ;
  assign g8904 = \DFF_955.Q ;
  assign g8905 = \DFF_960.Q ;
  assign g8908 = \DFF_1093.Q ;
  assign g8909 = \DFF_1307.Q ;
  assign g891 = \DFF_568.Q ;
  assign g8910 = \DFF_1312.Q ;
  assign g8911 = \DFF_1493.Q ;
  assign g8912 = \DFF_1504.Q ;
  assign g8915 = \DFF_19.Q ;
  assign g8918 = \DFF_1428.Q ;
  assign g8921 = \DFF_1427.Q ;
  assign g8924 = \DFF_264.Q ;
  assign g8925 = \DFF_1429.Q ;
  assign g8928 = \DFF_1427.Q ;
  assign g8931 = \DFF_611.Q ;
  assign g8933 = \DFF_744.Q ;
  assign g8934 = \DFF_1428.Q ;
  assign g8937 = \DFF_958.Q ;
  assign g8938 = \DFF_963.Q ;
  assign g894 = \DFF_569.Q ;
  assign g8940 = \DFF_3.Q ;
  assign g8941 = \DFF_1427.Q ;
  assign g8944 = \DFF_1305.Q ;
  assign g8945 = \DFF_1310.Q ;
  assign g8948 = \DFF_1443.Q ;
  assign g8949 = \DFF_1613.Q ;
  assign g8952 = \DFF_1429.Q ;
  assign g8955 = \DFF_1428.Q ;
  assign g8958 = \DFF_1428.Q ;
  assign g8961 = \DFF_1427.Q ;
  assign g8964 = \DFF_614.Q ;
  assign g8965 = \DFF_1429.Q ;
  assign g8968 = \DFF_1427.Q ;
  assign g897 = \DFF_570.Q ;
  assign g8971 = \DFF_961.Q ;
  assign g8973 = \DFF_1094.Q ;
  assign g8974 = \DFF_1428.Q ;
  assign g8977 = \DFF_1308.Q ;
  assign g8978 = \DFF_1313.Q ;
  assign g8980 = \DFF_1429.Q ;
  assign g8984 = \DFF_1429.Q ;
  assign g8987 = \DFF_1428.Q ;
  assign g8990 = \DFF_1428.Q ;
  assign g8993 = \DFF_1427.Q ;
  assign g8996 = \DFF_964.Q ;
  assign g8997 = \DFF_1429.Q ;
  assign g900 = \DFF_574.Q ;
  assign g9000 = \DFF_1427.Q ;
  assign g9003 = \DFF_1311.Q ;
  assign g9005 = \DFF_1444.Q ;
  assign g9006 = \DFF_1613.Q ;
  assign g9010 = \DFF_1429.Q ;
  assign g9013 = \DFF_1429.Q ;
  assign g9016 = \DFF_1428.Q ;
  assign g9019 = \DFF_1428.Q ;
  assign g9022 = \DFF_1427.Q ;
  assign g9025 = \DFF_1314.Q ;
  assign g9027 = \DFF_432.Q ;
  assign g903 = \DFF_575.Q ;
  assign g9035 = \DFF_1429.Q ;
  assign g9038 = \DFF_1429.Q ;
  assign g9041 = \DFF_1428.Q ;
  assign g9044 = \DFF_1613.Q ;
  assign g9050 = \DFF_782.Q ;
  assign g9058 = \DFF_1429.Q ;
  assign g906 = \DFF_576.Q ;
  assign g9067 = \DFF_1132.Q ;
  assign g9084 = \DFF_1482.Q ;
  assign g909 = \DFF_580.Q ;
  assign g912 = \DFF_581.Q ;
  assign g9128 = \DFF_1506.Q ;
  assign g9134 = \DFF_1506.Q ;
  assign g9140 = \DFF_1506.Q ;
  assign g9146 = \DFF_1506.Q ;
  assign g9149 = \DFF_3.Q ;
  assign g915 = \DFF_582.Q ;
  assign g9150 = \DFF_66.Q ;
  assign g9159 = \DFF_3.Q ;
  assign g9160 = \DFF_108.Q ;
  assign g9161 = \DFF_68.Q ;
  assign g9170 = \DFF_1427.Q ;
  assign g9173 = \DFF_1563.Q ;
  assign g9174 = \DFF_48.Q ;
  assign g918 = \DFF_559.Q ;
  assign g9183 = \DFF_3.Q ;
  assign g9184 = \DFF_157.Q ;
  assign g9187 = \DFF_70.Q ;
  assign g9196 = \DFF_1428.Q ;
  assign g9199 = \DFF_1427.Q ;
  assign g92 = \DFF_236.Q ;
  assign g9202 = \DFF_1563.Q ;
  assign g9203 = \DFF_50.Q ;
  assign g921 = \DFF_560.Q ;
  assign g9212 = \DFF_1427.Q ;
  assign g9215 = \DFF_1563.Q ;
  assign g9216 = \DFF_38.Q ;
  assign g9225 = \DFF_3.Q ;
  assign g9226 = \DFF_97.Q ;
  assign g9227 = \DFF_101.Q ;
  assign g9228 = \DFF_105.Q ;
  assign g9229 = \DFF_157.Q ;
  assign g9232 = \DFF_72.Q ;
  assign g924 = \DFF_561.Q ;
  assign g9242 = \DFF_1429.Q ;
  assign g9245 = \DFF_1428.Q ;
  assign g9248 = \DFF_52.Q ;
  assign g9257 = \DFF_1428.Q ;
  assign g9260 = \DFF_1427.Q ;
  assign g9263 = \DFF_1563.Q ;
  assign g9264 = \DFF_39.Q ;
  assign g927 = \DFF_565.Q ;
  assign g9273 = \DFF_1427.Q ;
  assign g9276 = \DFF_1563.Q ;
  assign g9277 = \DFF_83.Q ;
  assign g9286 = \DFF_109.Q ;
  assign g9287 = \DFF_113.Q ;
  assign g9288 = \DFF_117.Q ;
  assign g9289 = \DFF_118.Q ;
  assign g9290 = \DFF_157.Q ;
  assign g9293 = \DFF_74.Q ;
  assign g930 = \DFF_566.Q ;
  assign g9303 = \DFF_1429.Q ;
  assign g9306 = \DFF_1427.Q ;
  assign g9309 = \DFF_383.Q ;
  assign g9310 = \DFF_54.Q ;
  assign g9320 = \DFF_1429.Q ;
  assign g9323 = \DFF_1428.Q ;
  assign g9326 = \DFF_40.Q ;
  assign g933 = \DFF_567.Q ;
  assign g9335 = \DFF_1428.Q ;
  assign g9338 = \DFF_1427.Q ;
  assign g9341 = \DFF_1563.Q ;
  assign g9342 = \DFF_84.Q ;
  assign g9351 = \DFF_1427.Q ;
  assign g9354 = \DFF_1563.Q ;
  assign g9355 = \DFF_104.Q ;
  assign g9356 = \DFF_76.Q ;
  assign g936 = \DFF_571.Q ;
  assign g9368 = \DFF_1428.Q ;
  assign g9371 = \DFF_1427.Q ;
  assign g9374 = \DFF_56.Q ;
  assign g9384 = \DFF_1429.Q ;
  assign g9387 = \DFF_1427.Q ;
  assign g939 = \DFF_572.Q ;
  assign g9390 = \DFF_733.Q ;
  assign g9391 = \DFF_41.Q ;
  assign g9401 = \DFF_1429.Q ;
  assign g9404 = \DFF_1428.Q ;
  assign g9407 = \DFF_85.Q ;
  assign g9416 = \DFF_1428.Q ;
  assign g9419 = \DFF_1427.Q ;
  assign g942 = \DFF_573.Q ;
  assign g9422 = \DFF_1563.Q ;
  assign g9423 = \DFF_95.Q ;
  assign g9424 = \DFF_98.Q ;
  assign g9425 = \DFF_116.Q ;
  assign g9426 = \DFF_100.Q ;
  assign g9427 = \DFF_78.Q ;
  assign g9443 = \DFF_1429.Q ;
  assign g9446 = \DFF_1428.Q ;
  assign g9449 = \DFF_384.Q ;
  assign g945 = \DFF_577.Q ;
  assign g9450 = \DFF_1504.Q ;
  assign g9453 = \DFF_58.Q ;
  assign g9465 = \DFF_1428.Q ;
  assign g9468 = \DFF_1427.Q ;
  assign g9471 = \DFF_42.Q ;
  assign g948 = \DFF_578.Q ;
  assign g9481 = \DFF_1429.Q ;
  assign g9484 = \DFF_1427.Q ;
  assign g9487 = \DFF_1083.Q ;
  assign g9488 = \DFF_86.Q ;
  assign g9498 = \DFF_1429.Q ;
  assign g9501 = \DFF_1428.Q ;
  assign g9504 = \DFF_107.Q ;
  assign g9505 = \DFF_110.Q ;
  assign g9506 = \DFF_112.Q ;
  assign g9507 = \DFF_80.Q ;
  assign g951 = \DFF_579.Q ;
  assign g9524 = \DFF_1429.Q ;
  assign g9528 = \DFF_1505.Q ;
  assign g9531 = \DFF_1504.Q ;
  assign g954 = \DFF_583.Q ;
  assign g9569 = \DFF_60.Q ;
  assign g957 = \DFF_584.Q ;
  assign g9585 = \DFF_1429.Q ;
  assign g9588 = \DFF_1428.Q ;
  assign g9591 = \DFF_734.Q ;
  assign g9592 = \DFF_1504.Q ;
  assign g9595 = \DFF_43.Q ;
  assign g960 = \DFF_585.Q ;
  assign g9607 = \DFF_1428.Q ;
  assign g9610 = \DFF_1427.Q ;
  assign g9613 = \DFF_87.Q ;
  assign g9623 = \DFF_1429.Q ;
  assign g9626 = \DFF_1427.Q ;
  assign g9629 = \DFF_1433.Q ;
  assign g963 = \DFF_1427.Q ;
  assign g9640 = \DFF_385.Q ;
  assign g9641 = \DFF_1506.Q ;
  assign g9644 = \DFF_1505.Q ;
  assign g9649 = \DFF_62.Q ;
  assign g966 = \DFF_653.Q ;
  assign g9666 = \DFF_1429.Q ;
  assign g967 = \DFF_654.Q ;
  assign g9670 = \DFF_1505.Q ;
  assign g9673 = \DFF_1504.Q ;
  assign g968 = \DFF_655.Q ;
  assign g969 = \DFF_656.Q ;
  assign g97 = \DFF_80.Q ;
  assign g970 = \DFF_657.Q ;
  assign g971 = \DFF_658.Q ;
  assign g9711 = \DFF_44.Q ;
  assign g972 = \DFF_659.Q ;
  assign g9727 = \DFF_1429.Q ;
  assign g973 = \DFF_660.Q ;
  assign g9730 = \DFF_1428.Q ;
  assign g9733 = \DFF_1084.Q ;
  assign g9734 = \DFF_1504.Q ;
  assign g9737 = \DFF_88.Q ;
  assign g974 = \DFF_661.Q ;
  assign g9749 = \DFF_1428.Q ;
  assign g975 = \DFF_662.Q ;
  assign g9752 = \DFF_1427.Q ;
  assign g9755 = \DFF_96.Q ;
  assign g9756 = \DFF_99.Q ;
  assign g9757 = \DFF_102.Q ;
  assign g9758 = \DFF_103.Q ;
  assign g976 = \DFF_663.Q ;
  assign g9767 = \DFF_1506.Q ;
  assign g977 = \DFF_664.Q ;
  assign g9770 = \DFF_1504.Q ;
  assign g978 = \DFF_665.Q ;
  assign g9786 = \DFF_735.Q ;
  assign g9787 = \DFF_1506.Q ;
  assign g9790 = \DFF_1505.Q ;
  assign g9795 = \DFF_45.Q ;
  assign g9812 = \DFF_1429.Q ;
  assign g9816 = \DFF_1505.Q ;
  assign g9819 = \DFF_1504.Q ;
  assign g985 = \DFF_678.Q ;
  assign g9857 = \DFF_89.Q ;
  assign g986 = \DFF_666.Q ;
  assign g9873 = \DFF_1429.Q ;
  assign g9876 = \DFF_1428.Q ;
  assign g9879 = \DFF_1434.Q ;
  assign g9880 = \DFF_1504.Q ;
  assign g9884 = \DFF_111.Q ;
  assign g9885 = \DFF_114.Q ;
  assign g9886 = \DFF_115.Q ;
  assign g9895 = \DFF_1505.Q ;
  assign g9898 = \DFF_1504.Q ;
  assign g9913 = \DFF_1506.Q ;
  assign g9916 = \DFF_1504.Q ;
  assign g992 = \DFF_667.Q ;
  assign g9932 = \DFF_1085.Q ;
  assign g9933 = \DFF_1506.Q ;
  assign g9936 = \DFF_1505.Q ;
  assign g9941 = \DFF_90.Q ;
  assign g9958 = \DFF_1429.Q ;
  assign g996 = \DFF_1302.Q ;
  assign g9962 = \DFF_1505.Q ;
  assign g9965 = \DFF_1504.Q ;
  assign g999 = \DFF_633.Q ;
endmodule
