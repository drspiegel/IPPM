
module s35932(GND, VDD, CK, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, CRC_OUT_1_30, CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_2, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29, CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, CRC_OUT_3_31, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_3, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, CRC_OUT_5_1, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19, CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_2, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29, CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, CRC_OUT_8_31, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_3, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_0_0, DATA_0_1, DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13, DATA_0_14, DATA_0_15, DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19, DATA_0_2, DATA_0_20, DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24, DATA_0_25, DATA_0_26, DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3, DATA_0_30, DATA_0_31, DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7, DATA_0_8, DATA_0_9, DATA_9_0, DATA_9_1, DATA_9_10, DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, DATA_9_15, DATA_9_16, DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, DATA_9_20, DATA_9_21, DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, DATA_9_26, DATA_9_27, DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, DATA_9_31, DATA_9_4, DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, RESET, TM0, TM1);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  input CK;
  output CRC_OUT_1_0;
  output CRC_OUT_1_1;
  output CRC_OUT_1_10;
  output CRC_OUT_1_11;
  output CRC_OUT_1_12;
  output CRC_OUT_1_13;
  output CRC_OUT_1_14;
  output CRC_OUT_1_15;
  output CRC_OUT_1_16;
  output CRC_OUT_1_17;
  output CRC_OUT_1_18;
  output CRC_OUT_1_19;
  output CRC_OUT_1_2;
  output CRC_OUT_1_20;
  output CRC_OUT_1_21;
  output CRC_OUT_1_22;
  output CRC_OUT_1_23;
  output CRC_OUT_1_24;
  output CRC_OUT_1_25;
  output CRC_OUT_1_26;
  output CRC_OUT_1_27;
  output CRC_OUT_1_28;
  output CRC_OUT_1_29;
  output CRC_OUT_1_3;
  output CRC_OUT_1_30;
  output CRC_OUT_1_31;
  output CRC_OUT_1_4;
  output CRC_OUT_1_5;
  output CRC_OUT_1_6;
  output CRC_OUT_1_7;
  output CRC_OUT_1_8;
  output CRC_OUT_1_9;
  output CRC_OUT_2_0;
  output CRC_OUT_2_1;
  output CRC_OUT_2_10;
  output CRC_OUT_2_11;
  output CRC_OUT_2_12;
  output CRC_OUT_2_13;
  output CRC_OUT_2_14;
  output CRC_OUT_2_15;
  output CRC_OUT_2_16;
  output CRC_OUT_2_17;
  output CRC_OUT_2_18;
  output CRC_OUT_2_19;
  output CRC_OUT_2_2;
  output CRC_OUT_2_20;
  output CRC_OUT_2_21;
  output CRC_OUT_2_22;
  output CRC_OUT_2_23;
  output CRC_OUT_2_24;
  output CRC_OUT_2_25;
  output CRC_OUT_2_26;
  output CRC_OUT_2_27;
  output CRC_OUT_2_28;
  output CRC_OUT_2_29;
  output CRC_OUT_2_3;
  output CRC_OUT_2_30;
  output CRC_OUT_2_31;
  output CRC_OUT_2_4;
  output CRC_OUT_2_5;
  output CRC_OUT_2_6;
  output CRC_OUT_2_7;
  output CRC_OUT_2_8;
  output CRC_OUT_2_9;
  output CRC_OUT_3_0;
  output CRC_OUT_3_1;
  output CRC_OUT_3_10;
  output CRC_OUT_3_11;
  output CRC_OUT_3_12;
  output CRC_OUT_3_13;
  output CRC_OUT_3_14;
  output CRC_OUT_3_15;
  output CRC_OUT_3_16;
  output CRC_OUT_3_17;
  output CRC_OUT_3_18;
  output CRC_OUT_3_19;
  output CRC_OUT_3_2;
  output CRC_OUT_3_20;
  output CRC_OUT_3_21;
  output CRC_OUT_3_22;
  output CRC_OUT_3_23;
  output CRC_OUT_3_24;
  output CRC_OUT_3_25;
  output CRC_OUT_3_26;
  output CRC_OUT_3_27;
  output CRC_OUT_3_28;
  output CRC_OUT_3_29;
  output CRC_OUT_3_3;
  output CRC_OUT_3_30;
  output CRC_OUT_3_31;
  output CRC_OUT_3_4;
  output CRC_OUT_3_5;
  output CRC_OUT_3_6;
  output CRC_OUT_3_7;
  output CRC_OUT_3_8;
  output CRC_OUT_3_9;
  output CRC_OUT_4_0;
  output CRC_OUT_4_1;
  output CRC_OUT_4_10;
  output CRC_OUT_4_11;
  output CRC_OUT_4_12;
  output CRC_OUT_4_13;
  output CRC_OUT_4_14;
  output CRC_OUT_4_15;
  output CRC_OUT_4_16;
  output CRC_OUT_4_17;
  output CRC_OUT_4_18;
  output CRC_OUT_4_19;
  output CRC_OUT_4_2;
  output CRC_OUT_4_20;
  output CRC_OUT_4_21;
  output CRC_OUT_4_22;
  output CRC_OUT_4_23;
  output CRC_OUT_4_24;
  output CRC_OUT_4_25;
  output CRC_OUT_4_26;
  output CRC_OUT_4_27;
  output CRC_OUT_4_28;
  output CRC_OUT_4_29;
  output CRC_OUT_4_3;
  output CRC_OUT_4_30;
  output CRC_OUT_4_31;
  output CRC_OUT_4_4;
  output CRC_OUT_4_5;
  output CRC_OUT_4_6;
  output CRC_OUT_4_7;
  output CRC_OUT_4_8;
  output CRC_OUT_4_9;
  output CRC_OUT_5_0;
  output CRC_OUT_5_1;
  output CRC_OUT_5_10;
  output CRC_OUT_5_11;
  output CRC_OUT_5_12;
  output CRC_OUT_5_13;
  output CRC_OUT_5_14;
  output CRC_OUT_5_15;
  output CRC_OUT_5_16;
  output CRC_OUT_5_17;
  output CRC_OUT_5_18;
  output CRC_OUT_5_19;
  output CRC_OUT_5_2;
  output CRC_OUT_5_20;
  output CRC_OUT_5_21;
  output CRC_OUT_5_22;
  output CRC_OUT_5_23;
  output CRC_OUT_5_24;
  output CRC_OUT_5_25;
  output CRC_OUT_5_26;
  output CRC_OUT_5_27;
  output CRC_OUT_5_28;
  output CRC_OUT_5_29;
  output CRC_OUT_5_3;
  output CRC_OUT_5_30;
  output CRC_OUT_5_31;
  output CRC_OUT_5_4;
  output CRC_OUT_5_5;
  output CRC_OUT_5_6;
  output CRC_OUT_5_7;
  output CRC_OUT_5_8;
  output CRC_OUT_5_9;
  output CRC_OUT_6_0;
  output CRC_OUT_6_1;
  output CRC_OUT_6_10;
  output CRC_OUT_6_11;
  output CRC_OUT_6_12;
  output CRC_OUT_6_13;
  output CRC_OUT_6_14;
  output CRC_OUT_6_15;
  output CRC_OUT_6_16;
  output CRC_OUT_6_17;
  output CRC_OUT_6_18;
  output CRC_OUT_6_19;
  output CRC_OUT_6_2;
  output CRC_OUT_6_20;
  output CRC_OUT_6_21;
  output CRC_OUT_6_22;
  output CRC_OUT_6_23;
  output CRC_OUT_6_24;
  output CRC_OUT_6_25;
  output CRC_OUT_6_26;
  output CRC_OUT_6_27;
  output CRC_OUT_6_28;
  output CRC_OUT_6_29;
  output CRC_OUT_6_3;
  output CRC_OUT_6_30;
  output CRC_OUT_6_31;
  output CRC_OUT_6_4;
  output CRC_OUT_6_5;
  output CRC_OUT_6_6;
  output CRC_OUT_6_7;
  output CRC_OUT_6_8;
  output CRC_OUT_6_9;
  output CRC_OUT_7_0;
  output CRC_OUT_7_1;
  output CRC_OUT_7_10;
  output CRC_OUT_7_11;
  output CRC_OUT_7_12;
  output CRC_OUT_7_13;
  output CRC_OUT_7_14;
  output CRC_OUT_7_15;
  output CRC_OUT_7_16;
  output CRC_OUT_7_17;
  output CRC_OUT_7_18;
  output CRC_OUT_7_19;
  output CRC_OUT_7_2;
  output CRC_OUT_7_20;
  output CRC_OUT_7_21;
  output CRC_OUT_7_22;
  output CRC_OUT_7_23;
  output CRC_OUT_7_24;
  output CRC_OUT_7_25;
  output CRC_OUT_7_26;
  output CRC_OUT_7_27;
  output CRC_OUT_7_28;
  output CRC_OUT_7_29;
  output CRC_OUT_7_3;
  output CRC_OUT_7_30;
  output CRC_OUT_7_31;
  output CRC_OUT_7_4;
  output CRC_OUT_7_5;
  output CRC_OUT_7_6;
  output CRC_OUT_7_7;
  output CRC_OUT_7_8;
  output CRC_OUT_7_9;
  output CRC_OUT_8_0;
  output CRC_OUT_8_1;
  output CRC_OUT_8_10;
  output CRC_OUT_8_11;
  output CRC_OUT_8_12;
  output CRC_OUT_8_13;
  output CRC_OUT_8_14;
  output CRC_OUT_8_15;
  output CRC_OUT_8_16;
  output CRC_OUT_8_17;
  output CRC_OUT_8_18;
  output CRC_OUT_8_19;
  output CRC_OUT_8_2;
  output CRC_OUT_8_20;
  output CRC_OUT_8_21;
  output CRC_OUT_8_22;
  output CRC_OUT_8_23;
  output CRC_OUT_8_24;
  output CRC_OUT_8_25;
  output CRC_OUT_8_26;
  output CRC_OUT_8_27;
  output CRC_OUT_8_28;
  output CRC_OUT_8_29;
  output CRC_OUT_8_3;
  output CRC_OUT_8_30;
  output CRC_OUT_8_31;
  output CRC_OUT_8_4;
  output CRC_OUT_8_5;
  output CRC_OUT_8_6;
  output CRC_OUT_8_7;
  output CRC_OUT_8_8;
  output CRC_OUT_8_9;
  output CRC_OUT_9_0;
  output CRC_OUT_9_1;
  output CRC_OUT_9_10;
  output CRC_OUT_9_11;
  output CRC_OUT_9_12;
  output CRC_OUT_9_13;
  output CRC_OUT_9_14;
  output CRC_OUT_9_15;
  output CRC_OUT_9_16;
  output CRC_OUT_9_17;
  output CRC_OUT_9_18;
  output CRC_OUT_9_19;
  output CRC_OUT_9_2;
  output CRC_OUT_9_20;
  output CRC_OUT_9_21;
  output CRC_OUT_9_22;
  output CRC_OUT_9_23;
  output CRC_OUT_9_24;
  output CRC_OUT_9_25;
  output CRC_OUT_9_26;
  output CRC_OUT_9_27;
  output CRC_OUT_9_28;
  output CRC_OUT_9_29;
  output CRC_OUT_9_3;
  output CRC_OUT_9_30;
  output CRC_OUT_9_31;
  output CRC_OUT_9_4;
  output CRC_OUT_9_5;
  output CRC_OUT_9_6;
  output CRC_OUT_9_7;
  output CRC_OUT_9_8;
  output CRC_OUT_9_9;
  input DATA_0_0;
  input DATA_0_1;
  input DATA_0_10;
  input DATA_0_11;
  input DATA_0_12;
  input DATA_0_13;
  input DATA_0_14;
  input DATA_0_15;
  input DATA_0_16;
  input DATA_0_17;
  input DATA_0_18;
  input DATA_0_19;
  input DATA_0_2;
  input DATA_0_20;
  input DATA_0_21;
  input DATA_0_22;
  input DATA_0_23;
  input DATA_0_24;
  input DATA_0_25;
  input DATA_0_26;
  input DATA_0_27;
  input DATA_0_28;
  input DATA_0_29;
  input DATA_0_3;
  input DATA_0_30;
  input DATA_0_31;
  input DATA_0_4;
  input DATA_0_5;
  input DATA_0_6;
  input DATA_0_7;
  input DATA_0_8;
  input DATA_0_9;
  output DATA_9_0;
  output DATA_9_1;
  output DATA_9_10;
  output DATA_9_11;
  output DATA_9_12;
  output DATA_9_13;
  output DATA_9_14;
  output DATA_9_15;
  output DATA_9_16;
  output DATA_9_17;
  output DATA_9_18;
  output DATA_9_19;
  output DATA_9_2;
  output DATA_9_20;
  output DATA_9_21;
  output DATA_9_22;
  output DATA_9_23;
  output DATA_9_24;
  output DATA_9_25;
  output DATA_9_26;
  output DATA_9_27;
  output DATA_9_28;
  output DATA_9_29;
  output DATA_9_3;
  output DATA_9_30;
  output DATA_9_31;
  output DATA_9_4;
  output DATA_9_5;
  output DATA_9_6;
  output DATA_9_7;
  output DATA_9_8;
  output DATA_9_9;
  wire \DFF_0.CK ;
  wire \DFF_0.D ;
  wire \DFF_0.Q ;
  wire \DFF_1.CK ;
  wire \DFF_1.D ;
  wire \DFF_1.Q ;
  wire \DFF_10.CK ;
  wire \DFF_10.D ;
  wire \DFF_10.Q ;
  wire \DFF_100.CK ;
  wire \DFF_100.D ;
  wire \DFF_100.Q ;
  wire \DFF_1000.CK ;
  wire \DFF_1000.D ;
  wire \DFF_1000.Q ;
  wire \DFF_1001.CK ;
  wire \DFF_1001.D ;
  wire \DFF_1001.Q ;
  wire \DFF_1002.CK ;
  wire \DFF_1002.D ;
  wire \DFF_1002.Q ;
  wire \DFF_1003.CK ;
  wire \DFF_1003.D ;
  wire \DFF_1003.Q ;
  wire \DFF_1004.CK ;
  wire \DFF_1004.D ;
  wire \DFF_1004.Q ;
  wire \DFF_1005.CK ;
  wire \DFF_1005.D ;
  wire \DFF_1005.Q ;
  wire \DFF_1006.CK ;
  wire \DFF_1006.D ;
  wire \DFF_1006.Q ;
  wire \DFF_1007.CK ;
  wire \DFF_1007.D ;
  wire \DFF_1007.Q ;
  wire \DFF_1008.CK ;
  wire \DFF_1008.D ;
  wire \DFF_1008.Q ;
  wire \DFF_1009.CK ;
  wire \DFF_1009.D ;
  wire \DFF_1009.Q ;
  wire \DFF_101.CK ;
  wire \DFF_101.D ;
  wire \DFF_101.Q ;
  wire \DFF_1010.CK ;
  wire \DFF_1010.D ;
  wire \DFF_1010.Q ;
  wire \DFF_1011.CK ;
  wire \DFF_1011.D ;
  wire \DFF_1011.Q ;
  wire \DFF_1012.CK ;
  wire \DFF_1012.D ;
  wire \DFF_1012.Q ;
  wire \DFF_1013.CK ;
  wire \DFF_1013.D ;
  wire \DFF_1013.Q ;
  wire \DFF_1014.CK ;
  wire \DFF_1014.D ;
  wire \DFF_1014.Q ;
  wire \DFF_1015.CK ;
  wire \DFF_1015.D ;
  wire \DFF_1015.Q ;
  wire \DFF_1016.CK ;
  wire \DFF_1016.D ;
  wire \DFF_1016.Q ;
  wire \DFF_1017.CK ;
  wire \DFF_1017.D ;
  wire \DFF_1017.Q ;
  wire \DFF_1018.CK ;
  wire \DFF_1018.D ;
  wire \DFF_1018.Q ;
  wire \DFF_1019.CK ;
  wire \DFF_1019.D ;
  wire \DFF_1019.Q ;
  wire \DFF_102.CK ;
  wire \DFF_102.D ;
  wire \DFF_102.Q ;
  wire \DFF_1020.CK ;
  wire \DFF_1020.D ;
  wire \DFF_1020.Q ;
  wire \DFF_1021.CK ;
  wire \DFF_1021.D ;
  wire \DFF_1021.Q ;
  wire \DFF_1022.CK ;
  wire \DFF_1022.D ;
  wire \DFF_1022.Q ;
  wire \DFF_1023.CK ;
  wire \DFF_1023.D ;
  wire \DFF_1023.Q ;
  wire \DFF_1024.CK ;
  wire \DFF_1024.D ;
  wire \DFF_1024.Q ;
  wire \DFF_1025.CK ;
  wire \DFF_1025.D ;
  wire \DFF_1025.Q ;
  wire \DFF_1026.CK ;
  wire \DFF_1026.D ;
  wire \DFF_1026.Q ;
  wire \DFF_1027.CK ;
  wire \DFF_1027.D ;
  wire \DFF_1027.Q ;
  wire \DFF_1028.CK ;
  wire \DFF_1028.D ;
  wire \DFF_1028.Q ;
  wire \DFF_1029.CK ;
  wire \DFF_1029.D ;
  wire \DFF_1029.Q ;
  wire \DFF_103.CK ;
  wire \DFF_103.D ;
  wire \DFF_103.Q ;
  wire \DFF_1030.CK ;
  wire \DFF_1030.D ;
  wire \DFF_1030.Q ;
  wire \DFF_1031.CK ;
  wire \DFF_1031.D ;
  wire \DFF_1031.Q ;
  wire \DFF_1032.CK ;
  wire \DFF_1032.D ;
  wire \DFF_1032.Q ;
  wire \DFF_1033.CK ;
  wire \DFF_1033.D ;
  wire \DFF_1033.Q ;
  wire \DFF_1034.CK ;
  wire \DFF_1034.D ;
  wire \DFF_1034.Q ;
  wire \DFF_1035.CK ;
  wire \DFF_1035.D ;
  wire \DFF_1035.Q ;
  wire \DFF_1036.CK ;
  wire \DFF_1036.D ;
  wire \DFF_1036.Q ;
  wire \DFF_1037.CK ;
  wire \DFF_1037.D ;
  wire \DFF_1037.Q ;
  wire \DFF_1038.CK ;
  wire \DFF_1038.D ;
  wire \DFF_1038.Q ;
  wire \DFF_1039.CK ;
  wire \DFF_1039.D ;
  wire \DFF_1039.Q ;
  wire \DFF_104.CK ;
  wire \DFF_104.D ;
  wire \DFF_104.Q ;
  wire \DFF_1040.CK ;
  wire \DFF_1040.D ;
  wire \DFF_1040.Q ;
  wire \DFF_1041.CK ;
  wire \DFF_1041.D ;
  wire \DFF_1041.Q ;
  wire \DFF_1042.CK ;
  wire \DFF_1042.D ;
  wire \DFF_1042.Q ;
  wire \DFF_1043.CK ;
  wire \DFF_1043.D ;
  wire \DFF_1043.Q ;
  wire \DFF_1044.CK ;
  wire \DFF_1044.D ;
  wire \DFF_1044.Q ;
  wire \DFF_1045.CK ;
  wire \DFF_1045.D ;
  wire \DFF_1045.Q ;
  wire \DFF_1046.CK ;
  wire \DFF_1046.D ;
  wire \DFF_1046.Q ;
  wire \DFF_1047.CK ;
  wire \DFF_1047.D ;
  wire \DFF_1047.Q ;
  wire \DFF_1048.CK ;
  wire \DFF_1048.D ;
  wire \DFF_1048.Q ;
  wire \DFF_1049.CK ;
  wire \DFF_1049.D ;
  wire \DFF_1049.Q ;
  wire \DFF_105.CK ;
  wire \DFF_105.D ;
  wire \DFF_105.Q ;
  wire \DFF_1050.CK ;
  wire \DFF_1050.D ;
  wire \DFF_1050.Q ;
  wire \DFF_1051.CK ;
  wire \DFF_1051.D ;
  wire \DFF_1051.Q ;
  wire \DFF_1052.CK ;
  wire \DFF_1052.D ;
  wire \DFF_1052.Q ;
  wire \DFF_1053.CK ;
  wire \DFF_1053.D ;
  wire \DFF_1053.Q ;
  wire \DFF_1054.CK ;
  wire \DFF_1054.D ;
  wire \DFF_1054.Q ;
  wire \DFF_1055.CK ;
  wire \DFF_1055.D ;
  wire \DFF_1055.Q ;
  wire \DFF_1056.CK ;
  wire \DFF_1056.D ;
  wire \DFF_1056.Q ;
  wire \DFF_1057.CK ;
  wire \DFF_1057.D ;
  wire \DFF_1057.Q ;
  wire \DFF_1058.CK ;
  wire \DFF_1058.D ;
  wire \DFF_1058.Q ;
  wire \DFF_1059.CK ;
  wire \DFF_1059.D ;
  wire \DFF_1059.Q ;
  wire \DFF_106.CK ;
  wire \DFF_106.D ;
  wire \DFF_106.Q ;
  wire \DFF_1060.CK ;
  wire \DFF_1060.D ;
  wire \DFF_1060.Q ;
  wire \DFF_1061.CK ;
  wire \DFF_1061.D ;
  wire \DFF_1061.Q ;
  wire \DFF_1062.CK ;
  wire \DFF_1062.D ;
  wire \DFF_1062.Q ;
  wire \DFF_1063.CK ;
  wire \DFF_1063.D ;
  wire \DFF_1063.Q ;
  wire \DFF_1064.CK ;
  wire \DFF_1064.D ;
  wire \DFF_1064.Q ;
  wire \DFF_1065.CK ;
  wire \DFF_1065.D ;
  wire \DFF_1065.Q ;
  wire \DFF_1066.CK ;
  wire \DFF_1066.D ;
  wire \DFF_1066.Q ;
  wire \DFF_1067.CK ;
  wire \DFF_1067.D ;
  wire \DFF_1067.Q ;
  wire \DFF_1068.CK ;
  wire \DFF_1068.D ;
  wire \DFF_1068.Q ;
  wire \DFF_1069.CK ;
  wire \DFF_1069.D ;
  wire \DFF_1069.Q ;
  wire \DFF_107.CK ;
  wire \DFF_107.D ;
  wire \DFF_107.Q ;
  wire \DFF_1070.CK ;
  wire \DFF_1070.D ;
  wire \DFF_1070.Q ;
  wire \DFF_1071.CK ;
  wire \DFF_1071.D ;
  wire \DFF_1071.Q ;
  wire \DFF_1072.CK ;
  wire \DFF_1072.D ;
  wire \DFF_1072.Q ;
  wire \DFF_1073.CK ;
  wire \DFF_1073.D ;
  wire \DFF_1073.Q ;
  wire \DFF_1074.CK ;
  wire \DFF_1074.D ;
  wire \DFF_1074.Q ;
  wire \DFF_1075.CK ;
  wire \DFF_1075.D ;
  wire \DFF_1075.Q ;
  wire \DFF_1076.CK ;
  wire \DFF_1076.D ;
  wire \DFF_1076.Q ;
  wire \DFF_1077.CK ;
  wire \DFF_1077.D ;
  wire \DFF_1077.Q ;
  wire \DFF_1078.CK ;
  wire \DFF_1078.D ;
  wire \DFF_1078.Q ;
  wire \DFF_1079.CK ;
  wire \DFF_1079.D ;
  wire \DFF_1079.Q ;
  wire \DFF_108.CK ;
  wire \DFF_108.D ;
  wire \DFF_108.Q ;
  wire \DFF_1080.CK ;
  wire \DFF_1080.D ;
  wire \DFF_1080.Q ;
  wire \DFF_1081.CK ;
  wire \DFF_1081.D ;
  wire \DFF_1081.Q ;
  wire \DFF_1082.CK ;
  wire \DFF_1082.D ;
  wire \DFF_1082.Q ;
  wire \DFF_1083.CK ;
  wire \DFF_1083.D ;
  wire \DFF_1083.Q ;
  wire \DFF_1084.CK ;
  wire \DFF_1084.D ;
  wire \DFF_1084.Q ;
  wire \DFF_1085.CK ;
  wire \DFF_1085.D ;
  wire \DFF_1085.Q ;
  wire \DFF_1086.CK ;
  wire \DFF_1086.D ;
  wire \DFF_1086.Q ;
  wire \DFF_1087.CK ;
  wire \DFF_1087.D ;
  wire \DFF_1087.Q ;
  wire \DFF_1088.CK ;
  wire \DFF_1088.D ;
  wire \DFF_1088.Q ;
  wire \DFF_1089.CK ;
  wire \DFF_1089.D ;
  wire \DFF_1089.Q ;
  wire \DFF_109.CK ;
  wire \DFF_109.D ;
  wire \DFF_109.Q ;
  wire \DFF_1090.CK ;
  wire \DFF_1090.D ;
  wire \DFF_1090.Q ;
  wire \DFF_1091.CK ;
  wire \DFF_1091.D ;
  wire \DFF_1091.Q ;
  wire \DFF_1092.CK ;
  wire \DFF_1092.D ;
  wire \DFF_1092.Q ;
  wire \DFF_1093.CK ;
  wire \DFF_1093.D ;
  wire \DFF_1093.Q ;
  wire \DFF_1094.CK ;
  wire \DFF_1094.D ;
  wire \DFF_1094.Q ;
  wire \DFF_1095.CK ;
  wire \DFF_1095.D ;
  wire \DFF_1095.Q ;
  wire \DFF_1096.CK ;
  wire \DFF_1096.D ;
  wire \DFF_1096.Q ;
  wire \DFF_1097.CK ;
  wire \DFF_1097.D ;
  wire \DFF_1097.Q ;
  wire \DFF_1098.CK ;
  wire \DFF_1098.D ;
  wire \DFF_1098.Q ;
  wire \DFF_1099.CK ;
  wire \DFF_1099.D ;
  wire \DFF_1099.Q ;
  wire \DFF_11.CK ;
  wire \DFF_11.D ;
  wire \DFF_11.Q ;
  wire \DFF_110.CK ;
  wire \DFF_110.D ;
  wire \DFF_110.Q ;
  wire \DFF_1100.CK ;
  wire \DFF_1100.D ;
  wire \DFF_1100.Q ;
  wire \DFF_1101.CK ;
  wire \DFF_1101.D ;
  wire \DFF_1101.Q ;
  wire \DFF_1102.CK ;
  wire \DFF_1102.D ;
  wire \DFF_1102.Q ;
  wire \DFF_1103.CK ;
  wire \DFF_1103.D ;
  wire \DFF_1103.Q ;
  wire \DFF_1104.CK ;
  wire \DFF_1104.D ;
  wire \DFF_1104.Q ;
  wire \DFF_1105.CK ;
  wire \DFF_1105.D ;
  wire \DFF_1105.Q ;
  wire \DFF_1106.CK ;
  wire \DFF_1106.D ;
  wire \DFF_1106.Q ;
  wire \DFF_1107.CK ;
  wire \DFF_1107.D ;
  wire \DFF_1107.Q ;
  wire \DFF_1108.CK ;
  wire \DFF_1108.D ;
  wire \DFF_1108.Q ;
  wire \DFF_1109.CK ;
  wire \DFF_1109.D ;
  wire \DFF_1109.Q ;
  wire \DFF_111.CK ;
  wire \DFF_111.D ;
  wire \DFF_111.Q ;
  wire \DFF_1110.CK ;
  wire \DFF_1110.D ;
  wire \DFF_1110.Q ;
  wire \DFF_1111.CK ;
  wire \DFF_1111.D ;
  wire \DFF_1111.Q ;
  wire \DFF_1112.CK ;
  wire \DFF_1112.D ;
  wire \DFF_1112.Q ;
  wire \DFF_1113.CK ;
  wire \DFF_1113.D ;
  wire \DFF_1113.Q ;
  wire \DFF_1114.CK ;
  wire \DFF_1114.D ;
  wire \DFF_1114.Q ;
  wire \DFF_1115.CK ;
  wire \DFF_1115.D ;
  wire \DFF_1115.Q ;
  wire \DFF_1116.CK ;
  wire \DFF_1116.D ;
  wire \DFF_1116.Q ;
  wire \DFF_1117.CK ;
  wire \DFF_1117.D ;
  wire \DFF_1117.Q ;
  wire \DFF_1118.CK ;
  wire \DFF_1118.D ;
  wire \DFF_1118.Q ;
  wire \DFF_1119.CK ;
  wire \DFF_1119.D ;
  wire \DFF_1119.Q ;
  wire \DFF_112.CK ;
  wire \DFF_112.D ;
  wire \DFF_112.Q ;
  wire \DFF_1120.CK ;
  wire \DFF_1120.D ;
  wire \DFF_1120.Q ;
  wire \DFF_1121.CK ;
  wire \DFF_1121.D ;
  wire \DFF_1121.Q ;
  wire \DFF_1122.CK ;
  wire \DFF_1122.D ;
  wire \DFF_1122.Q ;
  wire \DFF_1123.CK ;
  wire \DFF_1123.D ;
  wire \DFF_1123.Q ;
  wire \DFF_1124.CK ;
  wire \DFF_1124.D ;
  wire \DFF_1124.Q ;
  wire \DFF_1125.CK ;
  wire \DFF_1125.D ;
  wire \DFF_1125.Q ;
  wire \DFF_1126.CK ;
  wire \DFF_1126.D ;
  wire \DFF_1126.Q ;
  wire \DFF_1127.CK ;
  wire \DFF_1127.D ;
  wire \DFF_1127.Q ;
  wire \DFF_1128.CK ;
  wire \DFF_1128.D ;
  wire \DFF_1128.Q ;
  wire \DFF_1129.CK ;
  wire \DFF_1129.D ;
  wire \DFF_1129.Q ;
  wire \DFF_113.CK ;
  wire \DFF_113.D ;
  wire \DFF_113.Q ;
  wire \DFF_1130.CK ;
  wire \DFF_1130.D ;
  wire \DFF_1130.Q ;
  wire \DFF_1131.CK ;
  wire \DFF_1131.D ;
  wire \DFF_1131.Q ;
  wire \DFF_1132.CK ;
  wire \DFF_1132.D ;
  wire \DFF_1132.Q ;
  wire \DFF_1133.CK ;
  wire \DFF_1133.D ;
  wire \DFF_1133.Q ;
  wire \DFF_1134.CK ;
  wire \DFF_1134.D ;
  wire \DFF_1134.Q ;
  wire \DFF_1135.CK ;
  wire \DFF_1135.D ;
  wire \DFF_1135.Q ;
  wire \DFF_1136.CK ;
  wire \DFF_1136.D ;
  wire \DFF_1136.Q ;
  wire \DFF_1137.CK ;
  wire \DFF_1137.D ;
  wire \DFF_1137.Q ;
  wire \DFF_1138.CK ;
  wire \DFF_1138.D ;
  wire \DFF_1138.Q ;
  wire \DFF_1139.CK ;
  wire \DFF_1139.D ;
  wire \DFF_1139.Q ;
  wire \DFF_114.CK ;
  wire \DFF_114.D ;
  wire \DFF_114.Q ;
  wire \DFF_1140.CK ;
  wire \DFF_1140.D ;
  wire \DFF_1140.Q ;
  wire \DFF_1141.CK ;
  wire \DFF_1141.D ;
  wire \DFF_1141.Q ;
  wire \DFF_1142.CK ;
  wire \DFF_1142.D ;
  wire \DFF_1142.Q ;
  wire \DFF_1143.CK ;
  wire \DFF_1143.D ;
  wire \DFF_1143.Q ;
  wire \DFF_1144.CK ;
  wire \DFF_1144.D ;
  wire \DFF_1144.Q ;
  wire \DFF_1145.CK ;
  wire \DFF_1145.D ;
  wire \DFF_1145.Q ;
  wire \DFF_1146.CK ;
  wire \DFF_1146.D ;
  wire \DFF_1146.Q ;
  wire \DFF_1147.CK ;
  wire \DFF_1147.D ;
  wire \DFF_1147.Q ;
  wire \DFF_1148.CK ;
  wire \DFF_1148.D ;
  wire \DFF_1148.Q ;
  wire \DFF_1149.CK ;
  wire \DFF_1149.D ;
  wire \DFF_1149.Q ;
  wire \DFF_115.CK ;
  wire \DFF_115.D ;
  wire \DFF_115.Q ;
  wire \DFF_1150.CK ;
  wire \DFF_1150.D ;
  wire \DFF_1150.Q ;
  wire \DFF_1151.CK ;
  wire \DFF_1151.D ;
  wire \DFF_1151.Q ;
  wire \DFF_1152.CK ;
  wire \DFF_1152.D ;
  wire \DFF_1152.Q ;
  wire \DFF_1153.CK ;
  wire \DFF_1153.D ;
  wire \DFF_1153.Q ;
  wire \DFF_1154.CK ;
  wire \DFF_1154.D ;
  wire \DFF_1154.Q ;
  wire \DFF_1155.CK ;
  wire \DFF_1155.D ;
  wire \DFF_1155.Q ;
  wire \DFF_1156.CK ;
  wire \DFF_1156.D ;
  wire \DFF_1156.Q ;
  wire \DFF_1157.CK ;
  wire \DFF_1157.D ;
  wire \DFF_1157.Q ;
  wire \DFF_1158.CK ;
  wire \DFF_1158.D ;
  wire \DFF_1158.Q ;
  wire \DFF_1159.CK ;
  wire \DFF_1159.D ;
  wire \DFF_1159.Q ;
  wire \DFF_116.CK ;
  wire \DFF_116.D ;
  wire \DFF_116.Q ;
  wire \DFF_1160.CK ;
  wire \DFF_1160.D ;
  wire \DFF_1160.Q ;
  wire \DFF_1161.CK ;
  wire \DFF_1161.D ;
  wire \DFF_1161.Q ;
  wire \DFF_1162.CK ;
  wire \DFF_1162.D ;
  wire \DFF_1162.Q ;
  wire \DFF_1163.CK ;
  wire \DFF_1163.D ;
  wire \DFF_1163.Q ;
  wire \DFF_1164.CK ;
  wire \DFF_1164.D ;
  wire \DFF_1164.Q ;
  wire \DFF_1165.CK ;
  wire \DFF_1165.D ;
  wire \DFF_1165.Q ;
  wire \DFF_1166.CK ;
  wire \DFF_1166.D ;
  wire \DFF_1166.Q ;
  wire \DFF_1167.CK ;
  wire \DFF_1167.D ;
  wire \DFF_1167.Q ;
  wire \DFF_1168.CK ;
  wire \DFF_1168.D ;
  wire \DFF_1168.Q ;
  wire \DFF_1169.CK ;
  wire \DFF_1169.D ;
  wire \DFF_1169.Q ;
  wire \DFF_117.CK ;
  wire \DFF_117.D ;
  wire \DFF_117.Q ;
  wire \DFF_1170.CK ;
  wire \DFF_1170.D ;
  wire \DFF_1170.Q ;
  wire \DFF_1171.CK ;
  wire \DFF_1171.D ;
  wire \DFF_1171.Q ;
  wire \DFF_1172.CK ;
  wire \DFF_1172.D ;
  wire \DFF_1172.Q ;
  wire \DFF_1173.CK ;
  wire \DFF_1173.D ;
  wire \DFF_1173.Q ;
  wire \DFF_1174.CK ;
  wire \DFF_1174.D ;
  wire \DFF_1174.Q ;
  wire \DFF_1175.CK ;
  wire \DFF_1175.D ;
  wire \DFF_1175.Q ;
  wire \DFF_1176.CK ;
  wire \DFF_1176.D ;
  wire \DFF_1176.Q ;
  wire \DFF_1177.CK ;
  wire \DFF_1177.D ;
  wire \DFF_1177.Q ;
  wire \DFF_1178.CK ;
  wire \DFF_1178.D ;
  wire \DFF_1178.Q ;
  wire \DFF_1179.CK ;
  wire \DFF_1179.D ;
  wire \DFF_1179.Q ;
  wire \DFF_118.CK ;
  wire \DFF_118.D ;
  wire \DFF_118.Q ;
  wire \DFF_1180.CK ;
  wire \DFF_1180.D ;
  wire \DFF_1180.Q ;
  wire \DFF_1181.CK ;
  wire \DFF_1181.D ;
  wire \DFF_1181.Q ;
  wire \DFF_1182.CK ;
  wire \DFF_1182.D ;
  wire \DFF_1182.Q ;
  wire \DFF_1183.CK ;
  wire \DFF_1183.D ;
  wire \DFF_1183.Q ;
  wire \DFF_1184.CK ;
  wire \DFF_1184.D ;
  wire \DFF_1184.Q ;
  wire \DFF_1185.CK ;
  wire \DFF_1185.D ;
  wire \DFF_1185.Q ;
  wire \DFF_1186.CK ;
  wire \DFF_1186.D ;
  wire \DFF_1186.Q ;
  wire \DFF_1187.CK ;
  wire \DFF_1187.D ;
  wire \DFF_1187.Q ;
  wire \DFF_1188.CK ;
  wire \DFF_1188.D ;
  wire \DFF_1188.Q ;
  wire \DFF_1189.CK ;
  wire \DFF_1189.D ;
  wire \DFF_1189.Q ;
  wire \DFF_119.CK ;
  wire \DFF_119.D ;
  wire \DFF_119.Q ;
  wire \DFF_1190.CK ;
  wire \DFF_1190.D ;
  wire \DFF_1190.Q ;
  wire \DFF_1191.CK ;
  wire \DFF_1191.D ;
  wire \DFF_1191.Q ;
  wire \DFF_1192.CK ;
  wire \DFF_1192.D ;
  wire \DFF_1192.Q ;
  wire \DFF_1193.CK ;
  wire \DFF_1193.D ;
  wire \DFF_1193.Q ;
  wire \DFF_1194.CK ;
  wire \DFF_1194.D ;
  wire \DFF_1194.Q ;
  wire \DFF_1195.CK ;
  wire \DFF_1195.D ;
  wire \DFF_1195.Q ;
  wire \DFF_1196.CK ;
  wire \DFF_1196.D ;
  wire \DFF_1196.Q ;
  wire \DFF_1197.CK ;
  wire \DFF_1197.D ;
  wire \DFF_1197.Q ;
  wire \DFF_1198.CK ;
  wire \DFF_1198.D ;
  wire \DFF_1198.Q ;
  wire \DFF_1199.CK ;
  wire \DFF_1199.D ;
  wire \DFF_1199.Q ;
  wire \DFF_12.CK ;
  wire \DFF_12.D ;
  wire \DFF_12.Q ;
  wire \DFF_120.CK ;
  wire \DFF_120.D ;
  wire \DFF_120.Q ;
  wire \DFF_1200.CK ;
  wire \DFF_1200.D ;
  wire \DFF_1200.Q ;
  wire \DFF_1201.CK ;
  wire \DFF_1201.D ;
  wire \DFF_1201.Q ;
  wire \DFF_1202.CK ;
  wire \DFF_1202.D ;
  wire \DFF_1202.Q ;
  wire \DFF_1203.CK ;
  wire \DFF_1203.D ;
  wire \DFF_1203.Q ;
  wire \DFF_1204.CK ;
  wire \DFF_1204.D ;
  wire \DFF_1204.Q ;
  wire \DFF_1205.CK ;
  wire \DFF_1205.D ;
  wire \DFF_1205.Q ;
  wire \DFF_1206.CK ;
  wire \DFF_1206.D ;
  wire \DFF_1206.Q ;
  wire \DFF_1207.CK ;
  wire \DFF_1207.D ;
  wire \DFF_1207.Q ;
  wire \DFF_1208.CK ;
  wire \DFF_1208.D ;
  wire \DFF_1208.Q ;
  wire \DFF_1209.CK ;
  wire \DFF_1209.D ;
  wire \DFF_1209.Q ;
  wire \DFF_121.CK ;
  wire \DFF_121.D ;
  wire \DFF_121.Q ;
  wire \DFF_1210.CK ;
  wire \DFF_1210.D ;
  wire \DFF_1210.Q ;
  wire \DFF_1211.CK ;
  wire \DFF_1211.D ;
  wire \DFF_1211.Q ;
  wire \DFF_1212.CK ;
  wire \DFF_1212.D ;
  wire \DFF_1212.Q ;
  wire \DFF_1213.CK ;
  wire \DFF_1213.D ;
  wire \DFF_1213.Q ;
  wire \DFF_1214.CK ;
  wire \DFF_1214.D ;
  wire \DFF_1214.Q ;
  wire \DFF_1215.CK ;
  wire \DFF_1215.D ;
  wire \DFF_1215.Q ;
  wire \DFF_1216.CK ;
  wire \DFF_1216.D ;
  wire \DFF_1216.Q ;
  wire \DFF_1217.CK ;
  wire \DFF_1217.D ;
  wire \DFF_1217.Q ;
  wire \DFF_1218.CK ;
  wire \DFF_1218.D ;
  wire \DFF_1218.Q ;
  wire \DFF_1219.CK ;
  wire \DFF_1219.D ;
  wire \DFF_1219.Q ;
  wire \DFF_122.CK ;
  wire \DFF_122.D ;
  wire \DFF_122.Q ;
  wire \DFF_1220.CK ;
  wire \DFF_1220.D ;
  wire \DFF_1220.Q ;
  wire \DFF_1221.CK ;
  wire \DFF_1221.D ;
  wire \DFF_1221.Q ;
  wire \DFF_1222.CK ;
  wire \DFF_1222.D ;
  wire \DFF_1222.Q ;
  wire \DFF_1223.CK ;
  wire \DFF_1223.D ;
  wire \DFF_1223.Q ;
  wire \DFF_1224.CK ;
  wire \DFF_1224.D ;
  wire \DFF_1224.Q ;
  wire \DFF_1225.CK ;
  wire \DFF_1225.D ;
  wire \DFF_1225.Q ;
  wire \DFF_1226.CK ;
  wire \DFF_1226.D ;
  wire \DFF_1226.Q ;
  wire \DFF_1227.CK ;
  wire \DFF_1227.D ;
  wire \DFF_1227.Q ;
  wire \DFF_1228.CK ;
  wire \DFF_1228.D ;
  wire \DFF_1228.Q ;
  wire \DFF_1229.CK ;
  wire \DFF_1229.D ;
  wire \DFF_1229.Q ;
  wire \DFF_123.CK ;
  wire \DFF_123.D ;
  wire \DFF_123.Q ;
  wire \DFF_1230.CK ;
  wire \DFF_1230.D ;
  wire \DFF_1230.Q ;
  wire \DFF_1231.CK ;
  wire \DFF_1231.D ;
  wire \DFF_1231.Q ;
  wire \DFF_1232.CK ;
  wire \DFF_1232.D ;
  wire \DFF_1232.Q ;
  wire \DFF_1233.CK ;
  wire \DFF_1233.D ;
  wire \DFF_1233.Q ;
  wire \DFF_1234.CK ;
  wire \DFF_1234.D ;
  wire \DFF_1234.Q ;
  wire \DFF_1235.CK ;
  wire \DFF_1235.D ;
  wire \DFF_1235.Q ;
  wire \DFF_1236.CK ;
  wire \DFF_1236.D ;
  wire \DFF_1236.Q ;
  wire \DFF_1237.CK ;
  wire \DFF_1237.D ;
  wire \DFF_1237.Q ;
  wire \DFF_1238.CK ;
  wire \DFF_1238.D ;
  wire \DFF_1238.Q ;
  wire \DFF_1239.CK ;
  wire \DFF_1239.D ;
  wire \DFF_1239.Q ;
  wire \DFF_124.CK ;
  wire \DFF_124.D ;
  wire \DFF_124.Q ;
  wire \DFF_1240.CK ;
  wire \DFF_1240.D ;
  wire \DFF_1240.Q ;
  wire \DFF_1241.CK ;
  wire \DFF_1241.D ;
  wire \DFF_1241.Q ;
  wire \DFF_1242.CK ;
  wire \DFF_1242.D ;
  wire \DFF_1242.Q ;
  wire \DFF_1243.CK ;
  wire \DFF_1243.D ;
  wire \DFF_1243.Q ;
  wire \DFF_1244.CK ;
  wire \DFF_1244.D ;
  wire \DFF_1244.Q ;
  wire \DFF_1245.CK ;
  wire \DFF_1245.D ;
  wire \DFF_1245.Q ;
  wire \DFF_1246.CK ;
  wire \DFF_1246.D ;
  wire \DFF_1246.Q ;
  wire \DFF_1247.CK ;
  wire \DFF_1247.D ;
  wire \DFF_1247.Q ;
  wire \DFF_1248.CK ;
  wire \DFF_1248.D ;
  wire \DFF_1248.Q ;
  wire \DFF_1249.CK ;
  wire \DFF_1249.D ;
  wire \DFF_1249.Q ;
  wire \DFF_125.CK ;
  wire \DFF_125.D ;
  wire \DFF_125.Q ;
  wire \DFF_1250.CK ;
  wire \DFF_1250.D ;
  wire \DFF_1250.Q ;
  wire \DFF_1251.CK ;
  wire \DFF_1251.D ;
  wire \DFF_1251.Q ;
  wire \DFF_1252.CK ;
  wire \DFF_1252.D ;
  wire \DFF_1252.Q ;
  wire \DFF_1253.CK ;
  wire \DFF_1253.D ;
  wire \DFF_1253.Q ;
  wire \DFF_1254.CK ;
  wire \DFF_1254.D ;
  wire \DFF_1254.Q ;
  wire \DFF_1255.CK ;
  wire \DFF_1255.D ;
  wire \DFF_1255.Q ;
  wire \DFF_1256.CK ;
  wire \DFF_1256.D ;
  wire \DFF_1256.Q ;
  wire \DFF_1257.CK ;
  wire \DFF_1257.D ;
  wire \DFF_1257.Q ;
  wire \DFF_1258.CK ;
  wire \DFF_1258.D ;
  wire \DFF_1258.Q ;
  wire \DFF_1259.CK ;
  wire \DFF_1259.D ;
  wire \DFF_1259.Q ;
  wire \DFF_126.CK ;
  wire \DFF_126.D ;
  wire \DFF_126.Q ;
  wire \DFF_1260.CK ;
  wire \DFF_1260.D ;
  wire \DFF_1260.Q ;
  wire \DFF_1261.CK ;
  wire \DFF_1261.D ;
  wire \DFF_1261.Q ;
  wire \DFF_1262.CK ;
  wire \DFF_1262.D ;
  wire \DFF_1262.Q ;
  wire \DFF_1263.CK ;
  wire \DFF_1263.D ;
  wire \DFF_1263.Q ;
  wire \DFF_1264.CK ;
  wire \DFF_1264.D ;
  wire \DFF_1264.Q ;
  wire \DFF_1265.CK ;
  wire \DFF_1265.D ;
  wire \DFF_1265.Q ;
  wire \DFF_1266.CK ;
  wire \DFF_1266.D ;
  wire \DFF_1266.Q ;
  wire \DFF_1267.CK ;
  wire \DFF_1267.D ;
  wire \DFF_1267.Q ;
  wire \DFF_1268.CK ;
  wire \DFF_1268.D ;
  wire \DFF_1268.Q ;
  wire \DFF_1269.CK ;
  wire \DFF_1269.D ;
  wire \DFF_1269.Q ;
  wire \DFF_127.CK ;
  wire \DFF_127.D ;
  wire \DFF_127.Q ;
  wire \DFF_1270.CK ;
  wire \DFF_1270.D ;
  wire \DFF_1270.Q ;
  wire \DFF_1271.CK ;
  wire \DFF_1271.D ;
  wire \DFF_1271.Q ;
  wire \DFF_1272.CK ;
  wire \DFF_1272.D ;
  wire \DFF_1272.Q ;
  wire \DFF_1273.CK ;
  wire \DFF_1273.D ;
  wire \DFF_1273.Q ;
  wire \DFF_1274.CK ;
  wire \DFF_1274.D ;
  wire \DFF_1274.Q ;
  wire \DFF_1275.CK ;
  wire \DFF_1275.D ;
  wire \DFF_1275.Q ;
  wire \DFF_1276.CK ;
  wire \DFF_1276.D ;
  wire \DFF_1276.Q ;
  wire \DFF_1277.CK ;
  wire \DFF_1277.D ;
  wire \DFF_1277.Q ;
  wire \DFF_1278.CK ;
  wire \DFF_1278.D ;
  wire \DFF_1278.Q ;
  wire \DFF_1279.CK ;
  wire \DFF_1279.D ;
  wire \DFF_1279.Q ;
  wire \DFF_128.CK ;
  wire \DFF_128.D ;
  wire \DFF_128.Q ;
  wire \DFF_1280.CK ;
  wire \DFF_1280.D ;
  wire \DFF_1280.Q ;
  wire \DFF_1281.CK ;
  wire \DFF_1281.D ;
  wire \DFF_1281.Q ;
  wire \DFF_1282.CK ;
  wire \DFF_1282.D ;
  wire \DFF_1282.Q ;
  wire \DFF_1283.CK ;
  wire \DFF_1283.D ;
  wire \DFF_1283.Q ;
  wire \DFF_1284.CK ;
  wire \DFF_1284.D ;
  wire \DFF_1284.Q ;
  wire \DFF_1285.CK ;
  wire \DFF_1285.D ;
  wire \DFF_1285.Q ;
  wire \DFF_1286.CK ;
  wire \DFF_1286.D ;
  wire \DFF_1286.Q ;
  wire \DFF_1287.CK ;
  wire \DFF_1287.D ;
  wire \DFF_1287.Q ;
  wire \DFF_1288.CK ;
  wire \DFF_1288.D ;
  wire \DFF_1288.Q ;
  wire \DFF_1289.CK ;
  wire \DFF_1289.D ;
  wire \DFF_1289.Q ;
  wire \DFF_129.CK ;
  wire \DFF_129.D ;
  wire \DFF_129.Q ;
  wire \DFF_1290.CK ;
  wire \DFF_1290.D ;
  wire \DFF_1290.Q ;
  wire \DFF_1291.CK ;
  wire \DFF_1291.D ;
  wire \DFF_1291.Q ;
  wire \DFF_1292.CK ;
  wire \DFF_1292.D ;
  wire \DFF_1292.Q ;
  wire \DFF_1293.CK ;
  wire \DFF_1293.D ;
  wire \DFF_1293.Q ;
  wire \DFF_1294.CK ;
  wire \DFF_1294.D ;
  wire \DFF_1294.Q ;
  wire \DFF_1295.CK ;
  wire \DFF_1295.D ;
  wire \DFF_1295.Q ;
  wire \DFF_1296.CK ;
  wire \DFF_1296.D ;
  wire \DFF_1296.Q ;
  wire \DFF_1297.CK ;
  wire \DFF_1297.D ;
  wire \DFF_1297.Q ;
  wire \DFF_1298.CK ;
  wire \DFF_1298.D ;
  wire \DFF_1298.Q ;
  wire \DFF_1299.CK ;
  wire \DFF_1299.D ;
  wire \DFF_1299.Q ;
  wire \DFF_13.CK ;
  wire \DFF_13.D ;
  wire \DFF_13.Q ;
  wire \DFF_130.CK ;
  wire \DFF_130.D ;
  wire \DFF_130.Q ;
  wire \DFF_1300.CK ;
  wire \DFF_1300.D ;
  wire \DFF_1300.Q ;
  wire \DFF_1301.CK ;
  wire \DFF_1301.D ;
  wire \DFF_1301.Q ;
  wire \DFF_1302.CK ;
  wire \DFF_1302.D ;
  wire \DFF_1302.Q ;
  wire \DFF_1303.CK ;
  wire \DFF_1303.D ;
  wire \DFF_1303.Q ;
  wire \DFF_1304.CK ;
  wire \DFF_1304.D ;
  wire \DFF_1304.Q ;
  wire \DFF_1305.CK ;
  wire \DFF_1305.D ;
  wire \DFF_1305.Q ;
  wire \DFF_1306.CK ;
  wire \DFF_1306.D ;
  wire \DFF_1306.Q ;
  wire \DFF_1307.CK ;
  wire \DFF_1307.D ;
  wire \DFF_1307.Q ;
  wire \DFF_1308.CK ;
  wire \DFF_1308.D ;
  wire \DFF_1308.Q ;
  wire \DFF_1309.CK ;
  wire \DFF_1309.D ;
  wire \DFF_1309.Q ;
  wire \DFF_131.CK ;
  wire \DFF_131.D ;
  wire \DFF_131.Q ;
  wire \DFF_1310.CK ;
  wire \DFF_1310.D ;
  wire \DFF_1310.Q ;
  wire \DFF_1311.CK ;
  wire \DFF_1311.D ;
  wire \DFF_1311.Q ;
  wire \DFF_1312.CK ;
  wire \DFF_1312.D ;
  wire \DFF_1312.Q ;
  wire \DFF_1313.CK ;
  wire \DFF_1313.D ;
  wire \DFF_1313.Q ;
  wire \DFF_1314.CK ;
  wire \DFF_1314.D ;
  wire \DFF_1314.Q ;
  wire \DFF_1315.CK ;
  wire \DFF_1315.D ;
  wire \DFF_1315.Q ;
  wire \DFF_1316.CK ;
  wire \DFF_1316.D ;
  wire \DFF_1316.Q ;
  wire \DFF_1317.CK ;
  wire \DFF_1317.D ;
  wire \DFF_1317.Q ;
  wire \DFF_1318.CK ;
  wire \DFF_1318.D ;
  wire \DFF_1318.Q ;
  wire \DFF_1319.CK ;
  wire \DFF_1319.D ;
  wire \DFF_1319.Q ;
  wire \DFF_132.CK ;
  wire \DFF_132.D ;
  wire \DFF_132.Q ;
  wire \DFF_1320.CK ;
  wire \DFF_1320.D ;
  wire \DFF_1320.Q ;
  wire \DFF_1321.CK ;
  wire \DFF_1321.D ;
  wire \DFF_1321.Q ;
  wire \DFF_1322.CK ;
  wire \DFF_1322.D ;
  wire \DFF_1322.Q ;
  wire \DFF_1323.CK ;
  wire \DFF_1323.D ;
  wire \DFF_1323.Q ;
  wire \DFF_1324.CK ;
  wire \DFF_1324.D ;
  wire \DFF_1324.Q ;
  wire \DFF_1325.CK ;
  wire \DFF_1325.D ;
  wire \DFF_1325.Q ;
  wire \DFF_1326.CK ;
  wire \DFF_1326.D ;
  wire \DFF_1326.Q ;
  wire \DFF_1327.CK ;
  wire \DFF_1327.D ;
  wire \DFF_1327.Q ;
  wire \DFF_1328.CK ;
  wire \DFF_1328.D ;
  wire \DFF_1328.Q ;
  wire \DFF_1329.CK ;
  wire \DFF_1329.D ;
  wire \DFF_1329.Q ;
  wire \DFF_133.CK ;
  wire \DFF_133.D ;
  wire \DFF_133.Q ;
  wire \DFF_1330.CK ;
  wire \DFF_1330.D ;
  wire \DFF_1330.Q ;
  wire \DFF_1331.CK ;
  wire \DFF_1331.D ;
  wire \DFF_1331.Q ;
  wire \DFF_1332.CK ;
  wire \DFF_1332.D ;
  wire \DFF_1332.Q ;
  wire \DFF_1333.CK ;
  wire \DFF_1333.D ;
  wire \DFF_1333.Q ;
  wire \DFF_1334.CK ;
  wire \DFF_1334.D ;
  wire \DFF_1334.Q ;
  wire \DFF_1335.CK ;
  wire \DFF_1335.D ;
  wire \DFF_1335.Q ;
  wire \DFF_1336.CK ;
  wire \DFF_1336.D ;
  wire \DFF_1336.Q ;
  wire \DFF_1337.CK ;
  wire \DFF_1337.D ;
  wire \DFF_1337.Q ;
  wire \DFF_1338.CK ;
  wire \DFF_1338.D ;
  wire \DFF_1338.Q ;
  wire \DFF_1339.CK ;
  wire \DFF_1339.D ;
  wire \DFF_1339.Q ;
  wire \DFF_134.CK ;
  wire \DFF_134.D ;
  wire \DFF_134.Q ;
  wire \DFF_1340.CK ;
  wire \DFF_1340.D ;
  wire \DFF_1340.Q ;
  wire \DFF_1341.CK ;
  wire \DFF_1341.D ;
  wire \DFF_1341.Q ;
  wire \DFF_1342.CK ;
  wire \DFF_1342.D ;
  wire \DFF_1342.Q ;
  wire \DFF_1343.CK ;
  wire \DFF_1343.D ;
  wire \DFF_1343.Q ;
  wire \DFF_1344.CK ;
  wire \DFF_1344.D ;
  wire \DFF_1344.Q ;
  wire \DFF_1345.CK ;
  wire \DFF_1345.D ;
  wire \DFF_1345.Q ;
  wire \DFF_1346.CK ;
  wire \DFF_1346.D ;
  wire \DFF_1346.Q ;
  wire \DFF_1347.CK ;
  wire \DFF_1347.D ;
  wire \DFF_1347.Q ;
  wire \DFF_1348.CK ;
  wire \DFF_1348.D ;
  wire \DFF_1348.Q ;
  wire \DFF_1349.CK ;
  wire \DFF_1349.D ;
  wire \DFF_1349.Q ;
  wire \DFF_135.CK ;
  wire \DFF_135.D ;
  wire \DFF_135.Q ;
  wire \DFF_1350.CK ;
  wire \DFF_1350.D ;
  wire \DFF_1350.Q ;
  wire \DFF_1351.CK ;
  wire \DFF_1351.D ;
  wire \DFF_1351.Q ;
  wire \DFF_1352.CK ;
  wire \DFF_1352.D ;
  wire \DFF_1352.Q ;
  wire \DFF_1353.CK ;
  wire \DFF_1353.D ;
  wire \DFF_1353.Q ;
  wire \DFF_1354.CK ;
  wire \DFF_1354.D ;
  wire \DFF_1354.Q ;
  wire \DFF_1355.CK ;
  wire \DFF_1355.D ;
  wire \DFF_1355.Q ;
  wire \DFF_1356.CK ;
  wire \DFF_1356.D ;
  wire \DFF_1356.Q ;
  wire \DFF_1357.CK ;
  wire \DFF_1357.D ;
  wire \DFF_1357.Q ;
  wire \DFF_1358.CK ;
  wire \DFF_1358.D ;
  wire \DFF_1358.Q ;
  wire \DFF_1359.CK ;
  wire \DFF_1359.D ;
  wire \DFF_1359.Q ;
  wire \DFF_136.CK ;
  wire \DFF_136.D ;
  wire \DFF_136.Q ;
  wire \DFF_1360.CK ;
  wire \DFF_1360.D ;
  wire \DFF_1360.Q ;
  wire \DFF_1361.CK ;
  wire \DFF_1361.D ;
  wire \DFF_1361.Q ;
  wire \DFF_1362.CK ;
  wire \DFF_1362.D ;
  wire \DFF_1362.Q ;
  wire \DFF_1363.CK ;
  wire \DFF_1363.D ;
  wire \DFF_1363.Q ;
  wire \DFF_1364.CK ;
  wire \DFF_1364.D ;
  wire \DFF_1364.Q ;
  wire \DFF_1365.CK ;
  wire \DFF_1365.D ;
  wire \DFF_1365.Q ;
  wire \DFF_1366.CK ;
  wire \DFF_1366.D ;
  wire \DFF_1366.Q ;
  wire \DFF_1367.CK ;
  wire \DFF_1367.D ;
  wire \DFF_1367.Q ;
  wire \DFF_1368.CK ;
  wire \DFF_1368.D ;
  wire \DFF_1368.Q ;
  wire \DFF_1369.CK ;
  wire \DFF_1369.D ;
  wire \DFF_1369.Q ;
  wire \DFF_137.CK ;
  wire \DFF_137.D ;
  wire \DFF_137.Q ;
  wire \DFF_1370.CK ;
  wire \DFF_1370.D ;
  wire \DFF_1370.Q ;
  wire \DFF_1371.CK ;
  wire \DFF_1371.D ;
  wire \DFF_1371.Q ;
  wire \DFF_1372.CK ;
  wire \DFF_1372.D ;
  wire \DFF_1372.Q ;
  wire \DFF_1373.CK ;
  wire \DFF_1373.D ;
  wire \DFF_1373.Q ;
  wire \DFF_1374.CK ;
  wire \DFF_1374.D ;
  wire \DFF_1374.Q ;
  wire \DFF_1375.CK ;
  wire \DFF_1375.D ;
  wire \DFF_1375.Q ;
  wire \DFF_1376.CK ;
  wire \DFF_1376.D ;
  wire \DFF_1376.Q ;
  wire \DFF_1377.CK ;
  wire \DFF_1377.D ;
  wire \DFF_1377.Q ;
  wire \DFF_1378.CK ;
  wire \DFF_1378.D ;
  wire \DFF_1378.Q ;
  wire \DFF_1379.CK ;
  wire \DFF_1379.D ;
  wire \DFF_1379.Q ;
  wire \DFF_138.CK ;
  wire \DFF_138.D ;
  wire \DFF_138.Q ;
  wire \DFF_1380.CK ;
  wire \DFF_1380.D ;
  wire \DFF_1380.Q ;
  wire \DFF_1381.CK ;
  wire \DFF_1381.D ;
  wire \DFF_1381.Q ;
  wire \DFF_1382.CK ;
  wire \DFF_1382.D ;
  wire \DFF_1382.Q ;
  wire \DFF_1383.CK ;
  wire \DFF_1383.D ;
  wire \DFF_1383.Q ;
  wire \DFF_1384.CK ;
  wire \DFF_1384.D ;
  wire \DFF_1384.Q ;
  wire \DFF_1385.CK ;
  wire \DFF_1385.D ;
  wire \DFF_1385.Q ;
  wire \DFF_1386.CK ;
  wire \DFF_1386.D ;
  wire \DFF_1386.Q ;
  wire \DFF_1387.CK ;
  wire \DFF_1387.D ;
  wire \DFF_1387.Q ;
  wire \DFF_1388.CK ;
  wire \DFF_1388.D ;
  wire \DFF_1388.Q ;
  wire \DFF_1389.CK ;
  wire \DFF_1389.D ;
  wire \DFF_1389.Q ;
  wire \DFF_139.CK ;
  wire \DFF_139.D ;
  wire \DFF_139.Q ;
  wire \DFF_1390.CK ;
  wire \DFF_1390.D ;
  wire \DFF_1390.Q ;
  wire \DFF_1391.CK ;
  wire \DFF_1391.D ;
  wire \DFF_1391.Q ;
  wire \DFF_1392.CK ;
  wire \DFF_1392.D ;
  wire \DFF_1392.Q ;
  wire \DFF_1393.CK ;
  wire \DFF_1393.D ;
  wire \DFF_1393.Q ;
  wire \DFF_1394.CK ;
  wire \DFF_1394.D ;
  wire \DFF_1394.Q ;
  wire \DFF_1395.CK ;
  wire \DFF_1395.D ;
  wire \DFF_1395.Q ;
  wire \DFF_1396.CK ;
  wire \DFF_1396.D ;
  wire \DFF_1396.Q ;
  wire \DFF_1397.CK ;
  wire \DFF_1397.D ;
  wire \DFF_1397.Q ;
  wire \DFF_1398.CK ;
  wire \DFF_1398.D ;
  wire \DFF_1398.Q ;
  wire \DFF_1399.CK ;
  wire \DFF_1399.D ;
  wire \DFF_1399.Q ;
  wire \DFF_14.CK ;
  wire \DFF_14.D ;
  wire \DFF_14.Q ;
  wire \DFF_140.CK ;
  wire \DFF_140.D ;
  wire \DFF_140.Q ;
  wire \DFF_1400.CK ;
  wire \DFF_1400.D ;
  wire \DFF_1400.Q ;
  wire \DFF_1401.CK ;
  wire \DFF_1401.D ;
  wire \DFF_1401.Q ;
  wire \DFF_1402.CK ;
  wire \DFF_1402.D ;
  wire \DFF_1402.Q ;
  wire \DFF_1403.CK ;
  wire \DFF_1403.D ;
  wire \DFF_1403.Q ;
  wire \DFF_1404.CK ;
  wire \DFF_1404.D ;
  wire \DFF_1404.Q ;
  wire \DFF_1405.CK ;
  wire \DFF_1405.D ;
  wire \DFF_1405.Q ;
  wire \DFF_1406.CK ;
  wire \DFF_1406.D ;
  wire \DFF_1406.Q ;
  wire \DFF_1407.CK ;
  wire \DFF_1407.D ;
  wire \DFF_1407.Q ;
  wire \DFF_1408.CK ;
  wire \DFF_1408.D ;
  wire \DFF_1408.Q ;
  wire \DFF_1409.CK ;
  wire \DFF_1409.D ;
  wire \DFF_1409.Q ;
  wire \DFF_141.CK ;
  wire \DFF_141.D ;
  wire \DFF_141.Q ;
  wire \DFF_1410.CK ;
  wire \DFF_1410.D ;
  wire \DFF_1410.Q ;
  wire \DFF_1411.CK ;
  wire \DFF_1411.D ;
  wire \DFF_1411.Q ;
  wire \DFF_1412.CK ;
  wire \DFF_1412.D ;
  wire \DFF_1412.Q ;
  wire \DFF_1413.CK ;
  wire \DFF_1413.D ;
  wire \DFF_1413.Q ;
  wire \DFF_1414.CK ;
  wire \DFF_1414.D ;
  wire \DFF_1414.Q ;
  wire \DFF_1415.CK ;
  wire \DFF_1415.D ;
  wire \DFF_1415.Q ;
  wire \DFF_1416.CK ;
  wire \DFF_1416.D ;
  wire \DFF_1416.Q ;
  wire \DFF_1417.CK ;
  wire \DFF_1417.D ;
  wire \DFF_1417.Q ;
  wire \DFF_1418.CK ;
  wire \DFF_1418.D ;
  wire \DFF_1418.Q ;
  wire \DFF_1419.CK ;
  wire \DFF_1419.D ;
  wire \DFF_1419.Q ;
  wire \DFF_142.CK ;
  wire \DFF_142.D ;
  wire \DFF_142.Q ;
  wire \DFF_1420.CK ;
  wire \DFF_1420.D ;
  wire \DFF_1420.Q ;
  wire \DFF_1421.CK ;
  wire \DFF_1421.D ;
  wire \DFF_1421.Q ;
  wire \DFF_1422.CK ;
  wire \DFF_1422.D ;
  wire \DFF_1422.Q ;
  wire \DFF_1423.CK ;
  wire \DFF_1423.D ;
  wire \DFF_1423.Q ;
  wire \DFF_1424.CK ;
  wire \DFF_1424.D ;
  wire \DFF_1424.Q ;
  wire \DFF_1425.CK ;
  wire \DFF_1425.D ;
  wire \DFF_1425.Q ;
  wire \DFF_1426.CK ;
  wire \DFF_1426.D ;
  wire \DFF_1426.Q ;
  wire \DFF_1427.CK ;
  wire \DFF_1427.D ;
  wire \DFF_1427.Q ;
  wire \DFF_1428.CK ;
  wire \DFF_1428.D ;
  wire \DFF_1428.Q ;
  wire \DFF_1429.CK ;
  wire \DFF_1429.D ;
  wire \DFF_1429.Q ;
  wire \DFF_143.CK ;
  wire \DFF_143.D ;
  wire \DFF_143.Q ;
  wire \DFF_1430.CK ;
  wire \DFF_1430.D ;
  wire \DFF_1430.Q ;
  wire \DFF_1431.CK ;
  wire \DFF_1431.D ;
  wire \DFF_1431.Q ;
  wire \DFF_1432.CK ;
  wire \DFF_1432.D ;
  wire \DFF_1432.Q ;
  wire \DFF_1433.CK ;
  wire \DFF_1433.D ;
  wire \DFF_1433.Q ;
  wire \DFF_1434.CK ;
  wire \DFF_1434.D ;
  wire \DFF_1434.Q ;
  wire \DFF_1435.CK ;
  wire \DFF_1435.D ;
  wire \DFF_1435.Q ;
  wire \DFF_1436.CK ;
  wire \DFF_1436.D ;
  wire \DFF_1436.Q ;
  wire \DFF_1437.CK ;
  wire \DFF_1437.D ;
  wire \DFF_1437.Q ;
  wire \DFF_1438.CK ;
  wire \DFF_1438.D ;
  wire \DFF_1438.Q ;
  wire \DFF_1439.CK ;
  wire \DFF_1439.D ;
  wire \DFF_1439.Q ;
  wire \DFF_144.CK ;
  wire \DFF_144.D ;
  wire \DFF_144.Q ;
  wire \DFF_1440.CK ;
  wire \DFF_1440.D ;
  wire \DFF_1440.Q ;
  wire \DFF_1441.CK ;
  wire \DFF_1441.D ;
  wire \DFF_1441.Q ;
  wire \DFF_1442.CK ;
  wire \DFF_1442.D ;
  wire \DFF_1442.Q ;
  wire \DFF_1443.CK ;
  wire \DFF_1443.D ;
  wire \DFF_1443.Q ;
  wire \DFF_1444.CK ;
  wire \DFF_1444.D ;
  wire \DFF_1444.Q ;
  wire \DFF_1445.CK ;
  wire \DFF_1445.D ;
  wire \DFF_1445.Q ;
  wire \DFF_1446.CK ;
  wire \DFF_1446.D ;
  wire \DFF_1446.Q ;
  wire \DFF_1447.CK ;
  wire \DFF_1447.D ;
  wire \DFF_1447.Q ;
  wire \DFF_1448.CK ;
  wire \DFF_1448.D ;
  wire \DFF_1448.Q ;
  wire \DFF_1449.CK ;
  wire \DFF_1449.D ;
  wire \DFF_1449.Q ;
  wire \DFF_145.CK ;
  wire \DFF_145.D ;
  wire \DFF_145.Q ;
  wire \DFF_1450.CK ;
  wire \DFF_1450.D ;
  wire \DFF_1450.Q ;
  wire \DFF_1451.CK ;
  wire \DFF_1451.D ;
  wire \DFF_1451.Q ;
  wire \DFF_1452.CK ;
  wire \DFF_1452.D ;
  wire \DFF_1452.Q ;
  wire \DFF_1453.CK ;
  wire \DFF_1453.D ;
  wire \DFF_1453.Q ;
  wire \DFF_1454.CK ;
  wire \DFF_1454.D ;
  wire \DFF_1454.Q ;
  wire \DFF_1455.CK ;
  wire \DFF_1455.D ;
  wire \DFF_1455.Q ;
  wire \DFF_1456.CK ;
  wire \DFF_1456.D ;
  wire \DFF_1456.Q ;
  wire \DFF_1457.CK ;
  wire \DFF_1457.D ;
  wire \DFF_1457.Q ;
  wire \DFF_1458.CK ;
  wire \DFF_1458.D ;
  wire \DFF_1458.Q ;
  wire \DFF_1459.CK ;
  wire \DFF_1459.D ;
  wire \DFF_1459.Q ;
  wire \DFF_146.CK ;
  wire \DFF_146.D ;
  wire \DFF_146.Q ;
  wire \DFF_1460.CK ;
  wire \DFF_1460.D ;
  wire \DFF_1460.Q ;
  wire \DFF_1461.CK ;
  wire \DFF_1461.D ;
  wire \DFF_1461.Q ;
  wire \DFF_1462.CK ;
  wire \DFF_1462.D ;
  wire \DFF_1462.Q ;
  wire \DFF_1463.CK ;
  wire \DFF_1463.D ;
  wire \DFF_1463.Q ;
  wire \DFF_1464.CK ;
  wire \DFF_1464.D ;
  wire \DFF_1464.Q ;
  wire \DFF_1465.CK ;
  wire \DFF_1465.D ;
  wire \DFF_1465.Q ;
  wire \DFF_1466.CK ;
  wire \DFF_1466.D ;
  wire \DFF_1466.Q ;
  wire \DFF_1467.CK ;
  wire \DFF_1467.D ;
  wire \DFF_1467.Q ;
  wire \DFF_1468.CK ;
  wire \DFF_1468.D ;
  wire \DFF_1468.Q ;
  wire \DFF_1469.CK ;
  wire \DFF_1469.D ;
  wire \DFF_1469.Q ;
  wire \DFF_147.CK ;
  wire \DFF_147.D ;
  wire \DFF_147.Q ;
  wire \DFF_1470.CK ;
  wire \DFF_1470.D ;
  wire \DFF_1470.Q ;
  wire \DFF_1471.CK ;
  wire \DFF_1471.D ;
  wire \DFF_1471.Q ;
  wire \DFF_1472.CK ;
  wire \DFF_1472.D ;
  wire \DFF_1472.Q ;
  wire \DFF_1473.CK ;
  wire \DFF_1473.D ;
  wire \DFF_1473.Q ;
  wire \DFF_1474.CK ;
  wire \DFF_1474.D ;
  wire \DFF_1474.Q ;
  wire \DFF_1475.CK ;
  wire \DFF_1475.D ;
  wire \DFF_1475.Q ;
  wire \DFF_1476.CK ;
  wire \DFF_1476.D ;
  wire \DFF_1476.Q ;
  wire \DFF_1477.CK ;
  wire \DFF_1477.D ;
  wire \DFF_1477.Q ;
  wire \DFF_1478.CK ;
  wire \DFF_1478.D ;
  wire \DFF_1478.Q ;
  wire \DFF_1479.CK ;
  wire \DFF_1479.D ;
  wire \DFF_1479.Q ;
  wire \DFF_148.CK ;
  wire \DFF_148.D ;
  wire \DFF_148.Q ;
  wire \DFF_1480.CK ;
  wire \DFF_1480.D ;
  wire \DFF_1480.Q ;
  wire \DFF_1481.CK ;
  wire \DFF_1481.D ;
  wire \DFF_1481.Q ;
  wire \DFF_1482.CK ;
  wire \DFF_1482.D ;
  wire \DFF_1482.Q ;
  wire \DFF_1483.CK ;
  wire \DFF_1483.D ;
  wire \DFF_1483.Q ;
  wire \DFF_1484.CK ;
  wire \DFF_1484.D ;
  wire \DFF_1484.Q ;
  wire \DFF_1485.CK ;
  wire \DFF_1485.D ;
  wire \DFF_1485.Q ;
  wire \DFF_1486.CK ;
  wire \DFF_1486.D ;
  wire \DFF_1486.Q ;
  wire \DFF_1487.CK ;
  wire \DFF_1487.D ;
  wire \DFF_1487.Q ;
  wire \DFF_1488.CK ;
  wire \DFF_1488.D ;
  wire \DFF_1488.Q ;
  wire \DFF_1489.CK ;
  wire \DFF_1489.D ;
  wire \DFF_1489.Q ;
  wire \DFF_149.CK ;
  wire \DFF_149.D ;
  wire \DFF_149.Q ;
  wire \DFF_1490.CK ;
  wire \DFF_1490.D ;
  wire \DFF_1490.Q ;
  wire \DFF_1491.CK ;
  wire \DFF_1491.D ;
  wire \DFF_1491.Q ;
  wire \DFF_1492.CK ;
  wire \DFF_1492.D ;
  wire \DFF_1492.Q ;
  wire \DFF_1493.CK ;
  wire \DFF_1493.D ;
  wire \DFF_1493.Q ;
  wire \DFF_1494.CK ;
  wire \DFF_1494.D ;
  wire \DFF_1494.Q ;
  wire \DFF_1495.CK ;
  wire \DFF_1495.D ;
  wire \DFF_1495.Q ;
  wire \DFF_1496.CK ;
  wire \DFF_1496.D ;
  wire \DFF_1496.Q ;
  wire \DFF_1497.CK ;
  wire \DFF_1497.D ;
  wire \DFF_1497.Q ;
  wire \DFF_1498.CK ;
  wire \DFF_1498.D ;
  wire \DFF_1498.Q ;
  wire \DFF_1499.CK ;
  wire \DFF_1499.D ;
  wire \DFF_1499.Q ;
  wire \DFF_15.CK ;
  wire \DFF_15.D ;
  wire \DFF_15.Q ;
  wire \DFF_150.CK ;
  wire \DFF_150.D ;
  wire \DFF_150.Q ;
  wire \DFF_1500.CK ;
  wire \DFF_1500.D ;
  wire \DFF_1500.Q ;
  wire \DFF_1501.CK ;
  wire \DFF_1501.D ;
  wire \DFF_1501.Q ;
  wire \DFF_1502.CK ;
  wire \DFF_1502.D ;
  wire \DFF_1502.Q ;
  wire \DFF_1503.CK ;
  wire \DFF_1503.D ;
  wire \DFF_1503.Q ;
  wire \DFF_1504.CK ;
  wire \DFF_1504.D ;
  wire \DFF_1504.Q ;
  wire \DFF_1505.CK ;
  wire \DFF_1505.D ;
  wire \DFF_1505.Q ;
  wire \DFF_1506.CK ;
  wire \DFF_1506.D ;
  wire \DFF_1506.Q ;
  wire \DFF_1507.CK ;
  wire \DFF_1507.D ;
  wire \DFF_1507.Q ;
  wire \DFF_1508.CK ;
  wire \DFF_1508.D ;
  wire \DFF_1508.Q ;
  wire \DFF_1509.CK ;
  wire \DFF_1509.D ;
  wire \DFF_1509.Q ;
  wire \DFF_151.CK ;
  wire \DFF_151.D ;
  wire \DFF_151.Q ;
  wire \DFF_1510.CK ;
  wire \DFF_1510.D ;
  wire \DFF_1510.Q ;
  wire \DFF_1511.CK ;
  wire \DFF_1511.D ;
  wire \DFF_1511.Q ;
  wire \DFF_1512.CK ;
  wire \DFF_1512.D ;
  wire \DFF_1512.Q ;
  wire \DFF_1513.CK ;
  wire \DFF_1513.D ;
  wire \DFF_1513.Q ;
  wire \DFF_1514.CK ;
  wire \DFF_1514.D ;
  wire \DFF_1514.Q ;
  wire \DFF_1515.CK ;
  wire \DFF_1515.D ;
  wire \DFF_1515.Q ;
  wire \DFF_1516.CK ;
  wire \DFF_1516.D ;
  wire \DFF_1516.Q ;
  wire \DFF_1517.CK ;
  wire \DFF_1517.D ;
  wire \DFF_1517.Q ;
  wire \DFF_1518.CK ;
  wire \DFF_1518.D ;
  wire \DFF_1518.Q ;
  wire \DFF_1519.CK ;
  wire \DFF_1519.D ;
  wire \DFF_1519.Q ;
  wire \DFF_152.CK ;
  wire \DFF_152.D ;
  wire \DFF_152.Q ;
  wire \DFF_1520.CK ;
  wire \DFF_1520.D ;
  wire \DFF_1520.Q ;
  wire \DFF_1521.CK ;
  wire \DFF_1521.D ;
  wire \DFF_1521.Q ;
  wire \DFF_1522.CK ;
  wire \DFF_1522.D ;
  wire \DFF_1522.Q ;
  wire \DFF_1523.CK ;
  wire \DFF_1523.D ;
  wire \DFF_1523.Q ;
  wire \DFF_1524.CK ;
  wire \DFF_1524.D ;
  wire \DFF_1524.Q ;
  wire \DFF_1525.CK ;
  wire \DFF_1525.D ;
  wire \DFF_1525.Q ;
  wire \DFF_1526.CK ;
  wire \DFF_1526.D ;
  wire \DFF_1526.Q ;
  wire \DFF_1527.CK ;
  wire \DFF_1527.D ;
  wire \DFF_1527.Q ;
  wire \DFF_1528.CK ;
  wire \DFF_1528.D ;
  wire \DFF_1528.Q ;
  wire \DFF_1529.CK ;
  wire \DFF_1529.D ;
  wire \DFF_1529.Q ;
  wire \DFF_153.CK ;
  wire \DFF_153.D ;
  wire \DFF_153.Q ;
  wire \DFF_1530.CK ;
  wire \DFF_1530.D ;
  wire \DFF_1530.Q ;
  wire \DFF_1531.CK ;
  wire \DFF_1531.D ;
  wire \DFF_1531.Q ;
  wire \DFF_1532.CK ;
  wire \DFF_1532.D ;
  wire \DFF_1532.Q ;
  wire \DFF_1533.CK ;
  wire \DFF_1533.D ;
  wire \DFF_1533.Q ;
  wire \DFF_1534.CK ;
  wire \DFF_1534.D ;
  wire \DFF_1534.Q ;
  wire \DFF_1535.CK ;
  wire \DFF_1535.D ;
  wire \DFF_1535.Q ;
  wire \DFF_1536.CK ;
  wire \DFF_1536.D ;
  wire \DFF_1536.Q ;
  wire \DFF_1537.CK ;
  wire \DFF_1537.D ;
  wire \DFF_1537.Q ;
  wire \DFF_1538.CK ;
  wire \DFF_1538.D ;
  wire \DFF_1538.Q ;
  wire \DFF_1539.CK ;
  wire \DFF_1539.D ;
  wire \DFF_1539.Q ;
  wire \DFF_154.CK ;
  wire \DFF_154.D ;
  wire \DFF_154.Q ;
  wire \DFF_1540.CK ;
  wire \DFF_1540.D ;
  wire \DFF_1540.Q ;
  wire \DFF_1541.CK ;
  wire \DFF_1541.D ;
  wire \DFF_1541.Q ;
  wire \DFF_1542.CK ;
  wire \DFF_1542.D ;
  wire \DFF_1542.Q ;
  wire \DFF_1543.CK ;
  wire \DFF_1543.D ;
  wire \DFF_1543.Q ;
  wire \DFF_1544.CK ;
  wire \DFF_1544.D ;
  wire \DFF_1544.Q ;
  wire \DFF_1545.CK ;
  wire \DFF_1545.D ;
  wire \DFF_1545.Q ;
  wire \DFF_1546.CK ;
  wire \DFF_1546.D ;
  wire \DFF_1546.Q ;
  wire \DFF_1547.CK ;
  wire \DFF_1547.D ;
  wire \DFF_1547.Q ;
  wire \DFF_1548.CK ;
  wire \DFF_1548.D ;
  wire \DFF_1548.Q ;
  wire \DFF_1549.CK ;
  wire \DFF_1549.D ;
  wire \DFF_1549.Q ;
  wire \DFF_155.CK ;
  wire \DFF_155.D ;
  wire \DFF_155.Q ;
  wire \DFF_1550.CK ;
  wire \DFF_1550.D ;
  wire \DFF_1550.Q ;
  wire \DFF_1551.CK ;
  wire \DFF_1551.D ;
  wire \DFF_1551.Q ;
  wire \DFF_1552.CK ;
  wire \DFF_1552.D ;
  wire \DFF_1552.Q ;
  wire \DFF_1553.CK ;
  wire \DFF_1553.D ;
  wire \DFF_1553.Q ;
  wire \DFF_1554.CK ;
  wire \DFF_1554.D ;
  wire \DFF_1554.Q ;
  wire \DFF_1555.CK ;
  wire \DFF_1555.D ;
  wire \DFF_1555.Q ;
  wire \DFF_1556.CK ;
  wire \DFF_1556.D ;
  wire \DFF_1556.Q ;
  wire \DFF_1557.CK ;
  wire \DFF_1557.D ;
  wire \DFF_1557.Q ;
  wire \DFF_1558.CK ;
  wire \DFF_1558.D ;
  wire \DFF_1558.Q ;
  wire \DFF_1559.CK ;
  wire \DFF_1559.D ;
  wire \DFF_1559.Q ;
  wire \DFF_156.CK ;
  wire \DFF_156.D ;
  wire \DFF_156.Q ;
  wire \DFF_1560.CK ;
  wire \DFF_1560.D ;
  wire \DFF_1560.Q ;
  wire \DFF_1561.CK ;
  wire \DFF_1561.D ;
  wire \DFF_1561.Q ;
  wire \DFF_1562.CK ;
  wire \DFF_1562.D ;
  wire \DFF_1562.Q ;
  wire \DFF_1563.CK ;
  wire \DFF_1563.D ;
  wire \DFF_1563.Q ;
  wire \DFF_1564.CK ;
  wire \DFF_1564.D ;
  wire \DFF_1564.Q ;
  wire \DFF_1565.CK ;
  wire \DFF_1565.D ;
  wire \DFF_1565.Q ;
  wire \DFF_1566.CK ;
  wire \DFF_1566.D ;
  wire \DFF_1566.Q ;
  wire \DFF_1567.CK ;
  wire \DFF_1567.D ;
  wire \DFF_1567.Q ;
  wire \DFF_1568.CK ;
  wire \DFF_1568.D ;
  wire \DFF_1568.Q ;
  wire \DFF_1569.CK ;
  wire \DFF_1569.D ;
  wire \DFF_1569.Q ;
  wire \DFF_157.CK ;
  wire \DFF_157.D ;
  wire \DFF_157.Q ;
  wire \DFF_1570.CK ;
  wire \DFF_1570.D ;
  wire \DFF_1570.Q ;
  wire \DFF_1571.CK ;
  wire \DFF_1571.D ;
  wire \DFF_1571.Q ;
  wire \DFF_1572.CK ;
  wire \DFF_1572.D ;
  wire \DFF_1572.Q ;
  wire \DFF_1573.CK ;
  wire \DFF_1573.D ;
  wire \DFF_1573.Q ;
  wire \DFF_1574.CK ;
  wire \DFF_1574.D ;
  wire \DFF_1574.Q ;
  wire \DFF_1575.CK ;
  wire \DFF_1575.D ;
  wire \DFF_1575.Q ;
  wire \DFF_1576.CK ;
  wire \DFF_1576.D ;
  wire \DFF_1576.Q ;
  wire \DFF_1577.CK ;
  wire \DFF_1577.D ;
  wire \DFF_1577.Q ;
  wire \DFF_1578.CK ;
  wire \DFF_1578.D ;
  wire \DFF_1578.Q ;
  wire \DFF_1579.CK ;
  wire \DFF_1579.D ;
  wire \DFF_1579.Q ;
  wire \DFF_158.CK ;
  wire \DFF_158.D ;
  wire \DFF_158.Q ;
  wire \DFF_1580.CK ;
  wire \DFF_1580.D ;
  wire \DFF_1580.Q ;
  wire \DFF_1581.CK ;
  wire \DFF_1581.D ;
  wire \DFF_1581.Q ;
  wire \DFF_1582.CK ;
  wire \DFF_1582.D ;
  wire \DFF_1582.Q ;
  wire \DFF_1583.CK ;
  wire \DFF_1583.D ;
  wire \DFF_1583.Q ;
  wire \DFF_1584.CK ;
  wire \DFF_1584.D ;
  wire \DFF_1584.Q ;
  wire \DFF_1585.CK ;
  wire \DFF_1585.D ;
  wire \DFF_1585.Q ;
  wire \DFF_1586.CK ;
  wire \DFF_1586.D ;
  wire \DFF_1586.Q ;
  wire \DFF_1587.CK ;
  wire \DFF_1587.D ;
  wire \DFF_1587.Q ;
  wire \DFF_1588.CK ;
  wire \DFF_1588.D ;
  wire \DFF_1588.Q ;
  wire \DFF_1589.CK ;
  wire \DFF_1589.D ;
  wire \DFF_1589.Q ;
  wire \DFF_159.CK ;
  wire \DFF_159.D ;
  wire \DFF_159.Q ;
  wire \DFF_1590.CK ;
  wire \DFF_1590.D ;
  wire \DFF_1590.Q ;
  wire \DFF_1591.CK ;
  wire \DFF_1591.D ;
  wire \DFF_1591.Q ;
  wire \DFF_1592.CK ;
  wire \DFF_1592.D ;
  wire \DFF_1592.Q ;
  wire \DFF_1593.CK ;
  wire \DFF_1593.D ;
  wire \DFF_1593.Q ;
  wire \DFF_1594.CK ;
  wire \DFF_1594.D ;
  wire \DFF_1594.Q ;
  wire \DFF_1595.CK ;
  wire \DFF_1595.D ;
  wire \DFF_1595.Q ;
  wire \DFF_1596.CK ;
  wire \DFF_1596.D ;
  wire \DFF_1596.Q ;
  wire \DFF_1597.CK ;
  wire \DFF_1597.D ;
  wire \DFF_1597.Q ;
  wire \DFF_1598.CK ;
  wire \DFF_1598.D ;
  wire \DFF_1598.Q ;
  wire \DFF_1599.CK ;
  wire \DFF_1599.D ;
  wire \DFF_1599.Q ;
  wire \DFF_16.CK ;
  wire \DFF_16.D ;
  wire \DFF_16.Q ;
  wire \DFF_160.CK ;
  wire \DFF_160.D ;
  wire \DFF_160.Q ;
  wire \DFF_1600.CK ;
  wire \DFF_1600.D ;
  wire \DFF_1600.Q ;
  wire \DFF_1601.CK ;
  wire \DFF_1601.D ;
  wire \DFF_1601.Q ;
  wire \DFF_1602.CK ;
  wire \DFF_1602.D ;
  wire \DFF_1602.Q ;
  wire \DFF_1603.CK ;
  wire \DFF_1603.D ;
  wire \DFF_1603.Q ;
  wire \DFF_1604.CK ;
  wire \DFF_1604.D ;
  wire \DFF_1604.Q ;
  wire \DFF_1605.CK ;
  wire \DFF_1605.D ;
  wire \DFF_1605.Q ;
  wire \DFF_1606.CK ;
  wire \DFF_1606.D ;
  wire \DFF_1606.Q ;
  wire \DFF_1607.CK ;
  wire \DFF_1607.D ;
  wire \DFF_1607.Q ;
  wire \DFF_1608.CK ;
  wire \DFF_1608.D ;
  wire \DFF_1608.Q ;
  wire \DFF_1609.CK ;
  wire \DFF_1609.D ;
  wire \DFF_1609.Q ;
  wire \DFF_161.CK ;
  wire \DFF_161.D ;
  wire \DFF_161.Q ;
  wire \DFF_1610.CK ;
  wire \DFF_1610.D ;
  wire \DFF_1610.Q ;
  wire \DFF_1611.CK ;
  wire \DFF_1611.D ;
  wire \DFF_1611.Q ;
  wire \DFF_1612.CK ;
  wire \DFF_1612.D ;
  wire \DFF_1612.Q ;
  wire \DFF_1613.CK ;
  wire \DFF_1613.D ;
  wire \DFF_1613.Q ;
  wire \DFF_1614.CK ;
  wire \DFF_1614.D ;
  wire \DFF_1614.Q ;
  wire \DFF_1615.CK ;
  wire \DFF_1615.D ;
  wire \DFF_1615.Q ;
  wire \DFF_1616.CK ;
  wire \DFF_1616.D ;
  wire \DFF_1616.Q ;
  wire \DFF_1617.CK ;
  wire \DFF_1617.D ;
  wire \DFF_1617.Q ;
  wire \DFF_1618.CK ;
  wire \DFF_1618.D ;
  wire \DFF_1618.Q ;
  wire \DFF_1619.CK ;
  wire \DFF_1619.D ;
  wire \DFF_1619.Q ;
  wire \DFF_162.CK ;
  wire \DFF_162.D ;
  wire \DFF_162.Q ;
  wire \DFF_1620.CK ;
  wire \DFF_1620.D ;
  wire \DFF_1620.Q ;
  wire \DFF_1621.CK ;
  wire \DFF_1621.D ;
  wire \DFF_1621.Q ;
  wire \DFF_1622.CK ;
  wire \DFF_1622.D ;
  wire \DFF_1622.Q ;
  wire \DFF_1623.CK ;
  wire \DFF_1623.D ;
  wire \DFF_1623.Q ;
  wire \DFF_1624.CK ;
  wire \DFF_1624.D ;
  wire \DFF_1624.Q ;
  wire \DFF_1625.CK ;
  wire \DFF_1625.D ;
  wire \DFF_1625.Q ;
  wire \DFF_1626.CK ;
  wire \DFF_1626.D ;
  wire \DFF_1626.Q ;
  wire \DFF_1627.CK ;
  wire \DFF_1627.D ;
  wire \DFF_1627.Q ;
  wire \DFF_1628.CK ;
  wire \DFF_1628.D ;
  wire \DFF_1628.Q ;
  wire \DFF_1629.CK ;
  wire \DFF_1629.D ;
  wire \DFF_1629.Q ;
  wire \DFF_163.CK ;
  wire \DFF_163.D ;
  wire \DFF_163.Q ;
  wire \DFF_1630.CK ;
  wire \DFF_1630.D ;
  wire \DFF_1630.Q ;
  wire \DFF_1631.CK ;
  wire \DFF_1631.D ;
  wire \DFF_1631.Q ;
  wire \DFF_1632.CK ;
  wire \DFF_1632.D ;
  wire \DFF_1632.Q ;
  wire \DFF_1633.CK ;
  wire \DFF_1633.D ;
  wire \DFF_1633.Q ;
  wire \DFF_1634.CK ;
  wire \DFF_1634.D ;
  wire \DFF_1634.Q ;
  wire \DFF_1635.CK ;
  wire \DFF_1635.D ;
  wire \DFF_1635.Q ;
  wire \DFF_1636.CK ;
  wire \DFF_1636.D ;
  wire \DFF_1636.Q ;
  wire \DFF_1637.CK ;
  wire \DFF_1637.D ;
  wire \DFF_1637.Q ;
  wire \DFF_1638.CK ;
  wire \DFF_1638.D ;
  wire \DFF_1638.Q ;
  wire \DFF_1639.CK ;
  wire \DFF_1639.D ;
  wire \DFF_1639.Q ;
  wire \DFF_164.CK ;
  wire \DFF_164.D ;
  wire \DFF_164.Q ;
  wire \DFF_1640.CK ;
  wire \DFF_1640.D ;
  wire \DFF_1640.Q ;
  wire \DFF_1641.CK ;
  wire \DFF_1641.D ;
  wire \DFF_1641.Q ;
  wire \DFF_1642.CK ;
  wire \DFF_1642.D ;
  wire \DFF_1642.Q ;
  wire \DFF_1643.CK ;
  wire \DFF_1643.D ;
  wire \DFF_1643.Q ;
  wire \DFF_1644.CK ;
  wire \DFF_1644.D ;
  wire \DFF_1644.Q ;
  wire \DFF_1645.CK ;
  wire \DFF_1645.D ;
  wire \DFF_1645.Q ;
  wire \DFF_1646.CK ;
  wire \DFF_1646.D ;
  wire \DFF_1646.Q ;
  wire \DFF_1647.CK ;
  wire \DFF_1647.D ;
  wire \DFF_1647.Q ;
  wire \DFF_1648.CK ;
  wire \DFF_1648.D ;
  wire \DFF_1648.Q ;
  wire \DFF_1649.CK ;
  wire \DFF_1649.D ;
  wire \DFF_1649.Q ;
  wire \DFF_165.CK ;
  wire \DFF_165.D ;
  wire \DFF_165.Q ;
  wire \DFF_1650.CK ;
  wire \DFF_1650.D ;
  wire \DFF_1650.Q ;
  wire \DFF_1651.CK ;
  wire \DFF_1651.D ;
  wire \DFF_1651.Q ;
  wire \DFF_1652.CK ;
  wire \DFF_1652.D ;
  wire \DFF_1652.Q ;
  wire \DFF_1653.CK ;
  wire \DFF_1653.D ;
  wire \DFF_1653.Q ;
  wire \DFF_1654.CK ;
  wire \DFF_1654.D ;
  wire \DFF_1654.Q ;
  wire \DFF_1655.CK ;
  wire \DFF_1655.D ;
  wire \DFF_1655.Q ;
  wire \DFF_1656.CK ;
  wire \DFF_1656.D ;
  wire \DFF_1656.Q ;
  wire \DFF_1657.CK ;
  wire \DFF_1657.D ;
  wire \DFF_1657.Q ;
  wire \DFF_1658.CK ;
  wire \DFF_1658.D ;
  wire \DFF_1658.Q ;
  wire \DFF_1659.CK ;
  wire \DFF_1659.D ;
  wire \DFF_1659.Q ;
  wire \DFF_166.CK ;
  wire \DFF_166.D ;
  wire \DFF_166.Q ;
  wire \DFF_1660.CK ;
  wire \DFF_1660.D ;
  wire \DFF_1660.Q ;
  wire \DFF_1661.CK ;
  wire \DFF_1661.D ;
  wire \DFF_1661.Q ;
  wire \DFF_1662.CK ;
  wire \DFF_1662.D ;
  wire \DFF_1662.Q ;
  wire \DFF_1663.CK ;
  wire \DFF_1663.D ;
  wire \DFF_1663.Q ;
  wire \DFF_1664.CK ;
  wire \DFF_1664.D ;
  wire \DFF_1664.Q ;
  wire \DFF_1665.CK ;
  wire \DFF_1665.D ;
  wire \DFF_1665.Q ;
  wire \DFF_1666.CK ;
  wire \DFF_1666.D ;
  wire \DFF_1666.Q ;
  wire \DFF_1667.CK ;
  wire \DFF_1667.D ;
  wire \DFF_1667.Q ;
  wire \DFF_1668.CK ;
  wire \DFF_1668.D ;
  wire \DFF_1668.Q ;
  wire \DFF_1669.CK ;
  wire \DFF_1669.D ;
  wire \DFF_1669.Q ;
  wire \DFF_167.CK ;
  wire \DFF_167.D ;
  wire \DFF_167.Q ;
  wire \DFF_1670.CK ;
  wire \DFF_1670.D ;
  wire \DFF_1670.Q ;
  wire \DFF_1671.CK ;
  wire \DFF_1671.D ;
  wire \DFF_1671.Q ;
  wire \DFF_1672.CK ;
  wire \DFF_1672.D ;
  wire \DFF_1672.Q ;
  wire \DFF_1673.CK ;
  wire \DFF_1673.D ;
  wire \DFF_1673.Q ;
  wire \DFF_1674.CK ;
  wire \DFF_1674.D ;
  wire \DFF_1674.Q ;
  wire \DFF_1675.CK ;
  wire \DFF_1675.D ;
  wire \DFF_1675.Q ;
  wire \DFF_1676.CK ;
  wire \DFF_1676.D ;
  wire \DFF_1676.Q ;
  wire \DFF_1677.CK ;
  wire \DFF_1677.D ;
  wire \DFF_1677.Q ;
  wire \DFF_1678.CK ;
  wire \DFF_1678.D ;
  wire \DFF_1678.Q ;
  wire \DFF_1679.CK ;
  wire \DFF_1679.D ;
  wire \DFF_1679.Q ;
  wire \DFF_168.CK ;
  wire \DFF_168.D ;
  wire \DFF_168.Q ;
  wire \DFF_1680.CK ;
  wire \DFF_1680.D ;
  wire \DFF_1680.Q ;
  wire \DFF_1681.CK ;
  wire \DFF_1681.D ;
  wire \DFF_1681.Q ;
  wire \DFF_1682.CK ;
  wire \DFF_1682.D ;
  wire \DFF_1682.Q ;
  wire \DFF_1683.CK ;
  wire \DFF_1683.D ;
  wire \DFF_1683.Q ;
  wire \DFF_1684.CK ;
  wire \DFF_1684.D ;
  wire \DFF_1684.Q ;
  wire \DFF_1685.CK ;
  wire \DFF_1685.D ;
  wire \DFF_1685.Q ;
  wire \DFF_1686.CK ;
  wire \DFF_1686.D ;
  wire \DFF_1686.Q ;
  wire \DFF_1687.CK ;
  wire \DFF_1687.D ;
  wire \DFF_1687.Q ;
  wire \DFF_1688.CK ;
  wire \DFF_1688.D ;
  wire \DFF_1688.Q ;
  wire \DFF_1689.CK ;
  wire \DFF_1689.D ;
  wire \DFF_1689.Q ;
  wire \DFF_169.CK ;
  wire \DFF_169.D ;
  wire \DFF_169.Q ;
  wire \DFF_1690.CK ;
  wire \DFF_1690.D ;
  wire \DFF_1690.Q ;
  wire \DFF_1691.CK ;
  wire \DFF_1691.D ;
  wire \DFF_1691.Q ;
  wire \DFF_1692.CK ;
  wire \DFF_1692.D ;
  wire \DFF_1692.Q ;
  wire \DFF_1693.CK ;
  wire \DFF_1693.D ;
  wire \DFF_1693.Q ;
  wire \DFF_1694.CK ;
  wire \DFF_1694.D ;
  wire \DFF_1694.Q ;
  wire \DFF_1695.CK ;
  wire \DFF_1695.D ;
  wire \DFF_1695.Q ;
  wire \DFF_1696.CK ;
  wire \DFF_1696.D ;
  wire \DFF_1696.Q ;
  wire \DFF_1697.CK ;
  wire \DFF_1697.D ;
  wire \DFF_1697.Q ;
  wire \DFF_1698.CK ;
  wire \DFF_1698.D ;
  wire \DFF_1698.Q ;
  wire \DFF_1699.CK ;
  wire \DFF_1699.D ;
  wire \DFF_1699.Q ;
  wire \DFF_17.CK ;
  wire \DFF_17.D ;
  wire \DFF_17.Q ;
  wire \DFF_170.CK ;
  wire \DFF_170.D ;
  wire \DFF_170.Q ;
  wire \DFF_1700.CK ;
  wire \DFF_1700.D ;
  wire \DFF_1700.Q ;
  wire \DFF_1701.CK ;
  wire \DFF_1701.D ;
  wire \DFF_1701.Q ;
  wire \DFF_1702.CK ;
  wire \DFF_1702.D ;
  wire \DFF_1702.Q ;
  wire \DFF_1703.CK ;
  wire \DFF_1703.D ;
  wire \DFF_1703.Q ;
  wire \DFF_1704.CK ;
  wire \DFF_1704.D ;
  wire \DFF_1704.Q ;
  wire \DFF_1705.CK ;
  wire \DFF_1705.D ;
  wire \DFF_1705.Q ;
  wire \DFF_1706.CK ;
  wire \DFF_1706.D ;
  wire \DFF_1706.Q ;
  wire \DFF_1707.CK ;
  wire \DFF_1707.D ;
  wire \DFF_1707.Q ;
  wire \DFF_1708.CK ;
  wire \DFF_1708.D ;
  wire \DFF_1708.Q ;
  wire \DFF_1709.CK ;
  wire \DFF_1709.D ;
  wire \DFF_1709.Q ;
  wire \DFF_171.CK ;
  wire \DFF_171.D ;
  wire \DFF_171.Q ;
  wire \DFF_1710.CK ;
  wire \DFF_1710.D ;
  wire \DFF_1710.Q ;
  wire \DFF_1711.CK ;
  wire \DFF_1711.D ;
  wire \DFF_1711.Q ;
  wire \DFF_1712.CK ;
  wire \DFF_1712.D ;
  wire \DFF_1712.Q ;
  wire \DFF_1713.CK ;
  wire \DFF_1713.D ;
  wire \DFF_1713.Q ;
  wire \DFF_1714.CK ;
  wire \DFF_1714.D ;
  wire \DFF_1714.Q ;
  wire \DFF_1715.CK ;
  wire \DFF_1715.D ;
  wire \DFF_1715.Q ;
  wire \DFF_1716.CK ;
  wire \DFF_1716.D ;
  wire \DFF_1716.Q ;
  wire \DFF_1717.CK ;
  wire \DFF_1717.D ;
  wire \DFF_1717.Q ;
  wire \DFF_1718.CK ;
  wire \DFF_1718.D ;
  wire \DFF_1718.Q ;
  wire \DFF_1719.CK ;
  wire \DFF_1719.D ;
  wire \DFF_1719.Q ;
  wire \DFF_172.CK ;
  wire \DFF_172.D ;
  wire \DFF_172.Q ;
  wire \DFF_1720.CK ;
  wire \DFF_1720.D ;
  wire \DFF_1720.Q ;
  wire \DFF_1721.CK ;
  wire \DFF_1721.D ;
  wire \DFF_1721.Q ;
  wire \DFF_1722.CK ;
  wire \DFF_1722.D ;
  wire \DFF_1722.Q ;
  wire \DFF_1723.CK ;
  wire \DFF_1723.D ;
  wire \DFF_1723.Q ;
  wire \DFF_1724.CK ;
  wire \DFF_1724.D ;
  wire \DFF_1724.Q ;
  wire \DFF_1725.CK ;
  wire \DFF_1725.D ;
  wire \DFF_1725.Q ;
  wire \DFF_1726.CK ;
  wire \DFF_1726.D ;
  wire \DFF_1726.Q ;
  wire \DFF_1727.CK ;
  wire \DFF_1727.D ;
  wire \DFF_1727.Q ;
  wire \DFF_173.CK ;
  wire \DFF_173.D ;
  wire \DFF_173.Q ;
  wire \DFF_174.CK ;
  wire \DFF_174.D ;
  wire \DFF_174.Q ;
  wire \DFF_175.CK ;
  wire \DFF_175.D ;
  wire \DFF_175.Q ;
  wire \DFF_176.CK ;
  wire \DFF_176.D ;
  wire \DFF_176.Q ;
  wire \DFF_177.CK ;
  wire \DFF_177.D ;
  wire \DFF_177.Q ;
  wire \DFF_178.CK ;
  wire \DFF_178.D ;
  wire \DFF_178.Q ;
  wire \DFF_179.CK ;
  wire \DFF_179.D ;
  wire \DFF_179.Q ;
  wire \DFF_18.CK ;
  wire \DFF_18.D ;
  wire \DFF_18.Q ;
  wire \DFF_180.CK ;
  wire \DFF_180.D ;
  wire \DFF_180.Q ;
  wire \DFF_181.CK ;
  wire \DFF_181.D ;
  wire \DFF_181.Q ;
  wire \DFF_182.CK ;
  wire \DFF_182.D ;
  wire \DFF_182.Q ;
  wire \DFF_183.CK ;
  wire \DFF_183.D ;
  wire \DFF_183.Q ;
  wire \DFF_184.CK ;
  wire \DFF_184.D ;
  wire \DFF_184.Q ;
  wire \DFF_185.CK ;
  wire \DFF_185.D ;
  wire \DFF_185.Q ;
  wire \DFF_186.CK ;
  wire \DFF_186.D ;
  wire \DFF_186.Q ;
  wire \DFF_187.CK ;
  wire \DFF_187.D ;
  wire \DFF_187.Q ;
  wire \DFF_188.CK ;
  wire \DFF_188.D ;
  wire \DFF_188.Q ;
  wire \DFF_189.CK ;
  wire \DFF_189.D ;
  wire \DFF_189.Q ;
  wire \DFF_19.CK ;
  wire \DFF_19.D ;
  wire \DFF_19.Q ;
  wire \DFF_190.CK ;
  wire \DFF_190.D ;
  wire \DFF_190.Q ;
  wire \DFF_191.CK ;
  wire \DFF_191.D ;
  wire \DFF_191.Q ;
  wire \DFF_192.CK ;
  wire \DFF_192.D ;
  wire \DFF_192.Q ;
  wire \DFF_193.CK ;
  wire \DFF_193.D ;
  wire \DFF_193.Q ;
  wire \DFF_194.CK ;
  wire \DFF_194.D ;
  wire \DFF_194.Q ;
  wire \DFF_195.CK ;
  wire \DFF_195.D ;
  wire \DFF_195.Q ;
  wire \DFF_196.CK ;
  wire \DFF_196.D ;
  wire \DFF_196.Q ;
  wire \DFF_197.CK ;
  wire \DFF_197.D ;
  wire \DFF_197.Q ;
  wire \DFF_198.CK ;
  wire \DFF_198.D ;
  wire \DFF_198.Q ;
  wire \DFF_199.CK ;
  wire \DFF_199.D ;
  wire \DFF_199.Q ;
  wire \DFF_2.CK ;
  wire \DFF_2.D ;
  wire \DFF_2.Q ;
  wire \DFF_20.CK ;
  wire \DFF_20.D ;
  wire \DFF_20.Q ;
  wire \DFF_200.CK ;
  wire \DFF_200.D ;
  wire \DFF_200.Q ;
  wire \DFF_201.CK ;
  wire \DFF_201.D ;
  wire \DFF_201.Q ;
  wire \DFF_202.CK ;
  wire \DFF_202.D ;
  wire \DFF_202.Q ;
  wire \DFF_203.CK ;
  wire \DFF_203.D ;
  wire \DFF_203.Q ;
  wire \DFF_204.CK ;
  wire \DFF_204.D ;
  wire \DFF_204.Q ;
  wire \DFF_205.CK ;
  wire \DFF_205.D ;
  wire \DFF_205.Q ;
  wire \DFF_206.CK ;
  wire \DFF_206.D ;
  wire \DFF_206.Q ;
  wire \DFF_207.CK ;
  wire \DFF_207.D ;
  wire \DFF_207.Q ;
  wire \DFF_208.CK ;
  wire \DFF_208.D ;
  wire \DFF_208.Q ;
  wire \DFF_209.CK ;
  wire \DFF_209.D ;
  wire \DFF_209.Q ;
  wire \DFF_21.CK ;
  wire \DFF_21.D ;
  wire \DFF_21.Q ;
  wire \DFF_210.CK ;
  wire \DFF_210.D ;
  wire \DFF_210.Q ;
  wire \DFF_211.CK ;
  wire \DFF_211.D ;
  wire \DFF_211.Q ;
  wire \DFF_212.CK ;
  wire \DFF_212.D ;
  wire \DFF_212.Q ;
  wire \DFF_213.CK ;
  wire \DFF_213.D ;
  wire \DFF_213.Q ;
  wire \DFF_214.CK ;
  wire \DFF_214.D ;
  wire \DFF_214.Q ;
  wire \DFF_215.CK ;
  wire \DFF_215.D ;
  wire \DFF_215.Q ;
  wire \DFF_216.CK ;
  wire \DFF_216.D ;
  wire \DFF_216.Q ;
  wire \DFF_217.CK ;
  wire \DFF_217.D ;
  wire \DFF_217.Q ;
  wire \DFF_218.CK ;
  wire \DFF_218.D ;
  wire \DFF_218.Q ;
  wire \DFF_219.CK ;
  wire \DFF_219.D ;
  wire \DFF_219.Q ;
  wire \DFF_22.CK ;
  wire \DFF_22.D ;
  wire \DFF_22.Q ;
  wire \DFF_220.CK ;
  wire \DFF_220.D ;
  wire \DFF_220.Q ;
  wire \DFF_221.CK ;
  wire \DFF_221.D ;
  wire \DFF_221.Q ;
  wire \DFF_222.CK ;
  wire \DFF_222.D ;
  wire \DFF_222.Q ;
  wire \DFF_223.CK ;
  wire \DFF_223.D ;
  wire \DFF_223.Q ;
  wire \DFF_224.CK ;
  wire \DFF_224.D ;
  wire \DFF_224.Q ;
  wire \DFF_225.CK ;
  wire \DFF_225.D ;
  wire \DFF_225.Q ;
  wire \DFF_226.CK ;
  wire \DFF_226.D ;
  wire \DFF_226.Q ;
  wire \DFF_227.CK ;
  wire \DFF_227.D ;
  wire \DFF_227.Q ;
  wire \DFF_228.CK ;
  wire \DFF_228.D ;
  wire \DFF_228.Q ;
  wire \DFF_229.CK ;
  wire \DFF_229.D ;
  wire \DFF_229.Q ;
  wire \DFF_23.CK ;
  wire \DFF_23.D ;
  wire \DFF_23.Q ;
  wire \DFF_230.CK ;
  wire \DFF_230.D ;
  wire \DFF_230.Q ;
  wire \DFF_231.CK ;
  wire \DFF_231.D ;
  wire \DFF_231.Q ;
  wire \DFF_232.CK ;
  wire \DFF_232.D ;
  wire \DFF_232.Q ;
  wire \DFF_233.CK ;
  wire \DFF_233.D ;
  wire \DFF_233.Q ;
  wire \DFF_234.CK ;
  wire \DFF_234.D ;
  wire \DFF_234.Q ;
  wire \DFF_235.CK ;
  wire \DFF_235.D ;
  wire \DFF_235.Q ;
  wire \DFF_236.CK ;
  wire \DFF_236.D ;
  wire \DFF_236.Q ;
  wire \DFF_237.CK ;
  wire \DFF_237.D ;
  wire \DFF_237.Q ;
  wire \DFF_238.CK ;
  wire \DFF_238.D ;
  wire \DFF_238.Q ;
  wire \DFF_239.CK ;
  wire \DFF_239.D ;
  wire \DFF_239.Q ;
  wire \DFF_24.CK ;
  wire \DFF_24.D ;
  wire \DFF_24.Q ;
  wire \DFF_240.CK ;
  wire \DFF_240.D ;
  wire \DFF_240.Q ;
  wire \DFF_241.CK ;
  wire \DFF_241.D ;
  wire \DFF_241.Q ;
  wire \DFF_242.CK ;
  wire \DFF_242.D ;
  wire \DFF_242.Q ;
  wire \DFF_243.CK ;
  wire \DFF_243.D ;
  wire \DFF_243.Q ;
  wire \DFF_244.CK ;
  wire \DFF_244.D ;
  wire \DFF_244.Q ;
  wire \DFF_245.CK ;
  wire \DFF_245.D ;
  wire \DFF_245.Q ;
  wire \DFF_246.CK ;
  wire \DFF_246.D ;
  wire \DFF_246.Q ;
  wire \DFF_247.CK ;
  wire \DFF_247.D ;
  wire \DFF_247.Q ;
  wire \DFF_248.CK ;
  wire \DFF_248.D ;
  wire \DFF_248.Q ;
  wire \DFF_249.CK ;
  wire \DFF_249.D ;
  wire \DFF_249.Q ;
  wire \DFF_25.CK ;
  wire \DFF_25.D ;
  wire \DFF_25.Q ;
  wire \DFF_250.CK ;
  wire \DFF_250.D ;
  wire \DFF_250.Q ;
  wire \DFF_251.CK ;
  wire \DFF_251.D ;
  wire \DFF_251.Q ;
  wire \DFF_252.CK ;
  wire \DFF_252.D ;
  wire \DFF_252.Q ;
  wire \DFF_253.CK ;
  wire \DFF_253.D ;
  wire \DFF_253.Q ;
  wire \DFF_254.CK ;
  wire \DFF_254.D ;
  wire \DFF_254.Q ;
  wire \DFF_255.CK ;
  wire \DFF_255.D ;
  wire \DFF_255.Q ;
  wire \DFF_256.CK ;
  wire \DFF_256.D ;
  wire \DFF_256.Q ;
  wire \DFF_257.CK ;
  wire \DFF_257.D ;
  wire \DFF_257.Q ;
  wire \DFF_258.CK ;
  wire \DFF_258.D ;
  wire \DFF_258.Q ;
  wire \DFF_259.CK ;
  wire \DFF_259.D ;
  wire \DFF_259.Q ;
  wire \DFF_26.CK ;
  wire \DFF_26.D ;
  wire \DFF_26.Q ;
  wire \DFF_260.CK ;
  wire \DFF_260.D ;
  wire \DFF_260.Q ;
  wire \DFF_261.CK ;
  wire \DFF_261.D ;
  wire \DFF_261.Q ;
  wire \DFF_262.CK ;
  wire \DFF_262.D ;
  wire \DFF_262.Q ;
  wire \DFF_263.CK ;
  wire \DFF_263.D ;
  wire \DFF_263.Q ;
  wire \DFF_264.CK ;
  wire \DFF_264.D ;
  wire \DFF_264.Q ;
  wire \DFF_265.CK ;
  wire \DFF_265.D ;
  wire \DFF_265.Q ;
  wire \DFF_266.CK ;
  wire \DFF_266.D ;
  wire \DFF_266.Q ;
  wire \DFF_267.CK ;
  wire \DFF_267.D ;
  wire \DFF_267.Q ;
  wire \DFF_268.CK ;
  wire \DFF_268.D ;
  wire \DFF_268.Q ;
  wire \DFF_269.CK ;
  wire \DFF_269.D ;
  wire \DFF_269.Q ;
  wire \DFF_27.CK ;
  wire \DFF_27.D ;
  wire \DFF_27.Q ;
  wire \DFF_270.CK ;
  wire \DFF_270.D ;
  wire \DFF_270.Q ;
  wire \DFF_271.CK ;
  wire \DFF_271.D ;
  wire \DFF_271.Q ;
  wire \DFF_272.CK ;
  wire \DFF_272.D ;
  wire \DFF_272.Q ;
  wire \DFF_273.CK ;
  wire \DFF_273.D ;
  wire \DFF_273.Q ;
  wire \DFF_274.CK ;
  wire \DFF_274.D ;
  wire \DFF_274.Q ;
  wire \DFF_275.CK ;
  wire \DFF_275.D ;
  wire \DFF_275.Q ;
  wire \DFF_276.CK ;
  wire \DFF_276.D ;
  wire \DFF_276.Q ;
  wire \DFF_277.CK ;
  wire \DFF_277.D ;
  wire \DFF_277.Q ;
  wire \DFF_278.CK ;
  wire \DFF_278.D ;
  wire \DFF_278.Q ;
  wire \DFF_279.CK ;
  wire \DFF_279.D ;
  wire \DFF_279.Q ;
  wire \DFF_28.CK ;
  wire \DFF_28.D ;
  wire \DFF_28.Q ;
  wire \DFF_280.CK ;
  wire \DFF_280.D ;
  wire \DFF_280.Q ;
  wire \DFF_281.CK ;
  wire \DFF_281.D ;
  wire \DFF_281.Q ;
  wire \DFF_282.CK ;
  wire \DFF_282.D ;
  wire \DFF_282.Q ;
  wire \DFF_283.CK ;
  wire \DFF_283.D ;
  wire \DFF_283.Q ;
  wire \DFF_284.CK ;
  wire \DFF_284.D ;
  wire \DFF_284.Q ;
  wire \DFF_285.CK ;
  wire \DFF_285.D ;
  wire \DFF_285.Q ;
  wire \DFF_286.CK ;
  wire \DFF_286.D ;
  wire \DFF_286.Q ;
  wire \DFF_287.CK ;
  wire \DFF_287.D ;
  wire \DFF_287.Q ;
  wire \DFF_288.CK ;
  wire \DFF_288.D ;
  wire \DFF_288.Q ;
  wire \DFF_289.CK ;
  wire \DFF_289.D ;
  wire \DFF_289.Q ;
  wire \DFF_29.CK ;
  wire \DFF_29.D ;
  wire \DFF_29.Q ;
  wire \DFF_290.CK ;
  wire \DFF_290.D ;
  wire \DFF_290.Q ;
  wire \DFF_291.CK ;
  wire \DFF_291.D ;
  wire \DFF_291.Q ;
  wire \DFF_292.CK ;
  wire \DFF_292.D ;
  wire \DFF_292.Q ;
  wire \DFF_293.CK ;
  wire \DFF_293.D ;
  wire \DFF_293.Q ;
  wire \DFF_294.CK ;
  wire \DFF_294.D ;
  wire \DFF_294.Q ;
  wire \DFF_295.CK ;
  wire \DFF_295.D ;
  wire \DFF_295.Q ;
  wire \DFF_296.CK ;
  wire \DFF_296.D ;
  wire \DFF_296.Q ;
  wire \DFF_297.CK ;
  wire \DFF_297.D ;
  wire \DFF_297.Q ;
  wire \DFF_298.CK ;
  wire \DFF_298.D ;
  wire \DFF_298.Q ;
  wire \DFF_299.CK ;
  wire \DFF_299.D ;
  wire \DFF_299.Q ;
  wire \DFF_3.CK ;
  wire \DFF_3.D ;
  wire \DFF_3.Q ;
  wire \DFF_30.CK ;
  wire \DFF_30.D ;
  wire \DFF_30.Q ;
  wire \DFF_300.CK ;
  wire \DFF_300.D ;
  wire \DFF_300.Q ;
  wire \DFF_301.CK ;
  wire \DFF_301.D ;
  wire \DFF_301.Q ;
  wire \DFF_302.CK ;
  wire \DFF_302.D ;
  wire \DFF_302.Q ;
  wire \DFF_303.CK ;
  wire \DFF_303.D ;
  wire \DFF_303.Q ;
  wire \DFF_304.CK ;
  wire \DFF_304.D ;
  wire \DFF_304.Q ;
  wire \DFF_305.CK ;
  wire \DFF_305.D ;
  wire \DFF_305.Q ;
  wire \DFF_306.CK ;
  wire \DFF_306.D ;
  wire \DFF_306.Q ;
  wire \DFF_307.CK ;
  wire \DFF_307.D ;
  wire \DFF_307.Q ;
  wire \DFF_308.CK ;
  wire \DFF_308.D ;
  wire \DFF_308.Q ;
  wire \DFF_309.CK ;
  wire \DFF_309.D ;
  wire \DFF_309.Q ;
  wire \DFF_31.CK ;
  wire \DFF_31.D ;
  wire \DFF_31.Q ;
  wire \DFF_310.CK ;
  wire \DFF_310.D ;
  wire \DFF_310.Q ;
  wire \DFF_311.CK ;
  wire \DFF_311.D ;
  wire \DFF_311.Q ;
  wire \DFF_312.CK ;
  wire \DFF_312.D ;
  wire \DFF_312.Q ;
  wire \DFF_313.CK ;
  wire \DFF_313.D ;
  wire \DFF_313.Q ;
  wire \DFF_314.CK ;
  wire \DFF_314.D ;
  wire \DFF_314.Q ;
  wire \DFF_315.CK ;
  wire \DFF_315.D ;
  wire \DFF_315.Q ;
  wire \DFF_316.CK ;
  wire \DFF_316.D ;
  wire \DFF_316.Q ;
  wire \DFF_317.CK ;
  wire \DFF_317.D ;
  wire \DFF_317.Q ;
  wire \DFF_318.CK ;
  wire \DFF_318.D ;
  wire \DFF_318.Q ;
  wire \DFF_319.CK ;
  wire \DFF_319.D ;
  wire \DFF_319.Q ;
  wire \DFF_32.CK ;
  wire \DFF_32.D ;
  wire \DFF_32.Q ;
  wire \DFF_320.CK ;
  wire \DFF_320.D ;
  wire \DFF_320.Q ;
  wire \DFF_321.CK ;
  wire \DFF_321.D ;
  wire \DFF_321.Q ;
  wire \DFF_322.CK ;
  wire \DFF_322.D ;
  wire \DFF_322.Q ;
  wire \DFF_323.CK ;
  wire \DFF_323.D ;
  wire \DFF_323.Q ;
  wire \DFF_324.CK ;
  wire \DFF_324.D ;
  wire \DFF_324.Q ;
  wire \DFF_325.CK ;
  wire \DFF_325.D ;
  wire \DFF_325.Q ;
  wire \DFF_326.CK ;
  wire \DFF_326.D ;
  wire \DFF_326.Q ;
  wire \DFF_327.CK ;
  wire \DFF_327.D ;
  wire \DFF_327.Q ;
  wire \DFF_328.CK ;
  wire \DFF_328.D ;
  wire \DFF_328.Q ;
  wire \DFF_329.CK ;
  wire \DFF_329.D ;
  wire \DFF_329.Q ;
  wire \DFF_33.CK ;
  wire \DFF_33.D ;
  wire \DFF_33.Q ;
  wire \DFF_330.CK ;
  wire \DFF_330.D ;
  wire \DFF_330.Q ;
  wire \DFF_331.CK ;
  wire \DFF_331.D ;
  wire \DFF_331.Q ;
  wire \DFF_332.CK ;
  wire \DFF_332.D ;
  wire \DFF_332.Q ;
  wire \DFF_333.CK ;
  wire \DFF_333.D ;
  wire \DFF_333.Q ;
  wire \DFF_334.CK ;
  wire \DFF_334.D ;
  wire \DFF_334.Q ;
  wire \DFF_335.CK ;
  wire \DFF_335.D ;
  wire \DFF_335.Q ;
  wire \DFF_336.CK ;
  wire \DFF_336.D ;
  wire \DFF_336.Q ;
  wire \DFF_337.CK ;
  wire \DFF_337.D ;
  wire \DFF_337.Q ;
  wire \DFF_338.CK ;
  wire \DFF_338.D ;
  wire \DFF_338.Q ;
  wire \DFF_339.CK ;
  wire \DFF_339.D ;
  wire \DFF_339.Q ;
  wire \DFF_34.CK ;
  wire \DFF_34.D ;
  wire \DFF_34.Q ;
  wire \DFF_340.CK ;
  wire \DFF_340.D ;
  wire \DFF_340.Q ;
  wire \DFF_341.CK ;
  wire \DFF_341.D ;
  wire \DFF_341.Q ;
  wire \DFF_342.CK ;
  wire \DFF_342.D ;
  wire \DFF_342.Q ;
  wire \DFF_343.CK ;
  wire \DFF_343.D ;
  wire \DFF_343.Q ;
  wire \DFF_344.CK ;
  wire \DFF_344.D ;
  wire \DFF_344.Q ;
  wire \DFF_345.CK ;
  wire \DFF_345.D ;
  wire \DFF_345.Q ;
  wire \DFF_346.CK ;
  wire \DFF_346.D ;
  wire \DFF_346.Q ;
  wire \DFF_347.CK ;
  wire \DFF_347.D ;
  wire \DFF_347.Q ;
  wire \DFF_348.CK ;
  wire \DFF_348.D ;
  wire \DFF_348.Q ;
  wire \DFF_349.CK ;
  wire \DFF_349.D ;
  wire \DFF_349.Q ;
  wire \DFF_35.CK ;
  wire \DFF_35.D ;
  wire \DFF_35.Q ;
  wire \DFF_350.CK ;
  wire \DFF_350.D ;
  wire \DFF_350.Q ;
  wire \DFF_351.CK ;
  wire \DFF_351.D ;
  wire \DFF_351.Q ;
  wire \DFF_352.CK ;
  wire \DFF_352.D ;
  wire \DFF_352.Q ;
  wire \DFF_353.CK ;
  wire \DFF_353.D ;
  wire \DFF_353.Q ;
  wire \DFF_354.CK ;
  wire \DFF_354.D ;
  wire \DFF_354.Q ;
  wire \DFF_355.CK ;
  wire \DFF_355.D ;
  wire \DFF_355.Q ;
  wire \DFF_356.CK ;
  wire \DFF_356.D ;
  wire \DFF_356.Q ;
  wire \DFF_357.CK ;
  wire \DFF_357.D ;
  wire \DFF_357.Q ;
  wire \DFF_358.CK ;
  wire \DFF_358.D ;
  wire \DFF_358.Q ;
  wire \DFF_359.CK ;
  wire \DFF_359.D ;
  wire \DFF_359.Q ;
  wire \DFF_36.CK ;
  wire \DFF_36.D ;
  wire \DFF_36.Q ;
  wire \DFF_360.CK ;
  wire \DFF_360.D ;
  wire \DFF_360.Q ;
  wire \DFF_361.CK ;
  wire \DFF_361.D ;
  wire \DFF_361.Q ;
  wire \DFF_362.CK ;
  wire \DFF_362.D ;
  wire \DFF_362.Q ;
  wire \DFF_363.CK ;
  wire \DFF_363.D ;
  wire \DFF_363.Q ;
  wire \DFF_364.CK ;
  wire \DFF_364.D ;
  wire \DFF_364.Q ;
  wire \DFF_365.CK ;
  wire \DFF_365.D ;
  wire \DFF_365.Q ;
  wire \DFF_366.CK ;
  wire \DFF_366.D ;
  wire \DFF_366.Q ;
  wire \DFF_367.CK ;
  wire \DFF_367.D ;
  wire \DFF_367.Q ;
  wire \DFF_368.CK ;
  wire \DFF_368.D ;
  wire \DFF_368.Q ;
  wire \DFF_369.CK ;
  wire \DFF_369.D ;
  wire \DFF_369.Q ;
  wire \DFF_37.CK ;
  wire \DFF_37.D ;
  wire \DFF_37.Q ;
  wire \DFF_370.CK ;
  wire \DFF_370.D ;
  wire \DFF_370.Q ;
  wire \DFF_371.CK ;
  wire \DFF_371.D ;
  wire \DFF_371.Q ;
  wire \DFF_372.CK ;
  wire \DFF_372.D ;
  wire \DFF_372.Q ;
  wire \DFF_373.CK ;
  wire \DFF_373.D ;
  wire \DFF_373.Q ;
  wire \DFF_374.CK ;
  wire \DFF_374.D ;
  wire \DFF_374.Q ;
  wire \DFF_375.CK ;
  wire \DFF_375.D ;
  wire \DFF_375.Q ;
  wire \DFF_376.CK ;
  wire \DFF_376.D ;
  wire \DFF_376.Q ;
  wire \DFF_377.CK ;
  wire \DFF_377.D ;
  wire \DFF_377.Q ;
  wire \DFF_378.CK ;
  wire \DFF_378.D ;
  wire \DFF_378.Q ;
  wire \DFF_379.CK ;
  wire \DFF_379.D ;
  wire \DFF_379.Q ;
  wire \DFF_38.CK ;
  wire \DFF_38.D ;
  wire \DFF_38.Q ;
  wire \DFF_380.CK ;
  wire \DFF_380.D ;
  wire \DFF_380.Q ;
  wire \DFF_381.CK ;
  wire \DFF_381.D ;
  wire \DFF_381.Q ;
  wire \DFF_382.CK ;
  wire \DFF_382.D ;
  wire \DFF_382.Q ;
  wire \DFF_383.CK ;
  wire \DFF_383.D ;
  wire \DFF_383.Q ;
  wire \DFF_384.CK ;
  wire \DFF_384.D ;
  wire \DFF_384.Q ;
  wire \DFF_385.CK ;
  wire \DFF_385.D ;
  wire \DFF_385.Q ;
  wire \DFF_386.CK ;
  wire \DFF_386.D ;
  wire \DFF_386.Q ;
  wire \DFF_387.CK ;
  wire \DFF_387.D ;
  wire \DFF_387.Q ;
  wire \DFF_388.CK ;
  wire \DFF_388.D ;
  wire \DFF_388.Q ;
  wire \DFF_389.CK ;
  wire \DFF_389.D ;
  wire \DFF_389.Q ;
  wire \DFF_39.CK ;
  wire \DFF_39.D ;
  wire \DFF_39.Q ;
  wire \DFF_390.CK ;
  wire \DFF_390.D ;
  wire \DFF_390.Q ;
  wire \DFF_391.CK ;
  wire \DFF_391.D ;
  wire \DFF_391.Q ;
  wire \DFF_392.CK ;
  wire \DFF_392.D ;
  wire \DFF_392.Q ;
  wire \DFF_393.CK ;
  wire \DFF_393.D ;
  wire \DFF_393.Q ;
  wire \DFF_394.CK ;
  wire \DFF_394.D ;
  wire \DFF_394.Q ;
  wire \DFF_395.CK ;
  wire \DFF_395.D ;
  wire \DFF_395.Q ;
  wire \DFF_396.CK ;
  wire \DFF_396.D ;
  wire \DFF_396.Q ;
  wire \DFF_397.CK ;
  wire \DFF_397.D ;
  wire \DFF_397.Q ;
  wire \DFF_398.CK ;
  wire \DFF_398.D ;
  wire \DFF_398.Q ;
  wire \DFF_399.CK ;
  wire \DFF_399.D ;
  wire \DFF_399.Q ;
  wire \DFF_4.CK ;
  wire \DFF_4.D ;
  wire \DFF_4.Q ;
  wire \DFF_40.CK ;
  wire \DFF_40.D ;
  wire \DFF_40.Q ;
  wire \DFF_400.CK ;
  wire \DFF_400.D ;
  wire \DFF_400.Q ;
  wire \DFF_401.CK ;
  wire \DFF_401.D ;
  wire \DFF_401.Q ;
  wire \DFF_402.CK ;
  wire \DFF_402.D ;
  wire \DFF_402.Q ;
  wire \DFF_403.CK ;
  wire \DFF_403.D ;
  wire \DFF_403.Q ;
  wire \DFF_404.CK ;
  wire \DFF_404.D ;
  wire \DFF_404.Q ;
  wire \DFF_405.CK ;
  wire \DFF_405.D ;
  wire \DFF_405.Q ;
  wire \DFF_406.CK ;
  wire \DFF_406.D ;
  wire \DFF_406.Q ;
  wire \DFF_407.CK ;
  wire \DFF_407.D ;
  wire \DFF_407.Q ;
  wire \DFF_408.CK ;
  wire \DFF_408.D ;
  wire \DFF_408.Q ;
  wire \DFF_409.CK ;
  wire \DFF_409.D ;
  wire \DFF_409.Q ;
  wire \DFF_41.CK ;
  wire \DFF_41.D ;
  wire \DFF_41.Q ;
  wire \DFF_410.CK ;
  wire \DFF_410.D ;
  wire \DFF_410.Q ;
  wire \DFF_411.CK ;
  wire \DFF_411.D ;
  wire \DFF_411.Q ;
  wire \DFF_412.CK ;
  wire \DFF_412.D ;
  wire \DFF_412.Q ;
  wire \DFF_413.CK ;
  wire \DFF_413.D ;
  wire \DFF_413.Q ;
  wire \DFF_414.CK ;
  wire \DFF_414.D ;
  wire \DFF_414.Q ;
  wire \DFF_415.CK ;
  wire \DFF_415.D ;
  wire \DFF_415.Q ;
  wire \DFF_416.CK ;
  wire \DFF_416.D ;
  wire \DFF_416.Q ;
  wire \DFF_417.CK ;
  wire \DFF_417.D ;
  wire \DFF_417.Q ;
  wire \DFF_418.CK ;
  wire \DFF_418.D ;
  wire \DFF_418.Q ;
  wire \DFF_419.CK ;
  wire \DFF_419.D ;
  wire \DFF_419.Q ;
  wire \DFF_42.CK ;
  wire \DFF_42.D ;
  wire \DFF_42.Q ;
  wire \DFF_420.CK ;
  wire \DFF_420.D ;
  wire \DFF_420.Q ;
  wire \DFF_421.CK ;
  wire \DFF_421.D ;
  wire \DFF_421.Q ;
  wire \DFF_422.CK ;
  wire \DFF_422.D ;
  wire \DFF_422.Q ;
  wire \DFF_423.CK ;
  wire \DFF_423.D ;
  wire \DFF_423.Q ;
  wire \DFF_424.CK ;
  wire \DFF_424.D ;
  wire \DFF_424.Q ;
  wire \DFF_425.CK ;
  wire \DFF_425.D ;
  wire \DFF_425.Q ;
  wire \DFF_426.CK ;
  wire \DFF_426.D ;
  wire \DFF_426.Q ;
  wire \DFF_427.CK ;
  wire \DFF_427.D ;
  wire \DFF_427.Q ;
  wire \DFF_428.CK ;
  wire \DFF_428.D ;
  wire \DFF_428.Q ;
  wire \DFF_429.CK ;
  wire \DFF_429.D ;
  wire \DFF_429.Q ;
  wire \DFF_43.CK ;
  wire \DFF_43.D ;
  wire \DFF_43.Q ;
  wire \DFF_430.CK ;
  wire \DFF_430.D ;
  wire \DFF_430.Q ;
  wire \DFF_431.CK ;
  wire \DFF_431.D ;
  wire \DFF_431.Q ;
  wire \DFF_432.CK ;
  wire \DFF_432.D ;
  wire \DFF_432.Q ;
  wire \DFF_433.CK ;
  wire \DFF_433.D ;
  wire \DFF_433.Q ;
  wire \DFF_434.CK ;
  wire \DFF_434.D ;
  wire \DFF_434.Q ;
  wire \DFF_435.CK ;
  wire \DFF_435.D ;
  wire \DFF_435.Q ;
  wire \DFF_436.CK ;
  wire \DFF_436.D ;
  wire \DFF_436.Q ;
  wire \DFF_437.CK ;
  wire \DFF_437.D ;
  wire \DFF_437.Q ;
  wire \DFF_438.CK ;
  wire \DFF_438.D ;
  wire \DFF_438.Q ;
  wire \DFF_439.CK ;
  wire \DFF_439.D ;
  wire \DFF_439.Q ;
  wire \DFF_44.CK ;
  wire \DFF_44.D ;
  wire \DFF_44.Q ;
  wire \DFF_440.CK ;
  wire \DFF_440.D ;
  wire \DFF_440.Q ;
  wire \DFF_441.CK ;
  wire \DFF_441.D ;
  wire \DFF_441.Q ;
  wire \DFF_442.CK ;
  wire \DFF_442.D ;
  wire \DFF_442.Q ;
  wire \DFF_443.CK ;
  wire \DFF_443.D ;
  wire \DFF_443.Q ;
  wire \DFF_444.CK ;
  wire \DFF_444.D ;
  wire \DFF_444.Q ;
  wire \DFF_445.CK ;
  wire \DFF_445.D ;
  wire \DFF_445.Q ;
  wire \DFF_446.CK ;
  wire \DFF_446.D ;
  wire \DFF_446.Q ;
  wire \DFF_447.CK ;
  wire \DFF_447.D ;
  wire \DFF_447.Q ;
  wire \DFF_448.CK ;
  wire \DFF_448.D ;
  wire \DFF_448.Q ;
  wire \DFF_449.CK ;
  wire \DFF_449.D ;
  wire \DFF_449.Q ;
  wire \DFF_45.CK ;
  wire \DFF_45.D ;
  wire \DFF_45.Q ;
  wire \DFF_450.CK ;
  wire \DFF_450.D ;
  wire \DFF_450.Q ;
  wire \DFF_451.CK ;
  wire \DFF_451.D ;
  wire \DFF_451.Q ;
  wire \DFF_452.CK ;
  wire \DFF_452.D ;
  wire \DFF_452.Q ;
  wire \DFF_453.CK ;
  wire \DFF_453.D ;
  wire \DFF_453.Q ;
  wire \DFF_454.CK ;
  wire \DFF_454.D ;
  wire \DFF_454.Q ;
  wire \DFF_455.CK ;
  wire \DFF_455.D ;
  wire \DFF_455.Q ;
  wire \DFF_456.CK ;
  wire \DFF_456.D ;
  wire \DFF_456.Q ;
  wire \DFF_457.CK ;
  wire \DFF_457.D ;
  wire \DFF_457.Q ;
  wire \DFF_458.CK ;
  wire \DFF_458.D ;
  wire \DFF_458.Q ;
  wire \DFF_459.CK ;
  wire \DFF_459.D ;
  wire \DFF_459.Q ;
  wire \DFF_46.CK ;
  wire \DFF_46.D ;
  wire \DFF_46.Q ;
  wire \DFF_460.CK ;
  wire \DFF_460.D ;
  wire \DFF_460.Q ;
  wire \DFF_461.CK ;
  wire \DFF_461.D ;
  wire \DFF_461.Q ;
  wire \DFF_462.CK ;
  wire \DFF_462.D ;
  wire \DFF_462.Q ;
  wire \DFF_463.CK ;
  wire \DFF_463.D ;
  wire \DFF_463.Q ;
  wire \DFF_464.CK ;
  wire \DFF_464.D ;
  wire \DFF_464.Q ;
  wire \DFF_465.CK ;
  wire \DFF_465.D ;
  wire \DFF_465.Q ;
  wire \DFF_466.CK ;
  wire \DFF_466.D ;
  wire \DFF_466.Q ;
  wire \DFF_467.CK ;
  wire \DFF_467.D ;
  wire \DFF_467.Q ;
  wire \DFF_468.CK ;
  wire \DFF_468.D ;
  wire \DFF_468.Q ;
  wire \DFF_469.CK ;
  wire \DFF_469.D ;
  wire \DFF_469.Q ;
  wire \DFF_47.CK ;
  wire \DFF_47.D ;
  wire \DFF_47.Q ;
  wire \DFF_470.CK ;
  wire \DFF_470.D ;
  wire \DFF_470.Q ;
  wire \DFF_471.CK ;
  wire \DFF_471.D ;
  wire \DFF_471.Q ;
  wire \DFF_472.CK ;
  wire \DFF_472.D ;
  wire \DFF_472.Q ;
  wire \DFF_473.CK ;
  wire \DFF_473.D ;
  wire \DFF_473.Q ;
  wire \DFF_474.CK ;
  wire \DFF_474.D ;
  wire \DFF_474.Q ;
  wire \DFF_475.CK ;
  wire \DFF_475.D ;
  wire \DFF_475.Q ;
  wire \DFF_476.CK ;
  wire \DFF_476.D ;
  wire \DFF_476.Q ;
  wire \DFF_477.CK ;
  wire \DFF_477.D ;
  wire \DFF_477.Q ;
  wire \DFF_478.CK ;
  wire \DFF_478.D ;
  wire \DFF_478.Q ;
  wire \DFF_479.CK ;
  wire \DFF_479.D ;
  wire \DFF_479.Q ;
  wire \DFF_48.CK ;
  wire \DFF_48.D ;
  wire \DFF_48.Q ;
  wire \DFF_480.CK ;
  wire \DFF_480.D ;
  wire \DFF_480.Q ;
  wire \DFF_481.CK ;
  wire \DFF_481.D ;
  wire \DFF_481.Q ;
  wire \DFF_482.CK ;
  wire \DFF_482.D ;
  wire \DFF_482.Q ;
  wire \DFF_483.CK ;
  wire \DFF_483.D ;
  wire \DFF_483.Q ;
  wire \DFF_484.CK ;
  wire \DFF_484.D ;
  wire \DFF_484.Q ;
  wire \DFF_485.CK ;
  wire \DFF_485.D ;
  wire \DFF_485.Q ;
  wire \DFF_486.CK ;
  wire \DFF_486.D ;
  wire \DFF_486.Q ;
  wire \DFF_487.CK ;
  wire \DFF_487.D ;
  wire \DFF_487.Q ;
  wire \DFF_488.CK ;
  wire \DFF_488.D ;
  wire \DFF_488.Q ;
  wire \DFF_489.CK ;
  wire \DFF_489.D ;
  wire \DFF_489.Q ;
  wire \DFF_49.CK ;
  wire \DFF_49.D ;
  wire \DFF_49.Q ;
  wire \DFF_490.CK ;
  wire \DFF_490.D ;
  wire \DFF_490.Q ;
  wire \DFF_491.CK ;
  wire \DFF_491.D ;
  wire \DFF_491.Q ;
  wire \DFF_492.CK ;
  wire \DFF_492.D ;
  wire \DFF_492.Q ;
  wire \DFF_493.CK ;
  wire \DFF_493.D ;
  wire \DFF_493.Q ;
  wire \DFF_494.CK ;
  wire \DFF_494.D ;
  wire \DFF_494.Q ;
  wire \DFF_495.CK ;
  wire \DFF_495.D ;
  wire \DFF_495.Q ;
  wire \DFF_496.CK ;
  wire \DFF_496.D ;
  wire \DFF_496.Q ;
  wire \DFF_497.CK ;
  wire \DFF_497.D ;
  wire \DFF_497.Q ;
  wire \DFF_498.CK ;
  wire \DFF_498.D ;
  wire \DFF_498.Q ;
  wire \DFF_499.CK ;
  wire \DFF_499.D ;
  wire \DFF_499.Q ;
  wire \DFF_5.CK ;
  wire \DFF_5.D ;
  wire \DFF_5.Q ;
  wire \DFF_50.CK ;
  wire \DFF_50.D ;
  wire \DFF_50.Q ;
  wire \DFF_500.CK ;
  wire \DFF_500.D ;
  wire \DFF_500.Q ;
  wire \DFF_501.CK ;
  wire \DFF_501.D ;
  wire \DFF_501.Q ;
  wire \DFF_502.CK ;
  wire \DFF_502.D ;
  wire \DFF_502.Q ;
  wire \DFF_503.CK ;
  wire \DFF_503.D ;
  wire \DFF_503.Q ;
  wire \DFF_504.CK ;
  wire \DFF_504.D ;
  wire \DFF_504.Q ;
  wire \DFF_505.CK ;
  wire \DFF_505.D ;
  wire \DFF_505.Q ;
  wire \DFF_506.CK ;
  wire \DFF_506.D ;
  wire \DFF_506.Q ;
  wire \DFF_507.CK ;
  wire \DFF_507.D ;
  wire \DFF_507.Q ;
  wire \DFF_508.CK ;
  wire \DFF_508.D ;
  wire \DFF_508.Q ;
  wire \DFF_509.CK ;
  wire \DFF_509.D ;
  wire \DFF_509.Q ;
  wire \DFF_51.CK ;
  wire \DFF_51.D ;
  wire \DFF_51.Q ;
  wire \DFF_510.CK ;
  wire \DFF_510.D ;
  wire \DFF_510.Q ;
  wire \DFF_511.CK ;
  wire \DFF_511.D ;
  wire \DFF_511.Q ;
  wire \DFF_512.CK ;
  wire \DFF_512.D ;
  wire \DFF_512.Q ;
  wire \DFF_513.CK ;
  wire \DFF_513.D ;
  wire \DFF_513.Q ;
  wire \DFF_514.CK ;
  wire \DFF_514.D ;
  wire \DFF_514.Q ;
  wire \DFF_515.CK ;
  wire \DFF_515.D ;
  wire \DFF_515.Q ;
  wire \DFF_516.CK ;
  wire \DFF_516.D ;
  wire \DFF_516.Q ;
  wire \DFF_517.CK ;
  wire \DFF_517.D ;
  wire \DFF_517.Q ;
  wire \DFF_518.CK ;
  wire \DFF_518.D ;
  wire \DFF_518.Q ;
  wire \DFF_519.CK ;
  wire \DFF_519.D ;
  wire \DFF_519.Q ;
  wire \DFF_52.CK ;
  wire \DFF_52.D ;
  wire \DFF_52.Q ;
  wire \DFF_520.CK ;
  wire \DFF_520.D ;
  wire \DFF_520.Q ;
  wire \DFF_521.CK ;
  wire \DFF_521.D ;
  wire \DFF_521.Q ;
  wire \DFF_522.CK ;
  wire \DFF_522.D ;
  wire \DFF_522.Q ;
  wire \DFF_523.CK ;
  wire \DFF_523.D ;
  wire \DFF_523.Q ;
  wire \DFF_524.CK ;
  wire \DFF_524.D ;
  wire \DFF_524.Q ;
  wire \DFF_525.CK ;
  wire \DFF_525.D ;
  wire \DFF_525.Q ;
  wire \DFF_526.CK ;
  wire \DFF_526.D ;
  wire \DFF_526.Q ;
  wire \DFF_527.CK ;
  wire \DFF_527.D ;
  wire \DFF_527.Q ;
  wire \DFF_528.CK ;
  wire \DFF_528.D ;
  wire \DFF_528.Q ;
  wire \DFF_529.CK ;
  wire \DFF_529.D ;
  wire \DFF_529.Q ;
  wire \DFF_53.CK ;
  wire \DFF_53.D ;
  wire \DFF_53.Q ;
  wire \DFF_530.CK ;
  wire \DFF_530.D ;
  wire \DFF_530.Q ;
  wire \DFF_531.CK ;
  wire \DFF_531.D ;
  wire \DFF_531.Q ;
  wire \DFF_532.CK ;
  wire \DFF_532.D ;
  wire \DFF_532.Q ;
  wire \DFF_533.CK ;
  wire \DFF_533.D ;
  wire \DFF_533.Q ;
  wire \DFF_534.CK ;
  wire \DFF_534.D ;
  wire \DFF_534.Q ;
  wire \DFF_535.CK ;
  wire \DFF_535.D ;
  wire \DFF_535.Q ;
  wire \DFF_536.CK ;
  wire \DFF_536.D ;
  wire \DFF_536.Q ;
  wire \DFF_537.CK ;
  wire \DFF_537.D ;
  wire \DFF_537.Q ;
  wire \DFF_538.CK ;
  wire \DFF_538.D ;
  wire \DFF_538.Q ;
  wire \DFF_539.CK ;
  wire \DFF_539.D ;
  wire \DFF_539.Q ;
  wire \DFF_54.CK ;
  wire \DFF_54.D ;
  wire \DFF_54.Q ;
  wire \DFF_540.CK ;
  wire \DFF_540.D ;
  wire \DFF_540.Q ;
  wire \DFF_541.CK ;
  wire \DFF_541.D ;
  wire \DFF_541.Q ;
  wire \DFF_542.CK ;
  wire \DFF_542.D ;
  wire \DFF_542.Q ;
  wire \DFF_543.CK ;
  wire \DFF_543.D ;
  wire \DFF_543.Q ;
  wire \DFF_544.CK ;
  wire \DFF_544.D ;
  wire \DFF_544.Q ;
  wire \DFF_545.CK ;
  wire \DFF_545.D ;
  wire \DFF_545.Q ;
  wire \DFF_546.CK ;
  wire \DFF_546.D ;
  wire \DFF_546.Q ;
  wire \DFF_547.CK ;
  wire \DFF_547.D ;
  wire \DFF_547.Q ;
  wire \DFF_548.CK ;
  wire \DFF_548.D ;
  wire \DFF_548.Q ;
  wire \DFF_549.CK ;
  wire \DFF_549.D ;
  wire \DFF_549.Q ;
  wire \DFF_55.CK ;
  wire \DFF_55.D ;
  wire \DFF_55.Q ;
  wire \DFF_550.CK ;
  wire \DFF_550.D ;
  wire \DFF_550.Q ;
  wire \DFF_551.CK ;
  wire \DFF_551.D ;
  wire \DFF_551.Q ;
  wire \DFF_552.CK ;
  wire \DFF_552.D ;
  wire \DFF_552.Q ;
  wire \DFF_553.CK ;
  wire \DFF_553.D ;
  wire \DFF_553.Q ;
  wire \DFF_554.CK ;
  wire \DFF_554.D ;
  wire \DFF_554.Q ;
  wire \DFF_555.CK ;
  wire \DFF_555.D ;
  wire \DFF_555.Q ;
  wire \DFF_556.CK ;
  wire \DFF_556.D ;
  wire \DFF_556.Q ;
  wire \DFF_557.CK ;
  wire \DFF_557.D ;
  wire \DFF_557.Q ;
  wire \DFF_558.CK ;
  wire \DFF_558.D ;
  wire \DFF_558.Q ;
  wire \DFF_559.CK ;
  wire \DFF_559.D ;
  wire \DFF_559.Q ;
  wire \DFF_56.CK ;
  wire \DFF_56.D ;
  wire \DFF_56.Q ;
  wire \DFF_560.CK ;
  wire \DFF_560.D ;
  wire \DFF_560.Q ;
  wire \DFF_561.CK ;
  wire \DFF_561.D ;
  wire \DFF_561.Q ;
  wire \DFF_562.CK ;
  wire \DFF_562.D ;
  wire \DFF_562.Q ;
  wire \DFF_563.CK ;
  wire \DFF_563.D ;
  wire \DFF_563.Q ;
  wire \DFF_564.CK ;
  wire \DFF_564.D ;
  wire \DFF_564.Q ;
  wire \DFF_565.CK ;
  wire \DFF_565.D ;
  wire \DFF_565.Q ;
  wire \DFF_566.CK ;
  wire \DFF_566.D ;
  wire \DFF_566.Q ;
  wire \DFF_567.CK ;
  wire \DFF_567.D ;
  wire \DFF_567.Q ;
  wire \DFF_568.CK ;
  wire \DFF_568.D ;
  wire \DFF_568.Q ;
  wire \DFF_569.CK ;
  wire \DFF_569.D ;
  wire \DFF_569.Q ;
  wire \DFF_57.CK ;
  wire \DFF_57.D ;
  wire \DFF_57.Q ;
  wire \DFF_570.CK ;
  wire \DFF_570.D ;
  wire \DFF_570.Q ;
  wire \DFF_571.CK ;
  wire \DFF_571.D ;
  wire \DFF_571.Q ;
  wire \DFF_572.CK ;
  wire \DFF_572.D ;
  wire \DFF_572.Q ;
  wire \DFF_573.CK ;
  wire \DFF_573.D ;
  wire \DFF_573.Q ;
  wire \DFF_574.CK ;
  wire \DFF_574.D ;
  wire \DFF_574.Q ;
  wire \DFF_575.CK ;
  wire \DFF_575.D ;
  wire \DFF_575.Q ;
  wire \DFF_576.CK ;
  wire \DFF_576.D ;
  wire \DFF_576.Q ;
  wire \DFF_577.CK ;
  wire \DFF_577.D ;
  wire \DFF_577.Q ;
  wire \DFF_578.CK ;
  wire \DFF_578.D ;
  wire \DFF_578.Q ;
  wire \DFF_579.CK ;
  wire \DFF_579.D ;
  wire \DFF_579.Q ;
  wire \DFF_58.CK ;
  wire \DFF_58.D ;
  wire \DFF_58.Q ;
  wire \DFF_580.CK ;
  wire \DFF_580.D ;
  wire \DFF_580.Q ;
  wire \DFF_581.CK ;
  wire \DFF_581.D ;
  wire \DFF_581.Q ;
  wire \DFF_582.CK ;
  wire \DFF_582.D ;
  wire \DFF_582.Q ;
  wire \DFF_583.CK ;
  wire \DFF_583.D ;
  wire \DFF_583.Q ;
  wire \DFF_584.CK ;
  wire \DFF_584.D ;
  wire \DFF_584.Q ;
  wire \DFF_585.CK ;
  wire \DFF_585.D ;
  wire \DFF_585.Q ;
  wire \DFF_586.CK ;
  wire \DFF_586.D ;
  wire \DFF_586.Q ;
  wire \DFF_587.CK ;
  wire \DFF_587.D ;
  wire \DFF_587.Q ;
  wire \DFF_588.CK ;
  wire \DFF_588.D ;
  wire \DFF_588.Q ;
  wire \DFF_589.CK ;
  wire \DFF_589.D ;
  wire \DFF_589.Q ;
  wire \DFF_59.CK ;
  wire \DFF_59.D ;
  wire \DFF_59.Q ;
  wire \DFF_590.CK ;
  wire \DFF_590.D ;
  wire \DFF_590.Q ;
  wire \DFF_591.CK ;
  wire \DFF_591.D ;
  wire \DFF_591.Q ;
  wire \DFF_592.CK ;
  wire \DFF_592.D ;
  wire \DFF_592.Q ;
  wire \DFF_593.CK ;
  wire \DFF_593.D ;
  wire \DFF_593.Q ;
  wire \DFF_594.CK ;
  wire \DFF_594.D ;
  wire \DFF_594.Q ;
  wire \DFF_595.CK ;
  wire \DFF_595.D ;
  wire \DFF_595.Q ;
  wire \DFF_596.CK ;
  wire \DFF_596.D ;
  wire \DFF_596.Q ;
  wire \DFF_597.CK ;
  wire \DFF_597.D ;
  wire \DFF_597.Q ;
  wire \DFF_598.CK ;
  wire \DFF_598.D ;
  wire \DFF_598.Q ;
  wire \DFF_599.CK ;
  wire \DFF_599.D ;
  wire \DFF_599.Q ;
  wire \DFF_6.CK ;
  wire \DFF_6.D ;
  wire \DFF_6.Q ;
  wire \DFF_60.CK ;
  wire \DFF_60.D ;
  wire \DFF_60.Q ;
  wire \DFF_600.CK ;
  wire \DFF_600.D ;
  wire \DFF_600.Q ;
  wire \DFF_601.CK ;
  wire \DFF_601.D ;
  wire \DFF_601.Q ;
  wire \DFF_602.CK ;
  wire \DFF_602.D ;
  wire \DFF_602.Q ;
  wire \DFF_603.CK ;
  wire \DFF_603.D ;
  wire \DFF_603.Q ;
  wire \DFF_604.CK ;
  wire \DFF_604.D ;
  wire \DFF_604.Q ;
  wire \DFF_605.CK ;
  wire \DFF_605.D ;
  wire \DFF_605.Q ;
  wire \DFF_606.CK ;
  wire \DFF_606.D ;
  wire \DFF_606.Q ;
  wire \DFF_607.CK ;
  wire \DFF_607.D ;
  wire \DFF_607.Q ;
  wire \DFF_608.CK ;
  wire \DFF_608.D ;
  wire \DFF_608.Q ;
  wire \DFF_609.CK ;
  wire \DFF_609.D ;
  wire \DFF_609.Q ;
  wire \DFF_61.CK ;
  wire \DFF_61.D ;
  wire \DFF_61.Q ;
  wire \DFF_610.CK ;
  wire \DFF_610.D ;
  wire \DFF_610.Q ;
  wire \DFF_611.CK ;
  wire \DFF_611.D ;
  wire \DFF_611.Q ;
  wire \DFF_612.CK ;
  wire \DFF_612.D ;
  wire \DFF_612.Q ;
  wire \DFF_613.CK ;
  wire \DFF_613.D ;
  wire \DFF_613.Q ;
  wire \DFF_614.CK ;
  wire \DFF_614.D ;
  wire \DFF_614.Q ;
  wire \DFF_615.CK ;
  wire \DFF_615.D ;
  wire \DFF_615.Q ;
  wire \DFF_616.CK ;
  wire \DFF_616.D ;
  wire \DFF_616.Q ;
  wire \DFF_617.CK ;
  wire \DFF_617.D ;
  wire \DFF_617.Q ;
  wire \DFF_618.CK ;
  wire \DFF_618.D ;
  wire \DFF_618.Q ;
  wire \DFF_619.CK ;
  wire \DFF_619.D ;
  wire \DFF_619.Q ;
  wire \DFF_62.CK ;
  wire \DFF_62.D ;
  wire \DFF_62.Q ;
  wire \DFF_620.CK ;
  wire \DFF_620.D ;
  wire \DFF_620.Q ;
  wire \DFF_621.CK ;
  wire \DFF_621.D ;
  wire \DFF_621.Q ;
  wire \DFF_622.CK ;
  wire \DFF_622.D ;
  wire \DFF_622.Q ;
  wire \DFF_623.CK ;
  wire \DFF_623.D ;
  wire \DFF_623.Q ;
  wire \DFF_624.CK ;
  wire \DFF_624.D ;
  wire \DFF_624.Q ;
  wire \DFF_625.CK ;
  wire \DFF_625.D ;
  wire \DFF_625.Q ;
  wire \DFF_626.CK ;
  wire \DFF_626.D ;
  wire \DFF_626.Q ;
  wire \DFF_627.CK ;
  wire \DFF_627.D ;
  wire \DFF_627.Q ;
  wire \DFF_628.CK ;
  wire \DFF_628.D ;
  wire \DFF_628.Q ;
  wire \DFF_629.CK ;
  wire \DFF_629.D ;
  wire \DFF_629.Q ;
  wire \DFF_63.CK ;
  wire \DFF_63.D ;
  wire \DFF_63.Q ;
  wire \DFF_630.CK ;
  wire \DFF_630.D ;
  wire \DFF_630.Q ;
  wire \DFF_631.CK ;
  wire \DFF_631.D ;
  wire \DFF_631.Q ;
  wire \DFF_632.CK ;
  wire \DFF_632.D ;
  wire \DFF_632.Q ;
  wire \DFF_633.CK ;
  wire \DFF_633.D ;
  wire \DFF_633.Q ;
  wire \DFF_634.CK ;
  wire \DFF_634.D ;
  wire \DFF_634.Q ;
  wire \DFF_635.CK ;
  wire \DFF_635.D ;
  wire \DFF_635.Q ;
  wire \DFF_636.CK ;
  wire \DFF_636.D ;
  wire \DFF_636.Q ;
  wire \DFF_637.CK ;
  wire \DFF_637.D ;
  wire \DFF_637.Q ;
  wire \DFF_638.CK ;
  wire \DFF_638.D ;
  wire \DFF_638.Q ;
  wire \DFF_639.CK ;
  wire \DFF_639.D ;
  wire \DFF_639.Q ;
  wire \DFF_64.CK ;
  wire \DFF_64.D ;
  wire \DFF_64.Q ;
  wire \DFF_640.CK ;
  wire \DFF_640.D ;
  wire \DFF_640.Q ;
  wire \DFF_641.CK ;
  wire \DFF_641.D ;
  wire \DFF_641.Q ;
  wire \DFF_642.CK ;
  wire \DFF_642.D ;
  wire \DFF_642.Q ;
  wire \DFF_643.CK ;
  wire \DFF_643.D ;
  wire \DFF_643.Q ;
  wire \DFF_644.CK ;
  wire \DFF_644.D ;
  wire \DFF_644.Q ;
  wire \DFF_645.CK ;
  wire \DFF_645.D ;
  wire \DFF_645.Q ;
  wire \DFF_646.CK ;
  wire \DFF_646.D ;
  wire \DFF_646.Q ;
  wire \DFF_647.CK ;
  wire \DFF_647.D ;
  wire \DFF_647.Q ;
  wire \DFF_648.CK ;
  wire \DFF_648.D ;
  wire \DFF_648.Q ;
  wire \DFF_649.CK ;
  wire \DFF_649.D ;
  wire \DFF_649.Q ;
  wire \DFF_65.CK ;
  wire \DFF_65.D ;
  wire \DFF_65.Q ;
  wire \DFF_650.CK ;
  wire \DFF_650.D ;
  wire \DFF_650.Q ;
  wire \DFF_651.CK ;
  wire \DFF_651.D ;
  wire \DFF_651.Q ;
  wire \DFF_652.CK ;
  wire \DFF_652.D ;
  wire \DFF_652.Q ;
  wire \DFF_653.CK ;
  wire \DFF_653.D ;
  wire \DFF_653.Q ;
  wire \DFF_654.CK ;
  wire \DFF_654.D ;
  wire \DFF_654.Q ;
  wire \DFF_655.CK ;
  wire \DFF_655.D ;
  wire \DFF_655.Q ;
  wire \DFF_656.CK ;
  wire \DFF_656.D ;
  wire \DFF_656.Q ;
  wire \DFF_657.CK ;
  wire \DFF_657.D ;
  wire \DFF_657.Q ;
  wire \DFF_658.CK ;
  wire \DFF_658.D ;
  wire \DFF_658.Q ;
  wire \DFF_659.CK ;
  wire \DFF_659.D ;
  wire \DFF_659.Q ;
  wire \DFF_66.CK ;
  wire \DFF_66.D ;
  wire \DFF_66.Q ;
  wire \DFF_660.CK ;
  wire \DFF_660.D ;
  wire \DFF_660.Q ;
  wire \DFF_661.CK ;
  wire \DFF_661.D ;
  wire \DFF_661.Q ;
  wire \DFF_662.CK ;
  wire \DFF_662.D ;
  wire \DFF_662.Q ;
  wire \DFF_663.CK ;
  wire \DFF_663.D ;
  wire \DFF_663.Q ;
  wire \DFF_664.CK ;
  wire \DFF_664.D ;
  wire \DFF_664.Q ;
  wire \DFF_665.CK ;
  wire \DFF_665.D ;
  wire \DFF_665.Q ;
  wire \DFF_666.CK ;
  wire \DFF_666.D ;
  wire \DFF_666.Q ;
  wire \DFF_667.CK ;
  wire \DFF_667.D ;
  wire \DFF_667.Q ;
  wire \DFF_668.CK ;
  wire \DFF_668.D ;
  wire \DFF_668.Q ;
  wire \DFF_669.CK ;
  wire \DFF_669.D ;
  wire \DFF_669.Q ;
  wire \DFF_67.CK ;
  wire \DFF_67.D ;
  wire \DFF_67.Q ;
  wire \DFF_670.CK ;
  wire \DFF_670.D ;
  wire \DFF_670.Q ;
  wire \DFF_671.CK ;
  wire \DFF_671.D ;
  wire \DFF_671.Q ;
  wire \DFF_672.CK ;
  wire \DFF_672.D ;
  wire \DFF_672.Q ;
  wire \DFF_673.CK ;
  wire \DFF_673.D ;
  wire \DFF_673.Q ;
  wire \DFF_674.CK ;
  wire \DFF_674.D ;
  wire \DFF_674.Q ;
  wire \DFF_675.CK ;
  wire \DFF_675.D ;
  wire \DFF_675.Q ;
  wire \DFF_676.CK ;
  wire \DFF_676.D ;
  wire \DFF_676.Q ;
  wire \DFF_677.CK ;
  wire \DFF_677.D ;
  wire \DFF_677.Q ;
  wire \DFF_678.CK ;
  wire \DFF_678.D ;
  wire \DFF_678.Q ;
  wire \DFF_679.CK ;
  wire \DFF_679.D ;
  wire \DFF_679.Q ;
  wire \DFF_68.CK ;
  wire \DFF_68.D ;
  wire \DFF_68.Q ;
  wire \DFF_680.CK ;
  wire \DFF_680.D ;
  wire \DFF_680.Q ;
  wire \DFF_681.CK ;
  wire \DFF_681.D ;
  wire \DFF_681.Q ;
  wire \DFF_682.CK ;
  wire \DFF_682.D ;
  wire \DFF_682.Q ;
  wire \DFF_683.CK ;
  wire \DFF_683.D ;
  wire \DFF_683.Q ;
  wire \DFF_684.CK ;
  wire \DFF_684.D ;
  wire \DFF_684.Q ;
  wire \DFF_685.CK ;
  wire \DFF_685.D ;
  wire \DFF_685.Q ;
  wire \DFF_686.CK ;
  wire \DFF_686.D ;
  wire \DFF_686.Q ;
  wire \DFF_687.CK ;
  wire \DFF_687.D ;
  wire \DFF_687.Q ;
  wire \DFF_688.CK ;
  wire \DFF_688.D ;
  wire \DFF_688.Q ;
  wire \DFF_689.CK ;
  wire \DFF_689.D ;
  wire \DFF_689.Q ;
  wire \DFF_69.CK ;
  wire \DFF_69.D ;
  wire \DFF_69.Q ;
  wire \DFF_690.CK ;
  wire \DFF_690.D ;
  wire \DFF_690.Q ;
  wire \DFF_691.CK ;
  wire \DFF_691.D ;
  wire \DFF_691.Q ;
  wire \DFF_692.CK ;
  wire \DFF_692.D ;
  wire \DFF_692.Q ;
  wire \DFF_693.CK ;
  wire \DFF_693.D ;
  wire \DFF_693.Q ;
  wire \DFF_694.CK ;
  wire \DFF_694.D ;
  wire \DFF_694.Q ;
  wire \DFF_695.CK ;
  wire \DFF_695.D ;
  wire \DFF_695.Q ;
  wire \DFF_696.CK ;
  wire \DFF_696.D ;
  wire \DFF_696.Q ;
  wire \DFF_697.CK ;
  wire \DFF_697.D ;
  wire \DFF_697.Q ;
  wire \DFF_698.CK ;
  wire \DFF_698.D ;
  wire \DFF_698.Q ;
  wire \DFF_699.CK ;
  wire \DFF_699.D ;
  wire \DFF_699.Q ;
  wire \DFF_7.CK ;
  wire \DFF_7.D ;
  wire \DFF_7.Q ;
  wire \DFF_70.CK ;
  wire \DFF_70.D ;
  wire \DFF_70.Q ;
  wire \DFF_700.CK ;
  wire \DFF_700.D ;
  wire \DFF_700.Q ;
  wire \DFF_701.CK ;
  wire \DFF_701.D ;
  wire \DFF_701.Q ;
  wire \DFF_702.CK ;
  wire \DFF_702.D ;
  wire \DFF_702.Q ;
  wire \DFF_703.CK ;
  wire \DFF_703.D ;
  wire \DFF_703.Q ;
  wire \DFF_704.CK ;
  wire \DFF_704.D ;
  wire \DFF_704.Q ;
  wire \DFF_705.CK ;
  wire \DFF_705.D ;
  wire \DFF_705.Q ;
  wire \DFF_706.CK ;
  wire \DFF_706.D ;
  wire \DFF_706.Q ;
  wire \DFF_707.CK ;
  wire \DFF_707.D ;
  wire \DFF_707.Q ;
  wire \DFF_708.CK ;
  wire \DFF_708.D ;
  wire \DFF_708.Q ;
  wire \DFF_709.CK ;
  wire \DFF_709.D ;
  wire \DFF_709.Q ;
  wire \DFF_71.CK ;
  wire \DFF_71.D ;
  wire \DFF_71.Q ;
  wire \DFF_710.CK ;
  wire \DFF_710.D ;
  wire \DFF_710.Q ;
  wire \DFF_711.CK ;
  wire \DFF_711.D ;
  wire \DFF_711.Q ;
  wire \DFF_712.CK ;
  wire \DFF_712.D ;
  wire \DFF_712.Q ;
  wire \DFF_713.CK ;
  wire \DFF_713.D ;
  wire \DFF_713.Q ;
  wire \DFF_714.CK ;
  wire \DFF_714.D ;
  wire \DFF_714.Q ;
  wire \DFF_715.CK ;
  wire \DFF_715.D ;
  wire \DFF_715.Q ;
  wire \DFF_716.CK ;
  wire \DFF_716.D ;
  wire \DFF_716.Q ;
  wire \DFF_717.CK ;
  wire \DFF_717.D ;
  wire \DFF_717.Q ;
  wire \DFF_718.CK ;
  wire \DFF_718.D ;
  wire \DFF_718.Q ;
  wire \DFF_719.CK ;
  wire \DFF_719.D ;
  wire \DFF_719.Q ;
  wire \DFF_72.CK ;
  wire \DFF_72.D ;
  wire \DFF_72.Q ;
  wire \DFF_720.CK ;
  wire \DFF_720.D ;
  wire \DFF_720.Q ;
  wire \DFF_721.CK ;
  wire \DFF_721.D ;
  wire \DFF_721.Q ;
  wire \DFF_722.CK ;
  wire \DFF_722.D ;
  wire \DFF_722.Q ;
  wire \DFF_723.CK ;
  wire \DFF_723.D ;
  wire \DFF_723.Q ;
  wire \DFF_724.CK ;
  wire \DFF_724.D ;
  wire \DFF_724.Q ;
  wire \DFF_725.CK ;
  wire \DFF_725.D ;
  wire \DFF_725.Q ;
  wire \DFF_726.CK ;
  wire \DFF_726.D ;
  wire \DFF_726.Q ;
  wire \DFF_727.CK ;
  wire \DFF_727.D ;
  wire \DFF_727.Q ;
  wire \DFF_728.CK ;
  wire \DFF_728.D ;
  wire \DFF_728.Q ;
  wire \DFF_729.CK ;
  wire \DFF_729.D ;
  wire \DFF_729.Q ;
  wire \DFF_73.CK ;
  wire \DFF_73.D ;
  wire \DFF_73.Q ;
  wire \DFF_730.CK ;
  wire \DFF_730.D ;
  wire \DFF_730.Q ;
  wire \DFF_731.CK ;
  wire \DFF_731.D ;
  wire \DFF_731.Q ;
  wire \DFF_732.CK ;
  wire \DFF_732.D ;
  wire \DFF_732.Q ;
  wire \DFF_733.CK ;
  wire \DFF_733.D ;
  wire \DFF_733.Q ;
  wire \DFF_734.CK ;
  wire \DFF_734.D ;
  wire \DFF_734.Q ;
  wire \DFF_735.CK ;
  wire \DFF_735.D ;
  wire \DFF_735.Q ;
  wire \DFF_736.CK ;
  wire \DFF_736.D ;
  wire \DFF_736.Q ;
  wire \DFF_737.CK ;
  wire \DFF_737.D ;
  wire \DFF_737.Q ;
  wire \DFF_738.CK ;
  wire \DFF_738.D ;
  wire \DFF_738.Q ;
  wire \DFF_739.CK ;
  wire \DFF_739.D ;
  wire \DFF_739.Q ;
  wire \DFF_74.CK ;
  wire \DFF_74.D ;
  wire \DFF_74.Q ;
  wire \DFF_740.CK ;
  wire \DFF_740.D ;
  wire \DFF_740.Q ;
  wire \DFF_741.CK ;
  wire \DFF_741.D ;
  wire \DFF_741.Q ;
  wire \DFF_742.CK ;
  wire \DFF_742.D ;
  wire \DFF_742.Q ;
  wire \DFF_743.CK ;
  wire \DFF_743.D ;
  wire \DFF_743.Q ;
  wire \DFF_744.CK ;
  wire \DFF_744.D ;
  wire \DFF_744.Q ;
  wire \DFF_745.CK ;
  wire \DFF_745.D ;
  wire \DFF_745.Q ;
  wire \DFF_746.CK ;
  wire \DFF_746.D ;
  wire \DFF_746.Q ;
  wire \DFF_747.CK ;
  wire \DFF_747.D ;
  wire \DFF_747.Q ;
  wire \DFF_748.CK ;
  wire \DFF_748.D ;
  wire \DFF_748.Q ;
  wire \DFF_749.CK ;
  wire \DFF_749.D ;
  wire \DFF_749.Q ;
  wire \DFF_75.CK ;
  wire \DFF_75.D ;
  wire \DFF_75.Q ;
  wire \DFF_750.CK ;
  wire \DFF_750.D ;
  wire \DFF_750.Q ;
  wire \DFF_751.CK ;
  wire \DFF_751.D ;
  wire \DFF_751.Q ;
  wire \DFF_752.CK ;
  wire \DFF_752.D ;
  wire \DFF_752.Q ;
  wire \DFF_753.CK ;
  wire \DFF_753.D ;
  wire \DFF_753.Q ;
  wire \DFF_754.CK ;
  wire \DFF_754.D ;
  wire \DFF_754.Q ;
  wire \DFF_755.CK ;
  wire \DFF_755.D ;
  wire \DFF_755.Q ;
  wire \DFF_756.CK ;
  wire \DFF_756.D ;
  wire \DFF_756.Q ;
  wire \DFF_757.CK ;
  wire \DFF_757.D ;
  wire \DFF_757.Q ;
  wire \DFF_758.CK ;
  wire \DFF_758.D ;
  wire \DFF_758.Q ;
  wire \DFF_759.CK ;
  wire \DFF_759.D ;
  wire \DFF_759.Q ;
  wire \DFF_76.CK ;
  wire \DFF_76.D ;
  wire \DFF_76.Q ;
  wire \DFF_760.CK ;
  wire \DFF_760.D ;
  wire \DFF_760.Q ;
  wire \DFF_761.CK ;
  wire \DFF_761.D ;
  wire \DFF_761.Q ;
  wire \DFF_762.CK ;
  wire \DFF_762.D ;
  wire \DFF_762.Q ;
  wire \DFF_763.CK ;
  wire \DFF_763.D ;
  wire \DFF_763.Q ;
  wire \DFF_764.CK ;
  wire \DFF_764.D ;
  wire \DFF_764.Q ;
  wire \DFF_765.CK ;
  wire \DFF_765.D ;
  wire \DFF_765.Q ;
  wire \DFF_766.CK ;
  wire \DFF_766.D ;
  wire \DFF_766.Q ;
  wire \DFF_767.CK ;
  wire \DFF_767.D ;
  wire \DFF_767.Q ;
  wire \DFF_768.CK ;
  wire \DFF_768.D ;
  wire \DFF_768.Q ;
  wire \DFF_769.CK ;
  wire \DFF_769.D ;
  wire \DFF_769.Q ;
  wire \DFF_77.CK ;
  wire \DFF_77.D ;
  wire \DFF_77.Q ;
  wire \DFF_770.CK ;
  wire \DFF_770.D ;
  wire \DFF_770.Q ;
  wire \DFF_771.CK ;
  wire \DFF_771.D ;
  wire \DFF_771.Q ;
  wire \DFF_772.CK ;
  wire \DFF_772.D ;
  wire \DFF_772.Q ;
  wire \DFF_773.CK ;
  wire \DFF_773.D ;
  wire \DFF_773.Q ;
  wire \DFF_774.CK ;
  wire \DFF_774.D ;
  wire \DFF_774.Q ;
  wire \DFF_775.CK ;
  wire \DFF_775.D ;
  wire \DFF_775.Q ;
  wire \DFF_776.CK ;
  wire \DFF_776.D ;
  wire \DFF_776.Q ;
  wire \DFF_777.CK ;
  wire \DFF_777.D ;
  wire \DFF_777.Q ;
  wire \DFF_778.CK ;
  wire \DFF_778.D ;
  wire \DFF_778.Q ;
  wire \DFF_779.CK ;
  wire \DFF_779.D ;
  wire \DFF_779.Q ;
  wire \DFF_78.CK ;
  wire \DFF_78.D ;
  wire \DFF_78.Q ;
  wire \DFF_780.CK ;
  wire \DFF_780.D ;
  wire \DFF_780.Q ;
  wire \DFF_781.CK ;
  wire \DFF_781.D ;
  wire \DFF_781.Q ;
  wire \DFF_782.CK ;
  wire \DFF_782.D ;
  wire \DFF_782.Q ;
  wire \DFF_783.CK ;
  wire \DFF_783.D ;
  wire \DFF_783.Q ;
  wire \DFF_784.CK ;
  wire \DFF_784.D ;
  wire \DFF_784.Q ;
  wire \DFF_785.CK ;
  wire \DFF_785.D ;
  wire \DFF_785.Q ;
  wire \DFF_786.CK ;
  wire \DFF_786.D ;
  wire \DFF_786.Q ;
  wire \DFF_787.CK ;
  wire \DFF_787.D ;
  wire \DFF_787.Q ;
  wire \DFF_788.CK ;
  wire \DFF_788.D ;
  wire \DFF_788.Q ;
  wire \DFF_789.CK ;
  wire \DFF_789.D ;
  wire \DFF_789.Q ;
  wire \DFF_79.CK ;
  wire \DFF_79.D ;
  wire \DFF_79.Q ;
  wire \DFF_790.CK ;
  wire \DFF_790.D ;
  wire \DFF_790.Q ;
  wire \DFF_791.CK ;
  wire \DFF_791.D ;
  wire \DFF_791.Q ;
  wire \DFF_792.CK ;
  wire \DFF_792.D ;
  wire \DFF_792.Q ;
  wire \DFF_793.CK ;
  wire \DFF_793.D ;
  wire \DFF_793.Q ;
  wire \DFF_794.CK ;
  wire \DFF_794.D ;
  wire \DFF_794.Q ;
  wire \DFF_795.CK ;
  wire \DFF_795.D ;
  wire \DFF_795.Q ;
  wire \DFF_796.CK ;
  wire \DFF_796.D ;
  wire \DFF_796.Q ;
  wire \DFF_797.CK ;
  wire \DFF_797.D ;
  wire \DFF_797.Q ;
  wire \DFF_798.CK ;
  wire \DFF_798.D ;
  wire \DFF_798.Q ;
  wire \DFF_799.CK ;
  wire \DFF_799.D ;
  wire \DFF_799.Q ;
  wire \DFF_8.CK ;
  wire \DFF_8.D ;
  wire \DFF_8.Q ;
  wire \DFF_80.CK ;
  wire \DFF_80.D ;
  wire \DFF_80.Q ;
  wire \DFF_800.CK ;
  wire \DFF_800.D ;
  wire \DFF_800.Q ;
  wire \DFF_801.CK ;
  wire \DFF_801.D ;
  wire \DFF_801.Q ;
  wire \DFF_802.CK ;
  wire \DFF_802.D ;
  wire \DFF_802.Q ;
  wire \DFF_803.CK ;
  wire \DFF_803.D ;
  wire \DFF_803.Q ;
  wire \DFF_804.CK ;
  wire \DFF_804.D ;
  wire \DFF_804.Q ;
  wire \DFF_805.CK ;
  wire \DFF_805.D ;
  wire \DFF_805.Q ;
  wire \DFF_806.CK ;
  wire \DFF_806.D ;
  wire \DFF_806.Q ;
  wire \DFF_807.CK ;
  wire \DFF_807.D ;
  wire \DFF_807.Q ;
  wire \DFF_808.CK ;
  wire \DFF_808.D ;
  wire \DFF_808.Q ;
  wire \DFF_809.CK ;
  wire \DFF_809.D ;
  wire \DFF_809.Q ;
  wire \DFF_81.CK ;
  wire \DFF_81.D ;
  wire \DFF_81.Q ;
  wire \DFF_810.CK ;
  wire \DFF_810.D ;
  wire \DFF_810.Q ;
  wire \DFF_811.CK ;
  wire \DFF_811.D ;
  wire \DFF_811.Q ;
  wire \DFF_812.CK ;
  wire \DFF_812.D ;
  wire \DFF_812.Q ;
  wire \DFF_813.CK ;
  wire \DFF_813.D ;
  wire \DFF_813.Q ;
  wire \DFF_814.CK ;
  wire \DFF_814.D ;
  wire \DFF_814.Q ;
  wire \DFF_815.CK ;
  wire \DFF_815.D ;
  wire \DFF_815.Q ;
  wire \DFF_816.CK ;
  wire \DFF_816.D ;
  wire \DFF_816.Q ;
  wire \DFF_817.CK ;
  wire \DFF_817.D ;
  wire \DFF_817.Q ;
  wire \DFF_818.CK ;
  wire \DFF_818.D ;
  wire \DFF_818.Q ;
  wire \DFF_819.CK ;
  wire \DFF_819.D ;
  wire \DFF_819.Q ;
  wire \DFF_82.CK ;
  wire \DFF_82.D ;
  wire \DFF_82.Q ;
  wire \DFF_820.CK ;
  wire \DFF_820.D ;
  wire \DFF_820.Q ;
  wire \DFF_821.CK ;
  wire \DFF_821.D ;
  wire \DFF_821.Q ;
  wire \DFF_822.CK ;
  wire \DFF_822.D ;
  wire \DFF_822.Q ;
  wire \DFF_823.CK ;
  wire \DFF_823.D ;
  wire \DFF_823.Q ;
  wire \DFF_824.CK ;
  wire \DFF_824.D ;
  wire \DFF_824.Q ;
  wire \DFF_825.CK ;
  wire \DFF_825.D ;
  wire \DFF_825.Q ;
  wire \DFF_826.CK ;
  wire \DFF_826.D ;
  wire \DFF_826.Q ;
  wire \DFF_827.CK ;
  wire \DFF_827.D ;
  wire \DFF_827.Q ;
  wire \DFF_828.CK ;
  wire \DFF_828.D ;
  wire \DFF_828.Q ;
  wire \DFF_829.CK ;
  wire \DFF_829.D ;
  wire \DFF_829.Q ;
  wire \DFF_83.CK ;
  wire \DFF_83.D ;
  wire \DFF_83.Q ;
  wire \DFF_830.CK ;
  wire \DFF_830.D ;
  wire \DFF_830.Q ;
  wire \DFF_831.CK ;
  wire \DFF_831.D ;
  wire \DFF_831.Q ;
  wire \DFF_832.CK ;
  wire \DFF_832.D ;
  wire \DFF_832.Q ;
  wire \DFF_833.CK ;
  wire \DFF_833.D ;
  wire \DFF_833.Q ;
  wire \DFF_834.CK ;
  wire \DFF_834.D ;
  wire \DFF_834.Q ;
  wire \DFF_835.CK ;
  wire \DFF_835.D ;
  wire \DFF_835.Q ;
  wire \DFF_836.CK ;
  wire \DFF_836.D ;
  wire \DFF_836.Q ;
  wire \DFF_837.CK ;
  wire \DFF_837.D ;
  wire \DFF_837.Q ;
  wire \DFF_838.CK ;
  wire \DFF_838.D ;
  wire \DFF_838.Q ;
  wire \DFF_839.CK ;
  wire \DFF_839.D ;
  wire \DFF_839.Q ;
  wire \DFF_84.CK ;
  wire \DFF_84.D ;
  wire \DFF_84.Q ;
  wire \DFF_840.CK ;
  wire \DFF_840.D ;
  wire \DFF_840.Q ;
  wire \DFF_841.CK ;
  wire \DFF_841.D ;
  wire \DFF_841.Q ;
  wire \DFF_842.CK ;
  wire \DFF_842.D ;
  wire \DFF_842.Q ;
  wire \DFF_843.CK ;
  wire \DFF_843.D ;
  wire \DFF_843.Q ;
  wire \DFF_844.CK ;
  wire \DFF_844.D ;
  wire \DFF_844.Q ;
  wire \DFF_845.CK ;
  wire \DFF_845.D ;
  wire \DFF_845.Q ;
  wire \DFF_846.CK ;
  wire \DFF_846.D ;
  wire \DFF_846.Q ;
  wire \DFF_847.CK ;
  wire \DFF_847.D ;
  wire \DFF_847.Q ;
  wire \DFF_848.CK ;
  wire \DFF_848.D ;
  wire \DFF_848.Q ;
  wire \DFF_849.CK ;
  wire \DFF_849.D ;
  wire \DFF_849.Q ;
  wire \DFF_85.CK ;
  wire \DFF_85.D ;
  wire \DFF_85.Q ;
  wire \DFF_850.CK ;
  wire \DFF_850.D ;
  wire \DFF_850.Q ;
  wire \DFF_851.CK ;
  wire \DFF_851.D ;
  wire \DFF_851.Q ;
  wire \DFF_852.CK ;
  wire \DFF_852.D ;
  wire \DFF_852.Q ;
  wire \DFF_853.CK ;
  wire \DFF_853.D ;
  wire \DFF_853.Q ;
  wire \DFF_854.CK ;
  wire \DFF_854.D ;
  wire \DFF_854.Q ;
  wire \DFF_855.CK ;
  wire \DFF_855.D ;
  wire \DFF_855.Q ;
  wire \DFF_856.CK ;
  wire \DFF_856.D ;
  wire \DFF_856.Q ;
  wire \DFF_857.CK ;
  wire \DFF_857.D ;
  wire \DFF_857.Q ;
  wire \DFF_858.CK ;
  wire \DFF_858.D ;
  wire \DFF_858.Q ;
  wire \DFF_859.CK ;
  wire \DFF_859.D ;
  wire \DFF_859.Q ;
  wire \DFF_86.CK ;
  wire \DFF_86.D ;
  wire \DFF_86.Q ;
  wire \DFF_860.CK ;
  wire \DFF_860.D ;
  wire \DFF_860.Q ;
  wire \DFF_861.CK ;
  wire \DFF_861.D ;
  wire \DFF_861.Q ;
  wire \DFF_862.CK ;
  wire \DFF_862.D ;
  wire \DFF_862.Q ;
  wire \DFF_863.CK ;
  wire \DFF_863.D ;
  wire \DFF_863.Q ;
  wire \DFF_864.CK ;
  wire \DFF_864.D ;
  wire \DFF_864.Q ;
  wire \DFF_865.CK ;
  wire \DFF_865.D ;
  wire \DFF_865.Q ;
  wire \DFF_866.CK ;
  wire \DFF_866.D ;
  wire \DFF_866.Q ;
  wire \DFF_867.CK ;
  wire \DFF_867.D ;
  wire \DFF_867.Q ;
  wire \DFF_868.CK ;
  wire \DFF_868.D ;
  wire \DFF_868.Q ;
  wire \DFF_869.CK ;
  wire \DFF_869.D ;
  wire \DFF_869.Q ;
  wire \DFF_87.CK ;
  wire \DFF_87.D ;
  wire \DFF_87.Q ;
  wire \DFF_870.CK ;
  wire \DFF_870.D ;
  wire \DFF_870.Q ;
  wire \DFF_871.CK ;
  wire \DFF_871.D ;
  wire \DFF_871.Q ;
  wire \DFF_872.CK ;
  wire \DFF_872.D ;
  wire \DFF_872.Q ;
  wire \DFF_873.CK ;
  wire \DFF_873.D ;
  wire \DFF_873.Q ;
  wire \DFF_874.CK ;
  wire \DFF_874.D ;
  wire \DFF_874.Q ;
  wire \DFF_875.CK ;
  wire \DFF_875.D ;
  wire \DFF_875.Q ;
  wire \DFF_876.CK ;
  wire \DFF_876.D ;
  wire \DFF_876.Q ;
  wire \DFF_877.CK ;
  wire \DFF_877.D ;
  wire \DFF_877.Q ;
  wire \DFF_878.CK ;
  wire \DFF_878.D ;
  wire \DFF_878.Q ;
  wire \DFF_879.CK ;
  wire \DFF_879.D ;
  wire \DFF_879.Q ;
  wire \DFF_88.CK ;
  wire \DFF_88.D ;
  wire \DFF_88.Q ;
  wire \DFF_880.CK ;
  wire \DFF_880.D ;
  wire \DFF_880.Q ;
  wire \DFF_881.CK ;
  wire \DFF_881.D ;
  wire \DFF_881.Q ;
  wire \DFF_882.CK ;
  wire \DFF_882.D ;
  wire \DFF_882.Q ;
  wire \DFF_883.CK ;
  wire \DFF_883.D ;
  wire \DFF_883.Q ;
  wire \DFF_884.CK ;
  wire \DFF_884.D ;
  wire \DFF_884.Q ;
  wire \DFF_885.CK ;
  wire \DFF_885.D ;
  wire \DFF_885.Q ;
  wire \DFF_886.CK ;
  wire \DFF_886.D ;
  wire \DFF_886.Q ;
  wire \DFF_887.CK ;
  wire \DFF_887.D ;
  wire \DFF_887.Q ;
  wire \DFF_888.CK ;
  wire \DFF_888.D ;
  wire \DFF_888.Q ;
  wire \DFF_889.CK ;
  wire \DFF_889.D ;
  wire \DFF_889.Q ;
  wire \DFF_89.CK ;
  wire \DFF_89.D ;
  wire \DFF_89.Q ;
  wire \DFF_890.CK ;
  wire \DFF_890.D ;
  wire \DFF_890.Q ;
  wire \DFF_891.CK ;
  wire \DFF_891.D ;
  wire \DFF_891.Q ;
  wire \DFF_892.CK ;
  wire \DFF_892.D ;
  wire \DFF_892.Q ;
  wire \DFF_893.CK ;
  wire \DFF_893.D ;
  wire \DFF_893.Q ;
  wire \DFF_894.CK ;
  wire \DFF_894.D ;
  wire \DFF_894.Q ;
  wire \DFF_895.CK ;
  wire \DFF_895.D ;
  wire \DFF_895.Q ;
  wire \DFF_896.CK ;
  wire \DFF_896.D ;
  wire \DFF_896.Q ;
  wire \DFF_897.CK ;
  wire \DFF_897.D ;
  wire \DFF_897.Q ;
  wire \DFF_898.CK ;
  wire \DFF_898.D ;
  wire \DFF_898.Q ;
  wire \DFF_899.CK ;
  wire \DFF_899.D ;
  wire \DFF_899.Q ;
  wire \DFF_9.CK ;
  wire \DFF_9.D ;
  wire \DFF_9.Q ;
  wire \DFF_90.CK ;
  wire \DFF_90.D ;
  wire \DFF_90.Q ;
  wire \DFF_900.CK ;
  wire \DFF_900.D ;
  wire \DFF_900.Q ;
  wire \DFF_901.CK ;
  wire \DFF_901.D ;
  wire \DFF_901.Q ;
  wire \DFF_902.CK ;
  wire \DFF_902.D ;
  wire \DFF_902.Q ;
  wire \DFF_903.CK ;
  wire \DFF_903.D ;
  wire \DFF_903.Q ;
  wire \DFF_904.CK ;
  wire \DFF_904.D ;
  wire \DFF_904.Q ;
  wire \DFF_905.CK ;
  wire \DFF_905.D ;
  wire \DFF_905.Q ;
  wire \DFF_906.CK ;
  wire \DFF_906.D ;
  wire \DFF_906.Q ;
  wire \DFF_907.CK ;
  wire \DFF_907.D ;
  wire \DFF_907.Q ;
  wire \DFF_908.CK ;
  wire \DFF_908.D ;
  wire \DFF_908.Q ;
  wire \DFF_909.CK ;
  wire \DFF_909.D ;
  wire \DFF_909.Q ;
  wire \DFF_91.CK ;
  wire \DFF_91.D ;
  wire \DFF_91.Q ;
  wire \DFF_910.CK ;
  wire \DFF_910.D ;
  wire \DFF_910.Q ;
  wire \DFF_911.CK ;
  wire \DFF_911.D ;
  wire \DFF_911.Q ;
  wire \DFF_912.CK ;
  wire \DFF_912.D ;
  wire \DFF_912.Q ;
  wire \DFF_913.CK ;
  wire \DFF_913.D ;
  wire \DFF_913.Q ;
  wire \DFF_914.CK ;
  wire \DFF_914.D ;
  wire \DFF_914.Q ;
  wire \DFF_915.CK ;
  wire \DFF_915.D ;
  wire \DFF_915.Q ;
  wire \DFF_916.CK ;
  wire \DFF_916.D ;
  wire \DFF_916.Q ;
  wire \DFF_917.CK ;
  wire \DFF_917.D ;
  wire \DFF_917.Q ;
  wire \DFF_918.CK ;
  wire \DFF_918.D ;
  wire \DFF_918.Q ;
  wire \DFF_919.CK ;
  wire \DFF_919.D ;
  wire \DFF_919.Q ;
  wire \DFF_92.CK ;
  wire \DFF_92.D ;
  wire \DFF_92.Q ;
  wire \DFF_920.CK ;
  wire \DFF_920.D ;
  wire \DFF_920.Q ;
  wire \DFF_921.CK ;
  wire \DFF_921.D ;
  wire \DFF_921.Q ;
  wire \DFF_922.CK ;
  wire \DFF_922.D ;
  wire \DFF_922.Q ;
  wire \DFF_923.CK ;
  wire \DFF_923.D ;
  wire \DFF_923.Q ;
  wire \DFF_924.CK ;
  wire \DFF_924.D ;
  wire \DFF_924.Q ;
  wire \DFF_925.CK ;
  wire \DFF_925.D ;
  wire \DFF_925.Q ;
  wire \DFF_926.CK ;
  wire \DFF_926.D ;
  wire \DFF_926.Q ;
  wire \DFF_927.CK ;
  wire \DFF_927.D ;
  wire \DFF_927.Q ;
  wire \DFF_928.CK ;
  wire \DFF_928.D ;
  wire \DFF_928.Q ;
  wire \DFF_929.CK ;
  wire \DFF_929.D ;
  wire \DFF_929.Q ;
  wire \DFF_93.CK ;
  wire \DFF_93.D ;
  wire \DFF_93.Q ;
  wire \DFF_930.CK ;
  wire \DFF_930.D ;
  wire \DFF_930.Q ;
  wire \DFF_931.CK ;
  wire \DFF_931.D ;
  wire \DFF_931.Q ;
  wire \DFF_932.CK ;
  wire \DFF_932.D ;
  wire \DFF_932.Q ;
  wire \DFF_933.CK ;
  wire \DFF_933.D ;
  wire \DFF_933.Q ;
  wire \DFF_934.CK ;
  wire \DFF_934.D ;
  wire \DFF_934.Q ;
  wire \DFF_935.CK ;
  wire \DFF_935.D ;
  wire \DFF_935.Q ;
  wire \DFF_936.CK ;
  wire \DFF_936.D ;
  wire \DFF_936.Q ;
  wire \DFF_937.CK ;
  wire \DFF_937.D ;
  wire \DFF_937.Q ;
  wire \DFF_938.CK ;
  wire \DFF_938.D ;
  wire \DFF_938.Q ;
  wire \DFF_939.CK ;
  wire \DFF_939.D ;
  wire \DFF_939.Q ;
  wire \DFF_94.CK ;
  wire \DFF_94.D ;
  wire \DFF_94.Q ;
  wire \DFF_940.CK ;
  wire \DFF_940.D ;
  wire \DFF_940.Q ;
  wire \DFF_941.CK ;
  wire \DFF_941.D ;
  wire \DFF_941.Q ;
  wire \DFF_942.CK ;
  wire \DFF_942.D ;
  wire \DFF_942.Q ;
  wire \DFF_943.CK ;
  wire \DFF_943.D ;
  wire \DFF_943.Q ;
  wire \DFF_944.CK ;
  wire \DFF_944.D ;
  wire \DFF_944.Q ;
  wire \DFF_945.CK ;
  wire \DFF_945.D ;
  wire \DFF_945.Q ;
  wire \DFF_946.CK ;
  wire \DFF_946.D ;
  wire \DFF_946.Q ;
  wire \DFF_947.CK ;
  wire \DFF_947.D ;
  wire \DFF_947.Q ;
  wire \DFF_948.CK ;
  wire \DFF_948.D ;
  wire \DFF_948.Q ;
  wire \DFF_949.CK ;
  wire \DFF_949.D ;
  wire \DFF_949.Q ;
  wire \DFF_95.CK ;
  wire \DFF_95.D ;
  wire \DFF_95.Q ;
  wire \DFF_950.CK ;
  wire \DFF_950.D ;
  wire \DFF_950.Q ;
  wire \DFF_951.CK ;
  wire \DFF_951.D ;
  wire \DFF_951.Q ;
  wire \DFF_952.CK ;
  wire \DFF_952.D ;
  wire \DFF_952.Q ;
  wire \DFF_953.CK ;
  wire \DFF_953.D ;
  wire \DFF_953.Q ;
  wire \DFF_954.CK ;
  wire \DFF_954.D ;
  wire \DFF_954.Q ;
  wire \DFF_955.CK ;
  wire \DFF_955.D ;
  wire \DFF_955.Q ;
  wire \DFF_956.CK ;
  wire \DFF_956.D ;
  wire \DFF_956.Q ;
  wire \DFF_957.CK ;
  wire \DFF_957.D ;
  wire \DFF_957.Q ;
  wire \DFF_958.CK ;
  wire \DFF_958.D ;
  wire \DFF_958.Q ;
  wire \DFF_959.CK ;
  wire \DFF_959.D ;
  wire \DFF_959.Q ;
  wire \DFF_96.CK ;
  wire \DFF_96.D ;
  wire \DFF_96.Q ;
  wire \DFF_960.CK ;
  wire \DFF_960.D ;
  wire \DFF_960.Q ;
  wire \DFF_961.CK ;
  wire \DFF_961.D ;
  wire \DFF_961.Q ;
  wire \DFF_962.CK ;
  wire \DFF_962.D ;
  wire \DFF_962.Q ;
  wire \DFF_963.CK ;
  wire \DFF_963.D ;
  wire \DFF_963.Q ;
  wire \DFF_964.CK ;
  wire \DFF_964.D ;
  wire \DFF_964.Q ;
  wire \DFF_965.CK ;
  wire \DFF_965.D ;
  wire \DFF_965.Q ;
  wire \DFF_966.CK ;
  wire \DFF_966.D ;
  wire \DFF_966.Q ;
  wire \DFF_967.CK ;
  wire \DFF_967.D ;
  wire \DFF_967.Q ;
  wire \DFF_968.CK ;
  wire \DFF_968.D ;
  wire \DFF_968.Q ;
  wire \DFF_969.CK ;
  wire \DFF_969.D ;
  wire \DFF_969.Q ;
  wire \DFF_97.CK ;
  wire \DFF_97.D ;
  wire \DFF_97.Q ;
  wire \DFF_970.CK ;
  wire \DFF_970.D ;
  wire \DFF_970.Q ;
  wire \DFF_971.CK ;
  wire \DFF_971.D ;
  wire \DFF_971.Q ;
  wire \DFF_972.CK ;
  wire \DFF_972.D ;
  wire \DFF_972.Q ;
  wire \DFF_973.CK ;
  wire \DFF_973.D ;
  wire \DFF_973.Q ;
  wire \DFF_974.CK ;
  wire \DFF_974.D ;
  wire \DFF_974.Q ;
  wire \DFF_975.CK ;
  wire \DFF_975.D ;
  wire \DFF_975.Q ;
  wire \DFF_976.CK ;
  wire \DFF_976.D ;
  wire \DFF_976.Q ;
  wire \DFF_977.CK ;
  wire \DFF_977.D ;
  wire \DFF_977.Q ;
  wire \DFF_978.CK ;
  wire \DFF_978.D ;
  wire \DFF_978.Q ;
  wire \DFF_979.CK ;
  wire \DFF_979.D ;
  wire \DFF_979.Q ;
  wire \DFF_98.CK ;
  wire \DFF_98.D ;
  wire \DFF_98.Q ;
  wire \DFF_980.CK ;
  wire \DFF_980.D ;
  wire \DFF_980.Q ;
  wire \DFF_981.CK ;
  wire \DFF_981.D ;
  wire \DFF_981.Q ;
  wire \DFF_982.CK ;
  wire \DFF_982.D ;
  wire \DFF_982.Q ;
  wire \DFF_983.CK ;
  wire \DFF_983.D ;
  wire \DFF_983.Q ;
  wire \DFF_984.CK ;
  wire \DFF_984.D ;
  wire \DFF_984.Q ;
  wire \DFF_985.CK ;
  wire \DFF_985.D ;
  wire \DFF_985.Q ;
  wire \DFF_986.CK ;
  wire \DFF_986.D ;
  wire \DFF_986.Q ;
  wire \DFF_987.CK ;
  wire \DFF_987.D ;
  wire \DFF_987.Q ;
  wire \DFF_988.CK ;
  wire \DFF_988.D ;
  wire \DFF_988.Q ;
  wire \DFF_989.CK ;
  wire \DFF_989.D ;
  wire \DFF_989.Q ;
  wire \DFF_99.CK ;
  wire \DFF_99.D ;
  wire \DFF_99.Q ;
  wire \DFF_990.CK ;
  wire \DFF_990.D ;
  wire \DFF_990.Q ;
  wire \DFF_991.CK ;
  wire \DFF_991.D ;
  wire \DFF_991.Q ;
  wire \DFF_992.CK ;
  wire \DFF_992.D ;
  wire \DFF_992.Q ;
  wire \DFF_993.CK ;
  wire \DFF_993.D ;
  wire \DFF_993.Q ;
  wire \DFF_994.CK ;
  wire \DFF_994.D ;
  wire \DFF_994.Q ;
  wire \DFF_995.CK ;
  wire \DFF_995.D ;
  wire \DFF_995.Q ;
  wire \DFF_996.CK ;
  wire \DFF_996.D ;
  wire \DFF_996.Q ;
  wire \DFF_997.CK ;
  wire \DFF_997.D ;
  wire \DFF_997.Q ;
  wire \DFF_998.CK ;
  wire \DFF_998.D ;
  wire \DFF_998.Q ;
  wire \DFF_999.CK ;
  wire \DFF_999.D ;
  wire \DFF_999.Q ;
  input GND;
  input RESET;
  input TM0;
  input TM1;
  input VDD;
  wire WX1001;
  wire WX1002;
  wire WX1003;
  wire WX1004;
  wire WX1005;
  wire WX10052;
  wire WX10053;
  wire WX10054;
  wire WX10055;
  wire WX10056;
  wire WX1010;
  wire WX1017;
  wire WX1024;
  wire WX1031;
  wire WX10314;
  wire WX10315;
  wire WX10317;
  wire WX10319;
  wire WX10321;
  wire WX10323;
  wire WX10325;
  wire WX10327;
  wire WX10329;
  wire WX10331;
  wire WX10333;
  wire WX10335;
  wire WX10337;
  wire WX10339;
  wire WX10341;
  wire WX10343;
  wire WX10345;
  wire WX10347;
  wire WX10349;
  wire WX10351;
  wire WX10353;
  wire WX10355;
  wire WX10357;
  wire WX10359;
  wire WX10361;
  wire WX10363;
  wire WX10365;
  wire WX10367;
  wire WX10369;
  wire WX10371;
  wire WX10373;
  wire WX10375;
  wire WX10377;
  wire WX1038;
  wire WX1045;
  wire WX1052;
  wire WX1059;
  wire WX1066;
  wire WX1073;
  wire WX1080;
  wire WX10828;
  wire WX10829;
  wire WX10830;
  wire WX10831;
  wire WX10832;
  wire WX10833;
  wire WX10834;
  wire WX10835;
  wire WX10836;
  wire WX10837;
  wire WX10838;
  wire WX10839;
  wire WX10840;
  wire WX10841;
  wire WX10842;
  wire WX10843;
  wire WX10844;
  wire WX10845;
  wire WX10846;
  wire WX10847;
  wire WX10848;
  wire WX10849;
  wire WX10850;
  wire WX10851;
  wire WX10852;
  wire WX10853;
  wire WX10854;
  wire WX10855;
  wire WX10856;
  wire WX10857;
  wire WX10858;
  wire WX10859;
  wire WX10860;
  wire WX10861;
  wire WX10862;
  wire WX10863;
  wire WX10864;
  wire WX10865;
  wire WX10866;
  wire WX10867;
  wire WX10868;
  wire WX10869;
  wire WX1087;
  wire WX10870;
  wire WX10871;
  wire WX10872;
  wire WX10873;
  wire WX10874;
  wire WX10875;
  wire WX10876;
  wire WX10877;
  wire WX10878;
  wire WX10879;
  wire WX10880;
  wire WX10881;
  wire WX10882;
  wire WX10883;
  wire WX10884;
  wire WX10885;
  wire WX10886;
  wire WX10887;
  wire WX10888;
  wire WX10889;
  wire WX10890;
  wire WX10891;
  wire WX1094;
  wire WX10988;
  wire WX10989;
  wire WX10990;
  wire WX10991;
  wire WX10992;
  wire WX10993;
  wire WX10994;
  wire WX10995;
  wire WX10996;
  wire WX10997;
  wire WX10998;
  wire WX10999;
  wire WX11000;
  wire WX11001;
  wire WX11002;
  wire WX11003;
  wire WX11004;
  wire WX11005;
  wire WX11006;
  wire WX11007;
  wire WX11008;
  wire WX11009;
  wire WX1101;
  wire WX11010;
  wire WX11011;
  wire WX11012;
  wire WX11013;
  wire WX11014;
  wire WX11015;
  wire WX11016;
  wire WX11017;
  wire WX11018;
  wire WX11019;
  wire WX11020;
  wire WX11021;
  wire WX11022;
  wire WX11023;
  wire WX11024;
  wire WX11025;
  wire WX11026;
  wire WX11027;
  wire WX11028;
  wire WX11029;
  wire WX11030;
  wire WX11031;
  wire WX11032;
  wire WX11033;
  wire WX11034;
  wire WX11035;
  wire WX11036;
  wire WX11037;
  wire WX11038;
  wire WX11039;
  wire WX11040;
  wire WX11041;
  wire WX11042;
  wire WX11043;
  wire WX11044;
  wire WX11045;
  wire WX11046;
  wire WX11047;
  wire WX11048;
  wire WX11049;
  wire WX11050;
  wire WX11051;
  wire WX11052;
  wire WX11053;
  wire WX11054;
  wire WX11055;
  wire WX11056;
  wire WX11057;
  wire WX11058;
  wire WX11059;
  wire WX11060;
  wire WX11061;
  wire WX11062;
  wire WX11063;
  wire WX11064;
  wire WX11065;
  wire WX11066;
  wire WX11067;
  wire WX11068;
  wire WX11069;
  wire WX11070;
  wire WX11071;
  wire WX11072;
  wire WX11073;
  wire WX11074;
  wire WX11075;
  wire WX11076;
  wire WX11077;
  wire WX11078;
  wire WX11079;
  wire WX1108;
  wire WX11080;
  wire WX11081;
  wire WX11082;
  wire WX11083;
  wire WX11084;
  wire WX11085;
  wire WX11086;
  wire WX11087;
  wire WX11088;
  wire WX11089;
  wire WX11090;
  wire WX11091;
  wire WX11092;
  wire WX11093;
  wire WX11094;
  wire WX11095;
  wire WX11096;
  wire WX11097;
  wire WX11098;
  wire WX11099;
  wire WX11100;
  wire WX11101;
  wire WX11102;
  wire WX11103;
  wire WX11104;
  wire WX11105;
  wire WX11106;
  wire WX11107;
  wire WX11108;
  wire WX11109;
  wire WX11110;
  wire WX11111;
  wire WX11112;
  wire WX11113;
  wire WX11114;
  wire WX11115;
  wire WX11116;
  wire WX11117;
  wire WX11118;
  wire WX11119;
  wire WX11120;
  wire WX11121;
  wire WX11122;
  wire WX11123;
  wire WX11124;
  wire WX11125;
  wire WX11126;
  wire WX11127;
  wire WX11128;
  wire WX11129;
  wire WX11130;
  wire WX11131;
  wire WX11132;
  wire WX11133;
  wire WX11134;
  wire WX11135;
  wire WX11136;
  wire WX11137;
  wire WX11138;
  wire WX11139;
  wire WX11140;
  wire WX11141;
  wire WX11142;
  wire WX11143;
  wire WX11144;
  wire WX11145;
  wire WX11146;
  wire WX11147;
  wire WX11148;
  wire WX11149;
  wire WX1115;
  wire WX11150;
  wire WX11151;
  wire WX11152;
  wire WX11153;
  wire WX11154;
  wire WX11155;
  wire WX11156;
  wire WX11157;
  wire WX11158;
  wire WX11159;
  wire WX11160;
  wire WX11161;
  wire WX11162;
  wire WX11163;
  wire WX11164;
  wire WX11165;
  wire WX11166;
  wire WX11167;
  wire WX11168;
  wire WX11169;
  wire WX11170;
  wire WX11171;
  wire WX11172;
  wire WX11173;
  wire WX11174;
  wire WX11175;
  wire WX11176;
  wire WX11177;
  wire WX11178;
  wire WX11179;
  wire WX11180;
  wire WX11181;
  wire WX11182;
  wire WX11183;
  wire WX11184;
  wire WX11185;
  wire WX11186;
  wire WX11187;
  wire WX11188;
  wire WX11189;
  wire WX11190;
  wire WX11191;
  wire WX11192;
  wire WX11193;
  wire WX11194;
  wire WX11195;
  wire WX11196;
  wire WX11197;
  wire WX11198;
  wire WX11199;
  wire WX11200;
  wire WX11201;
  wire WX11202;
  wire WX11203;
  wire WX11204;
  wire WX11205;
  wire WX11206;
  wire WX11207;
  wire WX11208;
  wire WX11209;
  wire WX11210;
  wire WX11211;
  wire WX11212;
  wire WX11213;
  wire WX11214;
  wire WX11215;
  wire WX11216;
  wire WX11217;
  wire WX11218;
  wire WX11219;
  wire WX1122;
  wire WX11220;
  wire WX11221;
  wire WX11222;
  wire WX11223;
  wire WX11224;
  wire WX11225;
  wire WX11226;
  wire WX11227;
  wire WX11228;
  wire WX11229;
  wire WX11230;
  wire WX11231;
  wire WX11232;
  wire WX11233;
  wire WX11234;
  wire WX11235;
  wire WX11236;
  wire WX11237;
  wire WX11238;
  wire WX11239;
  wire WX11240;
  wire WX11241;
  wire WX11242;
  wire WX11243;
  wire WX1129;
  wire WX11345;
  wire WX11346;
  wire WX11347;
  wire WX11348;
  wire WX11349;
  wire WX1136;
  wire WX1143;
  wire WX1150;
  wire WX1157;
  wire WX11607;
  wire WX11608;
  wire WX11610;
  wire WX11612;
  wire WX11614;
  wire WX11616;
  wire WX11618;
  wire WX11620;
  wire WX11622;
  wire WX11624;
  wire WX11626;
  wire WX11628;
  wire WX11630;
  wire WX11632;
  wire WX11634;
  wire WX11636;
  wire WX11638;
  wire WX1164;
  wire WX11640;
  wire WX11642;
  wire WX11644;
  wire WX11646;
  wire WX11648;
  wire WX11650;
  wire WX11652;
  wire WX11654;
  wire WX11656;
  wire WX11658;
  wire WX11660;
  wire WX11662;
  wire WX11664;
  wire WX11666;
  wire WX11668;
  wire WX11670;
  wire WX1171;
  wire WX1178;
  wire WX1185;
  wire WX1192;
  wire WX1199;
  wire WX1206;
  wire WX1213;
  wire WX1220;
  wire WX1227;
  wire WX1263;
  wire WX1264;
  wire WX1266;
  wire WX1268;
  wire WX1270;
  wire WX1272;
  wire WX1274;
  wire WX1276;
  wire WX1278;
  wire WX1280;
  wire WX1282;
  wire WX1284;
  wire WX1286;
  wire WX1288;
  wire WX1290;
  wire WX1292;
  wire WX1294;
  wire WX1296;
  wire WX1298;
  wire WX1300;
  wire WX1302;
  wire WX1304;
  wire WX1306;
  wire WX1308;
  wire WX1310;
  wire WX1312;
  wire WX1314;
  wire WX1316;
  wire WX1318;
  wire WX1320;
  wire WX1322;
  wire WX1324;
  wire WX1326;
  wire WX1777;
  wire WX1778;
  wire WX1779;
  wire WX1780;
  wire WX1781;
  wire WX1782;
  wire WX1783;
  wire WX1784;
  wire WX1785;
  wire WX1786;
  wire WX1787;
  wire WX1788;
  wire WX1789;
  wire WX1790;
  wire WX1791;
  wire WX1792;
  wire WX1793;
  wire WX1794;
  wire WX1795;
  wire WX1796;
  wire WX1797;
  wire WX1798;
  wire WX1799;
  wire WX1800;
  wire WX1801;
  wire WX1802;
  wire WX1803;
  wire WX1804;
  wire WX1805;
  wire WX1806;
  wire WX1807;
  wire WX1808;
  wire WX1809;
  wire WX1810;
  wire WX1811;
  wire WX1812;
  wire WX1813;
  wire WX1814;
  wire WX1815;
  wire WX1816;
  wire WX1817;
  wire WX1818;
  wire WX1819;
  wire WX1820;
  wire WX1821;
  wire WX1822;
  wire WX1823;
  wire WX1824;
  wire WX1825;
  wire WX1826;
  wire WX1827;
  wire WX1828;
  wire WX1829;
  wire WX1830;
  wire WX1831;
  wire WX1832;
  wire WX1833;
  wire WX1834;
  wire WX1835;
  wire WX1836;
  wire WX1837;
  wire WX1838;
  wire WX1839;
  wire WX1840;
  wire WX1937;
  wire WX1938;
  wire WX1939;
  wire WX1940;
  wire WX1941;
  wire WX1942;
  wire WX1943;
  wire WX1944;
  wire WX1945;
  wire WX1946;
  wire WX1947;
  wire WX1948;
  wire WX1949;
  wire WX1950;
  wire WX1951;
  wire WX1952;
  wire WX1953;
  wire WX1954;
  wire WX1955;
  wire WX1956;
  wire WX1957;
  wire WX1958;
  wire WX1959;
  wire WX1960;
  wire WX1961;
  wire WX1962;
  wire WX1963;
  wire WX1964;
  wire WX1965;
  wire WX1966;
  wire WX1967;
  wire WX1968;
  wire WX1969;
  wire WX1970;
  wire WX1971;
  wire WX1972;
  wire WX1973;
  wire WX1974;
  wire WX1975;
  wire WX1976;
  wire WX1977;
  wire WX1978;
  wire WX1979;
  wire WX1980;
  wire WX1981;
  wire WX1982;
  wire WX1983;
  wire WX1984;
  wire WX1985;
  wire WX1986;
  wire WX1987;
  wire WX1988;
  wire WX1989;
  wire WX1990;
  wire WX1991;
  wire WX1992;
  wire WX1993;
  wire WX1994;
  wire WX1995;
  wire WX1996;
  wire WX1997;
  wire WX1998;
  wire WX1999;
  wire WX2000;
  wire WX2001;
  wire WX2002;
  wire WX2003;
  wire WX2004;
  wire WX2005;
  wire WX2006;
  wire WX2007;
  wire WX2008;
  wire WX2009;
  wire WX2010;
  wire WX2011;
  wire WX2012;
  wire WX2013;
  wire WX2014;
  wire WX2015;
  wire WX2016;
  wire WX2017;
  wire WX2018;
  wire WX2019;
  wire WX2020;
  wire WX2021;
  wire WX2022;
  wire WX2023;
  wire WX2024;
  wire WX2025;
  wire WX2026;
  wire WX2027;
  wire WX2028;
  wire WX2029;
  wire WX2030;
  wire WX2031;
  wire WX2032;
  wire WX2033;
  wire WX2034;
  wire WX2035;
  wire WX2036;
  wire WX2037;
  wire WX2038;
  wire WX2039;
  wire WX2040;
  wire WX2041;
  wire WX2042;
  wire WX2043;
  wire WX2044;
  wire WX2045;
  wire WX2046;
  wire WX2047;
  wire WX2048;
  wire WX2049;
  wire WX2050;
  wire WX2051;
  wire WX2052;
  wire WX2053;
  wire WX2054;
  wire WX2055;
  wire WX2056;
  wire WX2057;
  wire WX2058;
  wire WX2059;
  wire WX2060;
  wire WX2061;
  wire WX2062;
  wire WX2063;
  wire WX2064;
  wire WX2065;
  wire WX2066;
  wire WX2067;
  wire WX2068;
  wire WX2069;
  wire WX2070;
  wire WX2071;
  wire WX2072;
  wire WX2073;
  wire WX2074;
  wire WX2075;
  wire WX2076;
  wire WX2077;
  wire WX2078;
  wire WX2079;
  wire WX2080;
  wire WX2081;
  wire WX2082;
  wire WX2083;
  wire WX2084;
  wire WX2085;
  wire WX2086;
  wire WX2087;
  wire WX2088;
  wire WX2089;
  wire WX2090;
  wire WX2091;
  wire WX2092;
  wire WX2093;
  wire WX2094;
  wire WX2095;
  wire WX2096;
  wire WX2097;
  wire WX2098;
  wire WX2099;
  wire WX2100;
  wire WX2101;
  wire WX2102;
  wire WX2103;
  wire WX2104;
  wire WX2105;
  wire WX2106;
  wire WX2107;
  wire WX2108;
  wire WX2109;
  wire WX2110;
  wire WX2111;
  wire WX2112;
  wire WX2113;
  wire WX2114;
  wire WX2115;
  wire WX2116;
  wire WX2117;
  wire WX2118;
  wire WX2119;
  wire WX2120;
  wire WX2121;
  wire WX2122;
  wire WX2123;
  wire WX2124;
  wire WX2125;
  wire WX2126;
  wire WX2127;
  wire WX2128;
  wire WX2129;
  wire WX2130;
  wire WX2131;
  wire WX2132;
  wire WX2133;
  wire WX2134;
  wire WX2135;
  wire WX2136;
  wire WX2137;
  wire WX2138;
  wire WX2139;
  wire WX2140;
  wire WX2141;
  wire WX2142;
  wire WX2143;
  wire WX2144;
  wire WX2145;
  wire WX2146;
  wire WX2147;
  wire WX2148;
  wire WX2149;
  wire WX2150;
  wire WX2151;
  wire WX2152;
  wire WX2153;
  wire WX2154;
  wire WX2155;
  wire WX2156;
  wire WX2157;
  wire WX2158;
  wire WX2159;
  wire WX2160;
  wire WX2161;
  wire WX2162;
  wire WX2163;
  wire WX2164;
  wire WX2165;
  wire WX2166;
  wire WX2167;
  wire WX2168;
  wire WX2169;
  wire WX2170;
  wire WX2171;
  wire WX2172;
  wire WX2173;
  wire WX2174;
  wire WX2175;
  wire WX2176;
  wire WX2177;
  wire WX2178;
  wire WX2179;
  wire WX2180;
  wire WX2181;
  wire WX2182;
  wire WX2183;
  wire WX2184;
  wire WX2185;
  wire WX2186;
  wire WX2187;
  wire WX2188;
  wire WX2189;
  wire WX2190;
  wire WX2191;
  wire WX2192;
  wire WX2294;
  wire WX2295;
  wire WX2296;
  wire WX2297;
  wire WX2298;
  wire WX2556;
  wire WX2557;
  wire WX2559;
  wire WX2561;
  wire WX2563;
  wire WX2565;
  wire WX2567;
  wire WX2569;
  wire WX2571;
  wire WX2573;
  wire WX2575;
  wire WX2577;
  wire WX2579;
  wire WX2581;
  wire WX2583;
  wire WX2585;
  wire WX2587;
  wire WX2589;
  wire WX2591;
  wire WX2593;
  wire WX2595;
  wire WX2597;
  wire WX2599;
  wire WX2601;
  wire WX2603;
  wire WX2605;
  wire WX2607;
  wire WX2609;
  wire WX2611;
  wire WX2613;
  wire WX2615;
  wire WX2617;
  wire WX2619;
  wire WX3070;
  wire WX3071;
  wire WX3072;
  wire WX3073;
  wire WX3074;
  wire WX3075;
  wire WX3076;
  wire WX3077;
  wire WX3078;
  wire WX3079;
  wire WX3080;
  wire WX3081;
  wire WX3082;
  wire WX3083;
  wire WX3084;
  wire WX3085;
  wire WX3086;
  wire WX3087;
  wire WX3088;
  wire WX3089;
  wire WX3090;
  wire WX3091;
  wire WX3092;
  wire WX3093;
  wire WX3094;
  wire WX3095;
  wire WX3096;
  wire WX3097;
  wire WX3098;
  wire WX3099;
  wire WX3100;
  wire WX3101;
  wire WX3102;
  wire WX3103;
  wire WX3104;
  wire WX3105;
  wire WX3106;
  wire WX3107;
  wire WX3108;
  wire WX3109;
  wire WX3110;
  wire WX3111;
  wire WX3112;
  wire WX3113;
  wire WX3114;
  wire WX3115;
  wire WX3116;
  wire WX3117;
  wire WX3118;
  wire WX3119;
  wire WX3120;
  wire WX3121;
  wire WX3122;
  wire WX3123;
  wire WX3124;
  wire WX3125;
  wire WX3126;
  wire WX3127;
  wire WX3128;
  wire WX3129;
  wire WX3130;
  wire WX3131;
  wire WX3132;
  wire WX3133;
  wire WX3230;
  wire WX3231;
  wire WX3232;
  wire WX3233;
  wire WX3234;
  wire WX3235;
  wire WX3236;
  wire WX3237;
  wire WX3238;
  wire WX3239;
  wire WX3240;
  wire WX3241;
  wire WX3242;
  wire WX3243;
  wire WX3244;
  wire WX3245;
  wire WX3246;
  wire WX3247;
  wire WX3248;
  wire WX3249;
  wire WX3250;
  wire WX3251;
  wire WX3252;
  wire WX3253;
  wire WX3254;
  wire WX3255;
  wire WX3256;
  wire WX3257;
  wire WX3258;
  wire WX3259;
  wire WX3260;
  wire WX3261;
  wire WX3262;
  wire WX3263;
  wire WX3264;
  wire WX3265;
  wire WX3266;
  wire WX3267;
  wire WX3268;
  wire WX3269;
  wire WX3270;
  wire WX3271;
  wire WX3272;
  wire WX3273;
  wire WX3274;
  wire WX3275;
  wire WX3276;
  wire WX3277;
  wire WX3278;
  wire WX3279;
  wire WX3280;
  wire WX3281;
  wire WX3282;
  wire WX3283;
  wire WX3284;
  wire WX3285;
  wire WX3286;
  wire WX3287;
  wire WX3288;
  wire WX3289;
  wire WX3290;
  wire WX3291;
  wire WX3292;
  wire WX3293;
  wire WX3294;
  wire WX3295;
  wire WX3296;
  wire WX3297;
  wire WX3298;
  wire WX3299;
  wire WX3300;
  wire WX3301;
  wire WX3302;
  wire WX3303;
  wire WX3304;
  wire WX3305;
  wire WX3306;
  wire WX3307;
  wire WX3308;
  wire WX3309;
  wire WX3310;
  wire WX3311;
  wire WX3312;
  wire WX3313;
  wire WX3314;
  wire WX3315;
  wire WX3316;
  wire WX3317;
  wire WX3318;
  wire WX3319;
  wire WX3320;
  wire WX3321;
  wire WX3322;
  wire WX3323;
  wire WX3324;
  wire WX3325;
  wire WX3326;
  wire WX3327;
  wire WX3328;
  wire WX3329;
  wire WX3330;
  wire WX3331;
  wire WX3332;
  wire WX3333;
  wire WX3334;
  wire WX3335;
  wire WX3336;
  wire WX3337;
  wire WX3338;
  wire WX3339;
  wire WX3340;
  wire WX3341;
  wire WX3342;
  wire WX3343;
  wire WX3344;
  wire WX3345;
  wire WX3346;
  wire WX3347;
  wire WX3348;
  wire WX3349;
  wire WX3350;
  wire WX3351;
  wire WX3352;
  wire WX3353;
  wire WX3354;
  wire WX3355;
  wire WX3356;
  wire WX3357;
  wire WX3358;
  wire WX3359;
  wire WX3360;
  wire WX3361;
  wire WX3362;
  wire WX3363;
  wire WX3364;
  wire WX3365;
  wire WX3366;
  wire WX3367;
  wire WX3368;
  wire WX3369;
  wire WX3370;
  wire WX3371;
  wire WX3372;
  wire WX3373;
  wire WX3374;
  wire WX3375;
  wire WX3376;
  wire WX3377;
  wire WX3378;
  wire WX3379;
  wire WX3380;
  wire WX3381;
  wire WX3382;
  wire WX3383;
  wire WX3384;
  wire WX3385;
  wire WX3386;
  wire WX3387;
  wire WX3388;
  wire WX3389;
  wire WX3390;
  wire WX3391;
  wire WX3392;
  wire WX3393;
  wire WX3394;
  wire WX3395;
  wire WX3396;
  wire WX3397;
  wire WX3398;
  wire WX3399;
  wire WX3400;
  wire WX3401;
  wire WX3402;
  wire WX3403;
  wire WX3404;
  wire WX3405;
  wire WX3406;
  wire WX3407;
  wire WX3408;
  wire WX3409;
  wire WX3410;
  wire WX3411;
  wire WX3412;
  wire WX3413;
  wire WX3414;
  wire WX3415;
  wire WX3416;
  wire WX3417;
  wire WX3418;
  wire WX3419;
  wire WX3420;
  wire WX3421;
  wire WX3422;
  wire WX3423;
  wire WX3424;
  wire WX3425;
  wire WX3426;
  wire WX3427;
  wire WX3428;
  wire WX3429;
  wire WX3430;
  wire WX3431;
  wire WX3432;
  wire WX3433;
  wire WX3434;
  wire WX3435;
  wire WX3436;
  wire WX3437;
  wire WX3438;
  wire WX3439;
  wire WX3440;
  wire WX3441;
  wire WX3442;
  wire WX3443;
  wire WX3444;
  wire WX3445;
  wire WX3446;
  wire WX3447;
  wire WX3448;
  wire WX3449;
  wire WX3450;
  wire WX3451;
  wire WX3452;
  wire WX3453;
  wire WX3454;
  wire WX3455;
  wire WX3456;
  wire WX3457;
  wire WX3458;
  wire WX3459;
  wire WX3460;
  wire WX3461;
  wire WX3462;
  wire WX3463;
  wire WX3464;
  wire WX3465;
  wire WX3466;
  wire WX3467;
  wire WX3468;
  wire WX3469;
  wire WX3470;
  wire WX3471;
  wire WX3472;
  wire WX3473;
  wire WX3474;
  wire WX3475;
  wire WX3476;
  wire WX3477;
  wire WX3478;
  wire WX3479;
  wire WX3480;
  wire WX3481;
  wire WX3482;
  wire WX3483;
  wire WX3484;
  wire WX3485;
  wire WX3587;
  wire WX3588;
  wire WX3589;
  wire WX3590;
  wire WX3591;
  wire WX3849;
  wire WX3850;
  wire WX3852;
  wire WX3854;
  wire WX3856;
  wire WX3858;
  wire WX3860;
  wire WX3862;
  wire WX3864;
  wire WX3866;
  wire WX3868;
  wire WX3870;
  wire WX3872;
  wire WX3874;
  wire WX3876;
  wire WX3878;
  wire WX3880;
  wire WX3882;
  wire WX3884;
  wire WX3886;
  wire WX3888;
  wire WX3890;
  wire WX3892;
  wire WX3894;
  wire WX3896;
  wire WX3898;
  wire WX3900;
  wire WX3902;
  wire WX3904;
  wire WX3906;
  wire WX3908;
  wire WX3910;
  wire WX3912;
  wire WX4363;
  wire WX4364;
  wire WX4365;
  wire WX4366;
  wire WX4367;
  wire WX4368;
  wire WX4369;
  wire WX4370;
  wire WX4371;
  wire WX4372;
  wire WX4373;
  wire WX4374;
  wire WX4375;
  wire WX4376;
  wire WX4377;
  wire WX4378;
  wire WX4379;
  wire WX4380;
  wire WX4381;
  wire WX4382;
  wire WX4383;
  wire WX4384;
  wire WX4385;
  wire WX4386;
  wire WX4387;
  wire WX4388;
  wire WX4389;
  wire WX4390;
  wire WX4391;
  wire WX4392;
  wire WX4393;
  wire WX4394;
  wire WX4395;
  wire WX4396;
  wire WX4397;
  wire WX4398;
  wire WX4399;
  wire WX4400;
  wire WX4401;
  wire WX4402;
  wire WX4403;
  wire WX4404;
  wire WX4405;
  wire WX4406;
  wire WX4407;
  wire WX4408;
  wire WX4409;
  wire WX4410;
  wire WX4411;
  wire WX4412;
  wire WX4413;
  wire WX4414;
  wire WX4415;
  wire WX4416;
  wire WX4417;
  wire WX4418;
  wire WX4419;
  wire WX4420;
  wire WX4421;
  wire WX4422;
  wire WX4423;
  wire WX4424;
  wire WX4425;
  wire WX4426;
  wire WX4523;
  wire WX4524;
  wire WX4525;
  wire WX4526;
  wire WX4527;
  wire WX4528;
  wire WX4529;
  wire WX4530;
  wire WX4531;
  wire WX4532;
  wire WX4533;
  wire WX4534;
  wire WX4535;
  wire WX4536;
  wire WX4537;
  wire WX4538;
  wire WX4539;
  wire WX4540;
  wire WX4541;
  wire WX4542;
  wire WX4543;
  wire WX4544;
  wire WX4545;
  wire WX4546;
  wire WX4547;
  wire WX4548;
  wire WX4549;
  wire WX4550;
  wire WX4551;
  wire WX4552;
  wire WX4553;
  wire WX4554;
  wire WX4555;
  wire WX4556;
  wire WX4557;
  wire WX4558;
  wire WX4559;
  wire WX4560;
  wire WX4561;
  wire WX4562;
  wire WX4563;
  wire WX4564;
  wire WX4565;
  wire WX4566;
  wire WX4567;
  wire WX4568;
  wire WX4569;
  wire WX4570;
  wire WX4571;
  wire WX4572;
  wire WX4573;
  wire WX4574;
  wire WX4575;
  wire WX4576;
  wire WX4577;
  wire WX4578;
  wire WX4579;
  wire WX4580;
  wire WX4581;
  wire WX4582;
  wire WX4583;
  wire WX4584;
  wire WX4585;
  wire WX4586;
  wire WX4587;
  wire WX4588;
  wire WX4589;
  wire WX4590;
  wire WX4591;
  wire WX4592;
  wire WX4593;
  wire WX4594;
  wire WX4595;
  wire WX4596;
  wire WX4597;
  wire WX4598;
  wire WX4599;
  wire WX4600;
  wire WX4601;
  wire WX4602;
  wire WX4603;
  wire WX4604;
  wire WX4605;
  wire WX4606;
  wire WX4607;
  wire WX4608;
  wire WX4609;
  wire WX4610;
  wire WX4611;
  wire WX4612;
  wire WX4613;
  wire WX4614;
  wire WX4615;
  wire WX4616;
  wire WX4617;
  wire WX4618;
  wire WX4619;
  wire WX4620;
  wire WX4621;
  wire WX4622;
  wire WX4623;
  wire WX4624;
  wire WX4625;
  wire WX4626;
  wire WX4627;
  wire WX4628;
  wire WX4629;
  wire WX4630;
  wire WX4631;
  wire WX4632;
  wire WX4633;
  wire WX4634;
  wire WX4635;
  wire WX4636;
  wire WX4637;
  wire WX4638;
  wire WX4639;
  wire WX4640;
  wire WX4641;
  wire WX4642;
  wire WX4643;
  wire WX4644;
  wire WX4645;
  wire WX4646;
  wire WX4647;
  wire WX4648;
  wire WX4649;
  wire WX4650;
  wire WX4651;
  wire WX4652;
  wire WX4653;
  wire WX4654;
  wire WX4655;
  wire WX4656;
  wire WX4657;
  wire WX4658;
  wire WX4659;
  wire WX4660;
  wire WX4661;
  wire WX4662;
  wire WX4663;
  wire WX4664;
  wire WX4665;
  wire WX4666;
  wire WX4667;
  wire WX4668;
  wire WX4669;
  wire WX4670;
  wire WX4671;
  wire WX4672;
  wire WX4673;
  wire WX4674;
  wire WX4675;
  wire WX4676;
  wire WX4677;
  wire WX4678;
  wire WX4679;
  wire WX4680;
  wire WX4681;
  wire WX4682;
  wire WX4683;
  wire WX4684;
  wire WX4685;
  wire WX4686;
  wire WX4687;
  wire WX4688;
  wire WX4689;
  wire WX4690;
  wire WX4691;
  wire WX4692;
  wire WX4693;
  wire WX4694;
  wire WX4695;
  wire WX4696;
  wire WX4697;
  wire WX4698;
  wire WX4699;
  wire WX4700;
  wire WX4701;
  wire WX4702;
  wire WX4703;
  wire WX4704;
  wire WX4705;
  wire WX4706;
  wire WX4707;
  wire WX4708;
  wire WX4709;
  wire WX4710;
  wire WX4711;
  wire WX4712;
  wire WX4713;
  wire WX4714;
  wire WX4715;
  wire WX4716;
  wire WX4717;
  wire WX4718;
  wire WX4719;
  wire WX4720;
  wire WX4721;
  wire WX4722;
  wire WX4723;
  wire WX4724;
  wire WX4725;
  wire WX4726;
  wire WX4727;
  wire WX4728;
  wire WX4729;
  wire WX4730;
  wire WX4731;
  wire WX4732;
  wire WX4733;
  wire WX4734;
  wire WX4735;
  wire WX4736;
  wire WX4737;
  wire WX4738;
  wire WX4739;
  wire WX4740;
  wire WX4741;
  wire WX4742;
  wire WX4743;
  wire WX4744;
  wire WX4745;
  wire WX4746;
  wire WX4747;
  wire WX4748;
  wire WX4749;
  wire WX4750;
  wire WX4751;
  wire WX4752;
  wire WX4753;
  wire WX4754;
  wire WX4755;
  wire WX4756;
  wire WX4757;
  wire WX4758;
  wire WX4759;
  wire WX4760;
  wire WX4761;
  wire WX4762;
  wire WX4763;
  wire WX4764;
  wire WX4765;
  wire WX4766;
  wire WX4767;
  wire WX4768;
  wire WX4769;
  wire WX4770;
  wire WX4771;
  wire WX4772;
  wire WX4773;
  wire WX4774;
  wire WX4775;
  wire WX4776;
  wire WX4777;
  wire WX4778;
  wire WX484;
  wire WX485;
  wire WX486;
  wire WX487;
  wire WX488;
  wire WX4880;
  wire WX4881;
  wire WX4882;
  wire WX4883;
  wire WX4884;
  wire WX489;
  wire WX490;
  wire WX491;
  wire WX492;
  wire WX493;
  wire WX494;
  wire WX495;
  wire WX496;
  wire WX497;
  wire WX498;
  wire WX499;
  wire WX500;
  wire WX501;
  wire WX502;
  wire WX503;
  wire WX504;
  wire WX505;
  wire WX506;
  wire WX507;
  wire WX508;
  wire WX509;
  wire WX510;
  wire WX511;
  wire WX512;
  wire WX513;
  wire WX514;
  wire WX5142;
  wire WX5143;
  wire WX5145;
  wire WX5147;
  wire WX5149;
  wire WX515;
  wire WX5151;
  wire WX5153;
  wire WX5155;
  wire WX5157;
  wire WX5159;
  wire WX516;
  wire WX5161;
  wire WX5163;
  wire WX5165;
  wire WX5167;
  wire WX5169;
  wire WX517;
  wire WX5171;
  wire WX5173;
  wire WX5175;
  wire WX5177;
  wire WX5179;
  wire WX518;
  wire WX5181;
  wire WX5183;
  wire WX5185;
  wire WX5187;
  wire WX5189;
  wire WX519;
  wire WX5191;
  wire WX5193;
  wire WX5195;
  wire WX5197;
  wire WX5199;
  wire WX520;
  wire WX5201;
  wire WX5203;
  wire WX5205;
  wire WX521;
  wire WX522;
  wire WX523;
  wire WX524;
  wire WX525;
  wire WX526;
  wire WX527;
  wire WX528;
  wire WX529;
  wire WX530;
  wire WX531;
  wire WX532;
  wire WX533;
  wire WX534;
  wire WX535;
  wire WX536;
  wire WX537;
  wire WX538;
  wire WX539;
  wire WX540;
  wire WX541;
  wire WX542;
  wire WX543;
  wire WX544;
  wire WX545;
  wire WX546;
  wire WX547;
  wire WX5656;
  wire WX5657;
  wire WX5658;
  wire WX5659;
  wire WX5660;
  wire WX5661;
  wire WX5662;
  wire WX5663;
  wire WX5664;
  wire WX5665;
  wire WX5666;
  wire WX5667;
  wire WX5668;
  wire WX5669;
  wire WX5670;
  wire WX5671;
  wire WX5672;
  wire WX5673;
  wire WX5674;
  wire WX5675;
  wire WX5676;
  wire WX5677;
  wire WX5678;
  wire WX5679;
  wire WX5680;
  wire WX5681;
  wire WX5682;
  wire WX5683;
  wire WX5684;
  wire WX5685;
  wire WX5686;
  wire WX5687;
  wire WX5688;
  wire WX5689;
  wire WX5690;
  wire WX5691;
  wire WX5692;
  wire WX5693;
  wire WX5694;
  wire WX5695;
  wire WX5696;
  wire WX5697;
  wire WX5698;
  wire WX5699;
  wire WX5700;
  wire WX5701;
  wire WX5702;
  wire WX5703;
  wire WX5704;
  wire WX5705;
  wire WX5706;
  wire WX5707;
  wire WX5708;
  wire WX5709;
  wire WX5710;
  wire WX5711;
  wire WX5712;
  wire WX5713;
  wire WX5714;
  wire WX5715;
  wire WX5716;
  wire WX5717;
  wire WX5718;
  wire WX5719;
  wire WX5816;
  wire WX5817;
  wire WX5818;
  wire WX5819;
  wire WX5820;
  wire WX5821;
  wire WX5822;
  wire WX5823;
  wire WX5824;
  wire WX5825;
  wire WX5826;
  wire WX5827;
  wire WX5828;
  wire WX5829;
  wire WX5830;
  wire WX5831;
  wire WX5832;
  wire WX5833;
  wire WX5834;
  wire WX5835;
  wire WX5836;
  wire WX5837;
  wire WX5838;
  wire WX5839;
  wire WX5840;
  wire WX5841;
  wire WX5842;
  wire WX5843;
  wire WX5844;
  wire WX5845;
  wire WX5846;
  wire WX5847;
  wire WX5848;
  wire WX5849;
  wire WX5850;
  wire WX5851;
  wire WX5852;
  wire WX5853;
  wire WX5854;
  wire WX5855;
  wire WX5856;
  wire WX5857;
  wire WX5858;
  wire WX5859;
  wire WX5860;
  wire WX5861;
  wire WX5862;
  wire WX5863;
  wire WX5864;
  wire WX5865;
  wire WX5866;
  wire WX5867;
  wire WX5868;
  wire WX5869;
  wire WX5870;
  wire WX5871;
  wire WX5872;
  wire WX5873;
  wire WX5874;
  wire WX5875;
  wire WX5876;
  wire WX5877;
  wire WX5878;
  wire WX5879;
  wire WX5880;
  wire WX5881;
  wire WX5882;
  wire WX5883;
  wire WX5884;
  wire WX5885;
  wire WX5886;
  wire WX5887;
  wire WX5888;
  wire WX5889;
  wire WX5890;
  wire WX5891;
  wire WX5892;
  wire WX5893;
  wire WX5894;
  wire WX5895;
  wire WX5896;
  wire WX5897;
  wire WX5898;
  wire WX5899;
  wire WX5900;
  wire WX5901;
  wire WX5902;
  wire WX5903;
  wire WX5904;
  wire WX5905;
  wire WX5906;
  wire WX5907;
  wire WX5908;
  wire WX5909;
  wire WX5910;
  wire WX5911;
  wire WX5912;
  wire WX5913;
  wire WX5914;
  wire WX5915;
  wire WX5916;
  wire WX5917;
  wire WX5918;
  wire WX5919;
  wire WX5920;
  wire WX5921;
  wire WX5922;
  wire WX5923;
  wire WX5924;
  wire WX5925;
  wire WX5926;
  wire WX5927;
  wire WX5928;
  wire WX5929;
  wire WX5930;
  wire WX5931;
  wire WX5932;
  wire WX5933;
  wire WX5934;
  wire WX5935;
  wire WX5936;
  wire WX5937;
  wire WX5938;
  wire WX5939;
  wire WX5940;
  wire WX5941;
  wire WX5942;
  wire WX5943;
  wire WX5944;
  wire WX5945;
  wire WX5946;
  wire WX5947;
  wire WX5948;
  wire WX5949;
  wire WX5950;
  wire WX5951;
  wire WX5952;
  wire WX5953;
  wire WX5954;
  wire WX5955;
  wire WX5956;
  wire WX5957;
  wire WX5958;
  wire WX5959;
  wire WX5960;
  wire WX5961;
  wire WX5962;
  wire WX5963;
  wire WX5964;
  wire WX5965;
  wire WX5966;
  wire WX5967;
  wire WX5968;
  wire WX5969;
  wire WX5970;
  wire WX5971;
  wire WX5972;
  wire WX5973;
  wire WX5974;
  wire WX5975;
  wire WX5976;
  wire WX5977;
  wire WX5978;
  wire WX5979;
  wire WX5980;
  wire WX5981;
  wire WX5982;
  wire WX5983;
  wire WX5984;
  wire WX5985;
  wire WX5986;
  wire WX5987;
  wire WX5988;
  wire WX5989;
  wire WX5990;
  wire WX5991;
  wire WX5992;
  wire WX5993;
  wire WX5994;
  wire WX5995;
  wire WX5996;
  wire WX5997;
  wire WX5998;
  wire WX5999;
  wire WX6000;
  wire WX6001;
  wire WX6002;
  wire WX6003;
  wire WX6004;
  wire WX6005;
  wire WX6006;
  wire WX6007;
  wire WX6008;
  wire WX6009;
  wire WX6010;
  wire WX6011;
  wire WX6012;
  wire WX6013;
  wire WX6014;
  wire WX6015;
  wire WX6016;
  wire WX6017;
  wire WX6018;
  wire WX6019;
  wire WX6020;
  wire WX6021;
  wire WX6022;
  wire WX6023;
  wire WX6024;
  wire WX6025;
  wire WX6026;
  wire WX6027;
  wire WX6028;
  wire WX6029;
  wire WX6030;
  wire WX6031;
  wire WX6032;
  wire WX6033;
  wire WX6034;
  wire WX6035;
  wire WX6036;
  wire WX6037;
  wire WX6038;
  wire WX6039;
  wire WX6040;
  wire WX6041;
  wire WX6042;
  wire WX6043;
  wire WX6044;
  wire WX6045;
  wire WX6046;
  wire WX6047;
  wire WX6048;
  wire WX6049;
  wire WX6050;
  wire WX6051;
  wire WX6052;
  wire WX6053;
  wire WX6054;
  wire WX6055;
  wire WX6056;
  wire WX6057;
  wire WX6058;
  wire WX6059;
  wire WX6060;
  wire WX6061;
  wire WX6062;
  wire WX6063;
  wire WX6064;
  wire WX6065;
  wire WX6066;
  wire WX6067;
  wire WX6068;
  wire WX6069;
  wire WX6070;
  wire WX6071;
  wire WX6173;
  wire WX6174;
  wire WX6175;
  wire WX6176;
  wire WX6177;
  wire WX6435;
  wire WX6436;
  wire WX6438;
  wire WX644;
  wire WX6440;
  wire WX6442;
  wire WX6444;
  wire WX6446;
  wire WX6448;
  wire WX645;
  wire WX6450;
  wire WX6452;
  wire WX6454;
  wire WX6456;
  wire WX6458;
  wire WX646;
  wire WX6460;
  wire WX6462;
  wire WX6464;
  wire WX6466;
  wire WX6468;
  wire WX647;
  wire WX6470;
  wire WX6472;
  wire WX6474;
  wire WX6476;
  wire WX6478;
  wire WX648;
  wire WX6480;
  wire WX6482;
  wire WX6484;
  wire WX6486;
  wire WX6488;
  wire WX649;
  wire WX6490;
  wire WX6492;
  wire WX6494;
  wire WX6496;
  wire WX6498;
  wire WX650;
  wire WX651;
  wire WX652;
  wire WX653;
  wire WX654;
  wire WX655;
  wire WX656;
  wire WX657;
  wire WX658;
  wire WX659;
  wire WX660;
  wire WX661;
  wire WX662;
  wire WX663;
  wire WX664;
  wire WX665;
  wire WX666;
  wire WX667;
  wire WX668;
  wire WX669;
  wire WX670;
  wire WX671;
  wire WX672;
  wire WX673;
  wire WX674;
  wire WX675;
  wire WX676;
  wire WX677;
  wire WX678;
  wire WX679;
  wire WX680;
  wire WX681;
  wire WX682;
  wire WX683;
  wire WX684;
  wire WX685;
  wire WX686;
  wire WX687;
  wire WX688;
  wire WX689;
  wire WX690;
  wire WX691;
  wire WX692;
  wire WX693;
  wire WX694;
  wire WX6949;
  wire WX695;
  wire WX6950;
  wire WX6951;
  wire WX6952;
  wire WX6953;
  wire WX6954;
  wire WX6955;
  wire WX6956;
  wire WX6957;
  wire WX6958;
  wire WX6959;
  wire WX696;
  wire WX6960;
  wire WX6961;
  wire WX6962;
  wire WX6963;
  wire WX6964;
  wire WX6965;
  wire WX6966;
  wire WX6967;
  wire WX6968;
  wire WX6969;
  wire WX697;
  wire WX6970;
  wire WX6971;
  wire WX6972;
  wire WX6973;
  wire WX6974;
  wire WX6975;
  wire WX6976;
  wire WX6977;
  wire WX6978;
  wire WX6979;
  wire WX698;
  wire WX6980;
  wire WX6981;
  wire WX6982;
  wire WX6983;
  wire WX6984;
  wire WX6985;
  wire WX6986;
  wire WX6987;
  wire WX6988;
  wire WX6989;
  wire WX699;
  wire WX6990;
  wire WX6991;
  wire WX6992;
  wire WX6993;
  wire WX6994;
  wire WX6995;
  wire WX6996;
  wire WX6997;
  wire WX6998;
  wire WX6999;
  wire WX700;
  wire WX7000;
  wire WX7001;
  wire WX7002;
  wire WX7003;
  wire WX7004;
  wire WX7005;
  wire WX7006;
  wire WX7007;
  wire WX7008;
  wire WX7009;
  wire WX701;
  wire WX7010;
  wire WX7011;
  wire WX7012;
  wire WX702;
  wire WX703;
  wire WX704;
  wire WX705;
  wire WX706;
  wire WX707;
  wire WX708;
  wire WX709;
  wire WX710;
  wire WX7109;
  wire WX711;
  wire WX7110;
  wire WX7111;
  wire WX7112;
  wire WX7113;
  wire WX7114;
  wire WX7115;
  wire WX7116;
  wire WX7117;
  wire WX7118;
  wire WX7119;
  wire WX712;
  wire WX7120;
  wire WX7121;
  wire WX7122;
  wire WX7123;
  wire WX7124;
  wire WX7125;
  wire WX7126;
  wire WX7127;
  wire WX7128;
  wire WX7129;
  wire WX713;
  wire WX7130;
  wire WX7131;
  wire WX7132;
  wire WX7133;
  wire WX7134;
  wire WX7135;
  wire WX7136;
  wire WX7137;
  wire WX7138;
  wire WX7139;
  wire WX714;
  wire WX7140;
  wire WX7141;
  wire WX7142;
  wire WX7143;
  wire WX7144;
  wire WX7145;
  wire WX7146;
  wire WX7147;
  wire WX7148;
  wire WX7149;
  wire WX715;
  wire WX7150;
  wire WX7151;
  wire WX7152;
  wire WX7153;
  wire WX7154;
  wire WX7155;
  wire WX7156;
  wire WX7157;
  wire WX7158;
  wire WX7159;
  wire WX716;
  wire WX7160;
  wire WX7161;
  wire WX7162;
  wire WX7163;
  wire WX7164;
  wire WX7165;
  wire WX7166;
  wire WX7167;
  wire WX7168;
  wire WX7169;
  wire WX717;
  wire WX7170;
  wire WX7171;
  wire WX7172;
  wire WX7173;
  wire WX7174;
  wire WX7175;
  wire WX7176;
  wire WX7177;
  wire WX7178;
  wire WX7179;
  wire WX718;
  wire WX7180;
  wire WX7181;
  wire WX7182;
  wire WX7183;
  wire WX7184;
  wire WX7185;
  wire WX7186;
  wire WX7187;
  wire WX7188;
  wire WX7189;
  wire WX719;
  wire WX7190;
  wire WX7191;
  wire WX7192;
  wire WX7193;
  wire WX7194;
  wire WX7195;
  wire WX7196;
  wire WX7197;
  wire WX7198;
  wire WX7199;
  wire WX720;
  wire WX7200;
  wire WX7201;
  wire WX7202;
  wire WX7203;
  wire WX7204;
  wire WX7205;
  wire WX7206;
  wire WX7207;
  wire WX7208;
  wire WX7209;
  wire WX721;
  wire WX7210;
  wire WX7211;
  wire WX7212;
  wire WX7213;
  wire WX7214;
  wire WX7215;
  wire WX7216;
  wire WX7217;
  wire WX7218;
  wire WX7219;
  wire WX722;
  wire WX7220;
  wire WX7221;
  wire WX7222;
  wire WX7223;
  wire WX7224;
  wire WX7225;
  wire WX7226;
  wire WX7227;
  wire WX7228;
  wire WX7229;
  wire WX723;
  wire WX7230;
  wire WX7231;
  wire WX7232;
  wire WX7233;
  wire WX7234;
  wire WX7235;
  wire WX7236;
  wire WX7237;
  wire WX7238;
  wire WX7239;
  wire WX724;
  wire WX7240;
  wire WX7241;
  wire WX7242;
  wire WX7243;
  wire WX7244;
  wire WX7245;
  wire WX7246;
  wire WX7247;
  wire WX7248;
  wire WX7249;
  wire WX725;
  wire WX7250;
  wire WX7251;
  wire WX7252;
  wire WX7253;
  wire WX7254;
  wire WX7255;
  wire WX7256;
  wire WX7257;
  wire WX7258;
  wire WX7259;
  wire WX726;
  wire WX7260;
  wire WX7261;
  wire WX7262;
  wire WX7263;
  wire WX7264;
  wire WX7265;
  wire WX7266;
  wire WX7267;
  wire WX7268;
  wire WX7269;
  wire WX727;
  wire WX7270;
  wire WX7271;
  wire WX7272;
  wire WX7273;
  wire WX7274;
  wire WX7275;
  wire WX7276;
  wire WX7277;
  wire WX7278;
  wire WX7279;
  wire WX728;
  wire WX7280;
  wire WX7281;
  wire WX7282;
  wire WX7283;
  wire WX7284;
  wire WX7285;
  wire WX7286;
  wire WX7287;
  wire WX7288;
  wire WX7289;
  wire WX729;
  wire WX7290;
  wire WX7291;
  wire WX7292;
  wire WX7293;
  wire WX7294;
  wire WX7295;
  wire WX7296;
  wire WX7297;
  wire WX7298;
  wire WX7299;
  wire WX730;
  wire WX7300;
  wire WX7301;
  wire WX7302;
  wire WX7303;
  wire WX7304;
  wire WX7305;
  wire WX7306;
  wire WX7307;
  wire WX7308;
  wire WX7309;
  wire WX731;
  wire WX7310;
  wire WX7311;
  wire WX7312;
  wire WX7313;
  wire WX7314;
  wire WX7315;
  wire WX7316;
  wire WX7317;
  wire WX7318;
  wire WX7319;
  wire WX732;
  wire WX7320;
  wire WX7321;
  wire WX7322;
  wire WX7323;
  wire WX7324;
  wire WX7325;
  wire WX7326;
  wire WX7327;
  wire WX7328;
  wire WX7329;
  wire WX733;
  wire WX7330;
  wire WX7331;
  wire WX7332;
  wire WX7333;
  wire WX7334;
  wire WX7335;
  wire WX7336;
  wire WX7337;
  wire WX7338;
  wire WX7339;
  wire WX734;
  wire WX7340;
  wire WX7341;
  wire WX7342;
  wire WX7343;
  wire WX7344;
  wire WX7345;
  wire WX7346;
  wire WX7347;
  wire WX7348;
  wire WX7349;
  wire WX735;
  wire WX7350;
  wire WX7351;
  wire WX7352;
  wire WX7353;
  wire WX7354;
  wire WX7355;
  wire WX7356;
  wire WX7357;
  wire WX7358;
  wire WX7359;
  wire WX736;
  wire WX7360;
  wire WX7361;
  wire WX7362;
  wire WX7363;
  wire WX7364;
  wire WX737;
  wire WX738;
  wire WX739;
  wire WX740;
  wire WX741;
  wire WX742;
  wire WX743;
  wire WX744;
  wire WX745;
  wire WX746;
  wire WX7466;
  wire WX7467;
  wire WX7468;
  wire WX7469;
  wire WX747;
  wire WX7470;
  wire WX748;
  wire WX749;
  wire WX750;
  wire WX751;
  wire WX752;
  wire WX753;
  wire WX754;
  wire WX755;
  wire WX756;
  wire WX757;
  wire WX758;
  wire WX759;
  wire WX760;
  wire WX761;
  wire WX762;
  wire WX763;
  wire WX764;
  wire WX765;
  wire WX766;
  wire WX767;
  wire WX768;
  wire WX769;
  wire WX770;
  wire WX771;
  wire WX772;
  wire WX7728;
  wire WX7729;
  wire WX773;
  wire WX7731;
  wire WX7733;
  wire WX7735;
  wire WX7737;
  wire WX7739;
  wire WX774;
  wire WX7741;
  wire WX7743;
  wire WX7745;
  wire WX7747;
  wire WX7749;
  wire WX775;
  wire WX7751;
  wire WX7753;
  wire WX7755;
  wire WX7757;
  wire WX7759;
  wire WX776;
  wire WX7761;
  wire WX7763;
  wire WX7765;
  wire WX7767;
  wire WX7769;
  wire WX777;
  wire WX7771;
  wire WX7773;
  wire WX7775;
  wire WX7777;
  wire WX7779;
  wire WX778;
  wire WX7781;
  wire WX7783;
  wire WX7785;
  wire WX7787;
  wire WX7789;
  wire WX779;
  wire WX7791;
  wire WX780;
  wire WX781;
  wire WX782;
  wire WX783;
  wire WX784;
  wire WX785;
  wire WX786;
  wire WX787;
  wire WX788;
  wire WX789;
  wire WX790;
  wire WX791;
  wire WX792;
  wire WX793;
  wire WX794;
  wire WX795;
  wire WX796;
  wire WX797;
  wire WX798;
  wire WX799;
  wire WX800;
  wire WX801;
  wire WX802;
  wire WX803;
  wire WX804;
  wire WX805;
  wire WX806;
  wire WX807;
  wire WX808;
  wire WX809;
  wire WX810;
  wire WX811;
  wire WX812;
  wire WX813;
  wire WX814;
  wire WX815;
  wire WX816;
  wire WX817;
  wire WX818;
  wire WX819;
  wire WX820;
  wire WX821;
  wire WX822;
  wire WX823;
  wire WX824;
  wire WX8242;
  wire WX8243;
  wire WX8244;
  wire WX8245;
  wire WX8246;
  wire WX8247;
  wire WX8248;
  wire WX8249;
  wire WX825;
  wire WX8250;
  wire WX8251;
  wire WX8252;
  wire WX8253;
  wire WX8254;
  wire WX8255;
  wire WX8256;
  wire WX8257;
  wire WX8258;
  wire WX8259;
  wire WX826;
  wire WX8260;
  wire WX8261;
  wire WX8262;
  wire WX8263;
  wire WX8264;
  wire WX8265;
  wire WX8266;
  wire WX8267;
  wire WX8268;
  wire WX8269;
  wire WX827;
  wire WX8270;
  wire WX8271;
  wire WX8272;
  wire WX8273;
  wire WX8274;
  wire WX8275;
  wire WX8276;
  wire WX8277;
  wire WX8278;
  wire WX8279;
  wire WX828;
  wire WX8280;
  wire WX8281;
  wire WX8282;
  wire WX8283;
  wire WX8284;
  wire WX8285;
  wire WX8286;
  wire WX8287;
  wire WX8288;
  wire WX8289;
  wire WX829;
  wire WX8290;
  wire WX8291;
  wire WX8292;
  wire WX8293;
  wire WX8294;
  wire WX8295;
  wire WX8296;
  wire WX8297;
  wire WX8298;
  wire WX8299;
  wire WX830;
  wire WX8300;
  wire WX8301;
  wire WX8302;
  wire WX8303;
  wire WX8304;
  wire WX8305;
  wire WX831;
  wire WX832;
  wire WX833;
  wire WX834;
  wire WX835;
  wire WX836;
  wire WX837;
  wire WX838;
  wire WX839;
  wire WX840;
  wire WX8402;
  wire WX8403;
  wire WX8404;
  wire WX8405;
  wire WX8406;
  wire WX8407;
  wire WX8408;
  wire WX8409;
  wire WX841;
  wire WX8410;
  wire WX8411;
  wire WX8412;
  wire WX8413;
  wire WX8414;
  wire WX8415;
  wire WX8416;
  wire WX8417;
  wire WX8418;
  wire WX8419;
  wire WX842;
  wire WX8420;
  wire WX8421;
  wire WX8422;
  wire WX8423;
  wire WX8424;
  wire WX8425;
  wire WX8426;
  wire WX8427;
  wire WX8428;
  wire WX8429;
  wire WX843;
  wire WX8430;
  wire WX8431;
  wire WX8432;
  wire WX8433;
  wire WX8434;
  wire WX8435;
  wire WX8436;
  wire WX8437;
  wire WX8438;
  wire WX8439;
  wire WX844;
  wire WX8440;
  wire WX8441;
  wire WX8442;
  wire WX8443;
  wire WX8444;
  wire WX8445;
  wire WX8446;
  wire WX8447;
  wire WX8448;
  wire WX8449;
  wire WX845;
  wire WX8450;
  wire WX8451;
  wire WX8452;
  wire WX8453;
  wire WX8454;
  wire WX8455;
  wire WX8456;
  wire WX8457;
  wire WX8458;
  wire WX8459;
  wire WX846;
  wire WX8460;
  wire WX8461;
  wire WX8462;
  wire WX8463;
  wire WX8464;
  wire WX8465;
  wire WX8466;
  wire WX8467;
  wire WX8468;
  wire WX8469;
  wire WX847;
  wire WX8470;
  wire WX8471;
  wire WX8472;
  wire WX8473;
  wire WX8474;
  wire WX8475;
  wire WX8476;
  wire WX8477;
  wire WX8478;
  wire WX8479;
  wire WX848;
  wire WX8480;
  wire WX8481;
  wire WX8482;
  wire WX8483;
  wire WX8484;
  wire WX8485;
  wire WX8486;
  wire WX8487;
  wire WX8488;
  wire WX8489;
  wire WX849;
  wire WX8490;
  wire WX8491;
  wire WX8492;
  wire WX8493;
  wire WX8494;
  wire WX8495;
  wire WX8496;
  wire WX8497;
  wire WX8498;
  wire WX8499;
  wire WX850;
  wire WX8500;
  wire WX8501;
  wire WX8502;
  wire WX8503;
  wire WX8504;
  wire WX8505;
  wire WX8506;
  wire WX8507;
  wire WX8508;
  wire WX8509;
  wire WX851;
  wire WX8510;
  wire WX8511;
  wire WX8512;
  wire WX8513;
  wire WX8514;
  wire WX8515;
  wire WX8516;
  wire WX8517;
  wire WX8518;
  wire WX8519;
  wire WX852;
  wire WX8520;
  wire WX8521;
  wire WX8522;
  wire WX8523;
  wire WX8524;
  wire WX8525;
  wire WX8526;
  wire WX8527;
  wire WX8528;
  wire WX8529;
  wire WX853;
  wire WX8530;
  wire WX8531;
  wire WX8532;
  wire WX8533;
  wire WX8534;
  wire WX8535;
  wire WX8536;
  wire WX8537;
  wire WX8538;
  wire WX8539;
  wire WX854;
  wire WX8540;
  wire WX8541;
  wire WX8542;
  wire WX8543;
  wire WX8544;
  wire WX8545;
  wire WX8546;
  wire WX8547;
  wire WX8548;
  wire WX8549;
  wire WX855;
  wire WX8550;
  wire WX8551;
  wire WX8552;
  wire WX8553;
  wire WX8554;
  wire WX8555;
  wire WX8556;
  wire WX8557;
  wire WX8558;
  wire WX8559;
  wire WX856;
  wire WX8560;
  wire WX8561;
  wire WX8562;
  wire WX8563;
  wire WX8564;
  wire WX8565;
  wire WX8566;
  wire WX8567;
  wire WX8568;
  wire WX8569;
  wire WX857;
  wire WX8570;
  wire WX8571;
  wire WX8572;
  wire WX8573;
  wire WX8574;
  wire WX8575;
  wire WX8576;
  wire WX8577;
  wire WX8578;
  wire WX8579;
  wire WX858;
  wire WX8580;
  wire WX8581;
  wire WX8582;
  wire WX8583;
  wire WX8584;
  wire WX8585;
  wire WX8586;
  wire WX8587;
  wire WX8588;
  wire WX8589;
  wire WX859;
  wire WX8590;
  wire WX8591;
  wire WX8592;
  wire WX8593;
  wire WX8594;
  wire WX8595;
  wire WX8596;
  wire WX8597;
  wire WX8598;
  wire WX8599;
  wire WX860;
  wire WX8600;
  wire WX8601;
  wire WX8602;
  wire WX8603;
  wire WX8604;
  wire WX8605;
  wire WX8606;
  wire WX8607;
  wire WX8608;
  wire WX8609;
  wire WX861;
  wire WX8610;
  wire WX8611;
  wire WX8612;
  wire WX8613;
  wire WX8614;
  wire WX8615;
  wire WX8616;
  wire WX8617;
  wire WX8618;
  wire WX8619;
  wire WX862;
  wire WX8620;
  wire WX8621;
  wire WX8622;
  wire WX8623;
  wire WX8624;
  wire WX8625;
  wire WX8626;
  wire WX8627;
  wire WX8628;
  wire WX8629;
  wire WX863;
  wire WX8630;
  wire WX8631;
  wire WX8632;
  wire WX8633;
  wire WX8634;
  wire WX8635;
  wire WX8636;
  wire WX8637;
  wire WX8638;
  wire WX8639;
  wire WX864;
  wire WX8640;
  wire WX8641;
  wire WX8642;
  wire WX8643;
  wire WX8644;
  wire WX8645;
  wire WX8646;
  wire WX8647;
  wire WX8648;
  wire WX8649;
  wire WX865;
  wire WX8650;
  wire WX8651;
  wire WX8652;
  wire WX8653;
  wire WX8654;
  wire WX8655;
  wire WX8656;
  wire WX8657;
  wire WX866;
  wire WX867;
  wire WX868;
  wire WX869;
  wire WX870;
  wire WX871;
  wire WX872;
  wire WX873;
  wire WX874;
  wire WX875;
  wire WX8759;
  wire WX876;
  wire WX8760;
  wire WX8761;
  wire WX8762;
  wire WX8763;
  wire WX877;
  wire WX878;
  wire WX879;
  wire WX880;
  wire WX881;
  wire WX882;
  wire WX883;
  wire WX884;
  wire WX885;
  wire WX886;
  wire WX887;
  wire WX888;
  wire WX889;
  wire WX890;
  wire WX891;
  wire WX892;
  wire WX893;
  wire WX894;
  wire WX895;
  wire WX896;
  wire WX897;
  wire WX898;
  wire WX899;
  wire WX9021;
  wire WX9022;
  wire WX9024;
  wire WX9026;
  wire WX9028;
  wire WX9030;
  wire WX9032;
  wire WX9034;
  wire WX9036;
  wire WX9038;
  wire WX9040;
  wire WX9042;
  wire WX9044;
  wire WX9046;
  wire WX9048;
  wire WX9050;
  wire WX9052;
  wire WX9054;
  wire WX9056;
  wire WX9058;
  wire WX9060;
  wire WX9062;
  wire WX9064;
  wire WX9066;
  wire WX9068;
  wire WX9070;
  wire WX9072;
  wire WX9074;
  wire WX9076;
  wire WX9078;
  wire WX9080;
  wire WX9082;
  wire WX9084;
  wire WX9535;
  wire WX9536;
  wire WX9537;
  wire WX9538;
  wire WX9539;
  wire WX9540;
  wire WX9541;
  wire WX9542;
  wire WX9543;
  wire WX9544;
  wire WX9545;
  wire WX9546;
  wire WX9547;
  wire WX9548;
  wire WX9549;
  wire WX9550;
  wire WX9551;
  wire WX9552;
  wire WX9553;
  wire WX9554;
  wire WX9555;
  wire WX9556;
  wire WX9557;
  wire WX9558;
  wire WX9559;
  wire WX9560;
  wire WX9561;
  wire WX9562;
  wire WX9563;
  wire WX9564;
  wire WX9565;
  wire WX9566;
  wire WX9567;
  wire WX9568;
  wire WX9569;
  wire WX9570;
  wire WX9571;
  wire WX9572;
  wire WX9573;
  wire WX9574;
  wire WX9575;
  wire WX9576;
  wire WX9577;
  wire WX9578;
  wire WX9579;
  wire WX9580;
  wire WX9581;
  wire WX9582;
  wire WX9583;
  wire WX9584;
  wire WX9585;
  wire WX9586;
  wire WX9587;
  wire WX9588;
  wire WX9589;
  wire WX9590;
  wire WX9591;
  wire WX9592;
  wire WX9593;
  wire WX9594;
  wire WX9595;
  wire WX9596;
  wire WX9597;
  wire WX9598;
  wire WX9695;
  wire WX9696;
  wire WX9697;
  wire WX9698;
  wire WX9699;
  wire WX9700;
  wire WX9701;
  wire WX9702;
  wire WX9703;
  wire WX9704;
  wire WX9705;
  wire WX9706;
  wire WX9707;
  wire WX9708;
  wire WX9709;
  wire WX9710;
  wire WX9711;
  wire WX9712;
  wire WX9713;
  wire WX9714;
  wire WX9715;
  wire WX9716;
  wire WX9717;
  wire WX9718;
  wire WX9719;
  wire WX9720;
  wire WX9721;
  wire WX9722;
  wire WX9723;
  wire WX9724;
  wire WX9725;
  wire WX9726;
  wire WX9727;
  wire WX9728;
  wire WX9729;
  wire WX9730;
  wire WX9731;
  wire WX9732;
  wire WX9733;
  wire WX9734;
  wire WX9735;
  wire WX9736;
  wire WX9737;
  wire WX9738;
  wire WX9739;
  wire WX9740;
  wire WX9741;
  wire WX9742;
  wire WX9743;
  wire WX9744;
  wire WX9745;
  wire WX9746;
  wire WX9747;
  wire WX9748;
  wire WX9749;
  wire WX9750;
  wire WX9751;
  wire WX9752;
  wire WX9753;
  wire WX9754;
  wire WX9755;
  wire WX9756;
  wire WX9757;
  wire WX9758;
  wire WX9759;
  wire WX9760;
  wire WX9761;
  wire WX9762;
  wire WX9763;
  wire WX9764;
  wire WX9765;
  wire WX9766;
  wire WX9767;
  wire WX9768;
  wire WX9769;
  wire WX9770;
  wire WX9771;
  wire WX9772;
  wire WX9773;
  wire WX9774;
  wire WX9775;
  wire WX9776;
  wire WX9777;
  wire WX9778;
  wire WX9779;
  wire WX9780;
  wire WX9781;
  wire WX9782;
  wire WX9783;
  wire WX9784;
  wire WX9785;
  wire WX9786;
  wire WX9787;
  wire WX9788;
  wire WX9789;
  wire WX9790;
  wire WX9791;
  wire WX9792;
  wire WX9793;
  wire WX9794;
  wire WX9795;
  wire WX9796;
  wire WX9797;
  wire WX9798;
  wire WX9799;
  wire WX9800;
  wire WX9801;
  wire WX9802;
  wire WX9803;
  wire WX9804;
  wire WX9805;
  wire WX9806;
  wire WX9807;
  wire WX9808;
  wire WX9809;
  wire WX9810;
  wire WX9811;
  wire WX9812;
  wire WX9813;
  wire WX9814;
  wire WX9815;
  wire WX9816;
  wire WX9817;
  wire WX9818;
  wire WX9819;
  wire WX9820;
  wire WX9821;
  wire WX9822;
  wire WX9823;
  wire WX9824;
  wire WX9825;
  wire WX9826;
  wire WX9827;
  wire WX9828;
  wire WX9829;
  wire WX9830;
  wire WX9831;
  wire WX9832;
  wire WX9833;
  wire WX9834;
  wire WX9835;
  wire WX9836;
  wire WX9837;
  wire WX9838;
  wire WX9839;
  wire WX9840;
  wire WX9841;
  wire WX9842;
  wire WX9843;
  wire WX9844;
  wire WX9845;
  wire WX9846;
  wire WX9847;
  wire WX9848;
  wire WX9849;
  wire WX9850;
  wire WX9851;
  wire WX9852;
  wire WX9853;
  wire WX9854;
  wire WX9855;
  wire WX9856;
  wire WX9857;
  wire WX9858;
  wire WX9859;
  wire WX9860;
  wire WX9861;
  wire WX9862;
  wire WX9863;
  wire WX9864;
  wire WX9865;
  wire WX9866;
  wire WX9867;
  wire WX9868;
  wire WX9869;
  wire WX9870;
  wire WX9871;
  wire WX9872;
  wire WX9873;
  wire WX9874;
  wire WX9875;
  wire WX9876;
  wire WX9877;
  wire WX9878;
  wire WX9879;
  wire WX9880;
  wire WX9881;
  wire WX9882;
  wire WX9883;
  wire WX9884;
  wire WX9885;
  wire WX9886;
  wire WX9887;
  wire WX9888;
  wire WX9889;
  wire WX9890;
  wire WX9891;
  wire WX9892;
  wire WX9893;
  wire WX9894;
  wire WX9895;
  wire WX9896;
  wire WX9897;
  wire WX9898;
  wire WX9899;
  wire WX9900;
  wire WX9901;
  wire WX9902;
  wire WX9903;
  wire WX9904;
  wire WX9905;
  wire WX9906;
  wire WX9907;
  wire WX9908;
  wire WX9909;
  wire WX9910;
  wire WX9911;
  wire WX9912;
  wire WX9913;
  wire WX9914;
  wire WX9915;
  wire WX9916;
  wire WX9917;
  wire WX9918;
  wire WX9919;
  wire WX9920;
  wire WX9921;
  wire WX9922;
  wire WX9923;
  wire WX9924;
  wire WX9925;
  wire WX9926;
  wire WX9927;
  wire WX9928;
  wire WX9929;
  wire WX9930;
  wire WX9931;
  wire WX9932;
  wire WX9933;
  wire WX9934;
  wire WX9935;
  wire WX9936;
  wire WX9937;
  wire WX9938;
  wire WX9939;
  wire WX9940;
  wire WX9941;
  wire WX9942;
  wire WX9943;
  wire WX9944;
  wire WX9945;
  wire WX9946;
  wire WX9947;
  wire WX9948;
  wire WX9949;
  wire WX9950;
  al_and2ft _04452_ (
    .a(\DFF_64.Q ),
    .b(\DFF_96.Q ),
    .y(_00000_)
  );
  al_and2ft _04453_ (
    .a(\DFF_96.Q ),
    .b(\DFF_64.Q ),
    .y(_00001_)
  );
  al_or2 _04454_ (
    .a(_00000_),
    .b(_00001_),
    .y(_00002_)
  );
  al_nand2ft _04455_ (
    .a(\DFF_32.Q ),
    .b(TM1),
    .y(_00003_)
  );
  al_nand2ft _04456_ (
    .a(TM1),
    .b(\DFF_32.Q ),
    .y(_00004_)
  );
  al_or3fft _04457_ (
    .a(_00003_),
    .b(_00004_),
    .c(_00002_),
    .y(_00005_)
  );
  al_ao21ttf _04458_ (
    .a(_00003_),
    .b(_00004_),
    .c(_00002_),
    .y(_00006_)
  );
  al_ao21ttf _04459_ (
    .a(\DFF_0.Q ),
    .b(TM0),
    .c(\DFF_128.Q ),
    .y(_00007_)
  );
  al_and3ftt _04460_ (
    .a(\DFF_128.Q ),
    .b(\DFF_0.Q ),
    .c(TM0),
    .y(_00008_)
  );
  al_and2ft _04461_ (
    .a(_00008_),
    .b(_00007_),
    .y(_00009_)
  );
  al_nand3ftt _04462_ (
    .a(_00009_),
    .b(_00006_),
    .c(_00005_),
    .y(_00010_)
  );
  al_ao21 _04463_ (
    .a(_00003_),
    .b(_00004_),
    .c(_00002_),
    .y(_00011_)
  );
  al_nand3 _04464_ (
    .a(_00003_),
    .b(_00004_),
    .c(_00002_),
    .y(_00012_)
  );
  al_nand3 _04465_ (
    .a(_00009_),
    .b(_00012_),
    .c(_00011_),
    .y(_00013_)
  );
  al_and2 _04466_ (
    .a(_00013_),
    .b(_00010_),
    .y(DATA_9_31)
  );
  al_and2ft _04467_ (
    .a(\DFF_65.Q ),
    .b(\DFF_97.Q ),
    .y(_00014_)
  );
  al_and2ft _04468_ (
    .a(\DFF_97.Q ),
    .b(\DFF_65.Q ),
    .y(_00015_)
  );
  al_or2 _04469_ (
    .a(_00014_),
    .b(_00015_),
    .y(_00016_)
  );
  al_nand2ft _04470_ (
    .a(\DFF_33.Q ),
    .b(TM1),
    .y(_00017_)
  );
  al_nand2ft _04471_ (
    .a(TM1),
    .b(\DFF_33.Q ),
    .y(_00018_)
  );
  al_or3fft _04472_ (
    .a(_00017_),
    .b(_00018_),
    .c(_00016_),
    .y(_00019_)
  );
  al_ao21ttf _04473_ (
    .a(_00017_),
    .b(_00018_),
    .c(_00016_),
    .y(_00020_)
  );
  al_ao21ttf _04474_ (
    .a(TM0),
    .b(\DFF_1.Q ),
    .c(\DFF_129.Q ),
    .y(_00021_)
  );
  al_and3ftt _04475_ (
    .a(\DFF_129.Q ),
    .b(TM0),
    .c(\DFF_1.Q ),
    .y(_00022_)
  );
  al_and2ft _04476_ (
    .a(_00022_),
    .b(_00021_),
    .y(_00023_)
  );
  al_nand3ftt _04477_ (
    .a(_00023_),
    .b(_00020_),
    .c(_00019_),
    .y(_00024_)
  );
  al_ao21 _04478_ (
    .a(_00017_),
    .b(_00018_),
    .c(_00016_),
    .y(_00025_)
  );
  al_nand3 _04479_ (
    .a(_00017_),
    .b(_00018_),
    .c(_00016_),
    .y(_00026_)
  );
  al_nand3 _04480_ (
    .a(_00023_),
    .b(_00026_),
    .c(_00025_),
    .y(_00027_)
  );
  al_and2 _04481_ (
    .a(_00027_),
    .b(_00024_),
    .y(DATA_9_30)
  );
  al_and2ft _04482_ (
    .a(\DFF_66.Q ),
    .b(\DFF_98.Q ),
    .y(_00028_)
  );
  al_and2ft _04483_ (
    .a(\DFF_98.Q ),
    .b(\DFF_66.Q ),
    .y(_00029_)
  );
  al_or2 _04484_ (
    .a(_00028_),
    .b(_00029_),
    .y(_00030_)
  );
  al_nand2ft _04485_ (
    .a(\DFF_34.Q ),
    .b(TM1),
    .y(_00031_)
  );
  al_nand2ft _04486_ (
    .a(TM1),
    .b(\DFF_34.Q ),
    .y(_00032_)
  );
  al_or3fft _04487_ (
    .a(_00031_),
    .b(_00032_),
    .c(_00030_),
    .y(_00033_)
  );
  al_ao21ttf _04488_ (
    .a(_00031_),
    .b(_00032_),
    .c(_00030_),
    .y(_00034_)
  );
  al_ao21ttf _04489_ (
    .a(TM0),
    .b(\DFF_2.Q ),
    .c(\DFF_130.Q ),
    .y(_00035_)
  );
  al_and3ftt _04490_ (
    .a(\DFF_130.Q ),
    .b(TM0),
    .c(\DFF_2.Q ),
    .y(_00036_)
  );
  al_and2ft _04491_ (
    .a(_00036_),
    .b(_00035_),
    .y(_00037_)
  );
  al_nand3ftt _04492_ (
    .a(_00037_),
    .b(_00034_),
    .c(_00033_),
    .y(_00038_)
  );
  al_ao21 _04493_ (
    .a(_00031_),
    .b(_00032_),
    .c(_00030_),
    .y(_00039_)
  );
  al_nand3 _04494_ (
    .a(_00031_),
    .b(_00032_),
    .c(_00030_),
    .y(_00040_)
  );
  al_nand3 _04495_ (
    .a(_00037_),
    .b(_00040_),
    .c(_00039_),
    .y(_00041_)
  );
  al_and2 _04496_ (
    .a(_00041_),
    .b(_00038_),
    .y(DATA_9_29)
  );
  al_and2ft _04497_ (
    .a(\DFF_67.Q ),
    .b(\DFF_99.Q ),
    .y(_00042_)
  );
  al_and2ft _04498_ (
    .a(\DFF_99.Q ),
    .b(\DFF_67.Q ),
    .y(_00043_)
  );
  al_or2 _04499_ (
    .a(_00042_),
    .b(_00043_),
    .y(_00044_)
  );
  al_nand2ft _04500_ (
    .a(\DFF_35.Q ),
    .b(TM1),
    .y(_00045_)
  );
  al_nand2ft _04501_ (
    .a(TM1),
    .b(\DFF_35.Q ),
    .y(_00046_)
  );
  al_or3fft _04502_ (
    .a(_00045_),
    .b(_00046_),
    .c(_00044_),
    .y(_00047_)
  );
  al_ao21ttf _04503_ (
    .a(_00045_),
    .b(_00046_),
    .c(_00044_),
    .y(_00048_)
  );
  al_ao21ttf _04504_ (
    .a(TM0),
    .b(\DFF_3.Q ),
    .c(\DFF_131.Q ),
    .y(_00049_)
  );
  al_and3ftt _04505_ (
    .a(\DFF_131.Q ),
    .b(TM0),
    .c(\DFF_3.Q ),
    .y(_00050_)
  );
  al_and2ft _04506_ (
    .a(_00050_),
    .b(_00049_),
    .y(_00051_)
  );
  al_nand3ftt _04507_ (
    .a(_00051_),
    .b(_00048_),
    .c(_00047_),
    .y(_00052_)
  );
  al_ao21 _04508_ (
    .a(_00045_),
    .b(_00046_),
    .c(_00044_),
    .y(_00053_)
  );
  al_nand3 _04509_ (
    .a(_00045_),
    .b(_00046_),
    .c(_00044_),
    .y(_00054_)
  );
  al_nand3 _04510_ (
    .a(_00051_),
    .b(_00054_),
    .c(_00053_),
    .y(_00055_)
  );
  al_and2 _04511_ (
    .a(_00055_),
    .b(_00052_),
    .y(DATA_9_28)
  );
  al_and2ft _04512_ (
    .a(\DFF_68.Q ),
    .b(\DFF_100.Q ),
    .y(_00056_)
  );
  al_and2ft _04513_ (
    .a(\DFF_100.Q ),
    .b(\DFF_68.Q ),
    .y(_00057_)
  );
  al_or2 _04514_ (
    .a(_00056_),
    .b(_00057_),
    .y(_00058_)
  );
  al_nand2ft _04515_ (
    .a(\DFF_36.Q ),
    .b(TM1),
    .y(_00059_)
  );
  al_nand2ft _04516_ (
    .a(TM1),
    .b(\DFF_36.Q ),
    .y(_00060_)
  );
  al_or3fft _04517_ (
    .a(_00059_),
    .b(_00060_),
    .c(_00058_),
    .y(_00061_)
  );
  al_ao21ttf _04518_ (
    .a(_00059_),
    .b(_00060_),
    .c(_00058_),
    .y(_00062_)
  );
  al_ao21ttf _04519_ (
    .a(TM0),
    .b(\DFF_4.Q ),
    .c(\DFF_132.Q ),
    .y(_00063_)
  );
  al_and3ftt _04520_ (
    .a(\DFF_132.Q ),
    .b(TM0),
    .c(\DFF_4.Q ),
    .y(_00064_)
  );
  al_and2ft _04521_ (
    .a(_00064_),
    .b(_00063_),
    .y(_00065_)
  );
  al_nand3ftt _04522_ (
    .a(_00065_),
    .b(_00062_),
    .c(_00061_),
    .y(_00066_)
  );
  al_ao21 _04523_ (
    .a(_00059_),
    .b(_00060_),
    .c(_00058_),
    .y(_00067_)
  );
  al_nand3 _04524_ (
    .a(_00059_),
    .b(_00060_),
    .c(_00058_),
    .y(_00068_)
  );
  al_nand3 _04525_ (
    .a(_00065_),
    .b(_00068_),
    .c(_00067_),
    .y(_00069_)
  );
  al_and2 _04526_ (
    .a(_00069_),
    .b(_00066_),
    .y(DATA_9_27)
  );
  al_and2ft _04527_ (
    .a(\DFF_69.Q ),
    .b(\DFF_101.Q ),
    .y(_00070_)
  );
  al_and2ft _04528_ (
    .a(\DFF_101.Q ),
    .b(\DFF_69.Q ),
    .y(_00071_)
  );
  al_or2 _04529_ (
    .a(_00070_),
    .b(_00071_),
    .y(_00072_)
  );
  al_nand2ft _04530_ (
    .a(\DFF_37.Q ),
    .b(TM1),
    .y(_00073_)
  );
  al_nand2ft _04531_ (
    .a(TM1),
    .b(\DFF_37.Q ),
    .y(_00074_)
  );
  al_or3fft _04532_ (
    .a(_00073_),
    .b(_00074_),
    .c(_00072_),
    .y(_00075_)
  );
  al_ao21ttf _04533_ (
    .a(_00073_),
    .b(_00074_),
    .c(_00072_),
    .y(_00076_)
  );
  al_ao21ttf _04534_ (
    .a(TM0),
    .b(\DFF_5.Q ),
    .c(\DFF_133.Q ),
    .y(_00077_)
  );
  al_and3ftt _04535_ (
    .a(\DFF_133.Q ),
    .b(TM0),
    .c(\DFF_5.Q ),
    .y(_00078_)
  );
  al_and2ft _04536_ (
    .a(_00078_),
    .b(_00077_),
    .y(_00079_)
  );
  al_nand3ftt _04537_ (
    .a(_00079_),
    .b(_00076_),
    .c(_00075_),
    .y(_00080_)
  );
  al_ao21 _04538_ (
    .a(_00073_),
    .b(_00074_),
    .c(_00072_),
    .y(_00081_)
  );
  al_nand3 _04539_ (
    .a(_00073_),
    .b(_00074_),
    .c(_00072_),
    .y(_00082_)
  );
  al_nand3 _04540_ (
    .a(_00079_),
    .b(_00082_),
    .c(_00081_),
    .y(_00083_)
  );
  al_and2 _04541_ (
    .a(_00083_),
    .b(_00080_),
    .y(DATA_9_26)
  );
  al_and2ft _04542_ (
    .a(\DFF_70.Q ),
    .b(\DFF_102.Q ),
    .y(_00084_)
  );
  al_and2ft _04543_ (
    .a(\DFF_102.Q ),
    .b(\DFF_70.Q ),
    .y(_00085_)
  );
  al_or2 _04544_ (
    .a(_00084_),
    .b(_00085_),
    .y(_00086_)
  );
  al_nand2ft _04545_ (
    .a(\DFF_38.Q ),
    .b(TM1),
    .y(_00087_)
  );
  al_nand2ft _04546_ (
    .a(TM1),
    .b(\DFF_38.Q ),
    .y(_00088_)
  );
  al_or3fft _04547_ (
    .a(_00087_),
    .b(_00088_),
    .c(_00086_),
    .y(_00089_)
  );
  al_ao21ttf _04548_ (
    .a(_00087_),
    .b(_00088_),
    .c(_00086_),
    .y(_00090_)
  );
  al_ao21ttf _04549_ (
    .a(TM0),
    .b(\DFF_6.Q ),
    .c(\DFF_134.Q ),
    .y(_00091_)
  );
  al_and3ftt _04550_ (
    .a(\DFF_134.Q ),
    .b(TM0),
    .c(\DFF_6.Q ),
    .y(_00092_)
  );
  al_and2ft _04551_ (
    .a(_00092_),
    .b(_00091_),
    .y(_00093_)
  );
  al_nand3ftt _04552_ (
    .a(_00093_),
    .b(_00090_),
    .c(_00089_),
    .y(_00094_)
  );
  al_ao21 _04553_ (
    .a(_00087_),
    .b(_00088_),
    .c(_00086_),
    .y(_00095_)
  );
  al_nand3 _04554_ (
    .a(_00087_),
    .b(_00088_),
    .c(_00086_),
    .y(_00096_)
  );
  al_nand3 _04555_ (
    .a(_00093_),
    .b(_00096_),
    .c(_00095_),
    .y(_00097_)
  );
  al_and2 _04556_ (
    .a(_00097_),
    .b(_00094_),
    .y(DATA_9_25)
  );
  al_and2ft _04557_ (
    .a(\DFF_71.Q ),
    .b(\DFF_103.Q ),
    .y(_00098_)
  );
  al_and2ft _04558_ (
    .a(\DFF_103.Q ),
    .b(\DFF_71.Q ),
    .y(_00099_)
  );
  al_or2 _04559_ (
    .a(_00098_),
    .b(_00099_),
    .y(_00100_)
  );
  al_nand2ft _04560_ (
    .a(\DFF_39.Q ),
    .b(TM1),
    .y(_00101_)
  );
  al_nand2ft _04561_ (
    .a(TM1),
    .b(\DFF_39.Q ),
    .y(_00102_)
  );
  al_or3fft _04562_ (
    .a(_00101_),
    .b(_00102_),
    .c(_00100_),
    .y(_00103_)
  );
  al_ao21ttf _04563_ (
    .a(_00101_),
    .b(_00102_),
    .c(_00100_),
    .y(_00104_)
  );
  al_ao21ttf _04564_ (
    .a(TM0),
    .b(\DFF_7.Q ),
    .c(\DFF_135.Q ),
    .y(_00105_)
  );
  al_and3ftt _04565_ (
    .a(\DFF_135.Q ),
    .b(TM0),
    .c(\DFF_7.Q ),
    .y(_00106_)
  );
  al_and2ft _04566_ (
    .a(_00106_),
    .b(_00105_),
    .y(_00107_)
  );
  al_nand3ftt _04567_ (
    .a(_00107_),
    .b(_00104_),
    .c(_00103_),
    .y(_00108_)
  );
  al_ao21 _04568_ (
    .a(_00101_),
    .b(_00102_),
    .c(_00100_),
    .y(_00109_)
  );
  al_nand3 _04569_ (
    .a(_00101_),
    .b(_00102_),
    .c(_00100_),
    .y(_00110_)
  );
  al_nand3 _04570_ (
    .a(_00107_),
    .b(_00110_),
    .c(_00109_),
    .y(_00111_)
  );
  al_and2 _04571_ (
    .a(_00111_),
    .b(_00108_),
    .y(DATA_9_24)
  );
  al_and2ft _04572_ (
    .a(\DFF_72.Q ),
    .b(\DFF_104.Q ),
    .y(_00112_)
  );
  al_and2ft _04573_ (
    .a(\DFF_104.Q ),
    .b(\DFF_72.Q ),
    .y(_00113_)
  );
  al_or2 _04574_ (
    .a(_00112_),
    .b(_00113_),
    .y(_00114_)
  );
  al_nand2ft _04575_ (
    .a(\DFF_40.Q ),
    .b(TM1),
    .y(_00115_)
  );
  al_nand2ft _04576_ (
    .a(TM1),
    .b(\DFF_40.Q ),
    .y(_00116_)
  );
  al_or3fft _04577_ (
    .a(_00115_),
    .b(_00116_),
    .c(_00114_),
    .y(_00117_)
  );
  al_ao21ttf _04578_ (
    .a(_00115_),
    .b(_00116_),
    .c(_00114_),
    .y(_00118_)
  );
  al_ao21ttf _04579_ (
    .a(TM0),
    .b(\DFF_8.Q ),
    .c(\DFF_136.Q ),
    .y(_00119_)
  );
  al_and3ftt _04580_ (
    .a(\DFF_136.Q ),
    .b(TM0),
    .c(\DFF_8.Q ),
    .y(_00120_)
  );
  al_and2ft _04581_ (
    .a(_00120_),
    .b(_00119_),
    .y(_00121_)
  );
  al_nand3ftt _04582_ (
    .a(_00121_),
    .b(_00118_),
    .c(_00117_),
    .y(_00122_)
  );
  al_ao21 _04583_ (
    .a(_00115_),
    .b(_00116_),
    .c(_00114_),
    .y(_00123_)
  );
  al_nand3 _04584_ (
    .a(_00115_),
    .b(_00116_),
    .c(_00114_),
    .y(_00124_)
  );
  al_nand3 _04585_ (
    .a(_00121_),
    .b(_00124_),
    .c(_00123_),
    .y(_00125_)
  );
  al_and2 _04586_ (
    .a(_00125_),
    .b(_00122_),
    .y(DATA_9_23)
  );
  al_and2ft _04587_ (
    .a(\DFF_73.Q ),
    .b(\DFF_105.Q ),
    .y(_00126_)
  );
  al_and2ft _04588_ (
    .a(\DFF_105.Q ),
    .b(\DFF_73.Q ),
    .y(_00127_)
  );
  al_or2 _04589_ (
    .a(_00126_),
    .b(_00127_),
    .y(_00128_)
  );
  al_nand2ft _04590_ (
    .a(\DFF_41.Q ),
    .b(TM1),
    .y(_00129_)
  );
  al_nand2ft _04591_ (
    .a(TM1),
    .b(\DFF_41.Q ),
    .y(_00130_)
  );
  al_or3fft _04592_ (
    .a(_00129_),
    .b(_00130_),
    .c(_00128_),
    .y(_00131_)
  );
  al_ao21ttf _04593_ (
    .a(_00129_),
    .b(_00130_),
    .c(_00128_),
    .y(_00132_)
  );
  al_ao21ttf _04594_ (
    .a(TM0),
    .b(\DFF_9.Q ),
    .c(\DFF_137.Q ),
    .y(_00133_)
  );
  al_and3ftt _04595_ (
    .a(\DFF_137.Q ),
    .b(TM0),
    .c(\DFF_9.Q ),
    .y(_00134_)
  );
  al_and2ft _04596_ (
    .a(_00134_),
    .b(_00133_),
    .y(_00135_)
  );
  al_nand3ftt _04597_ (
    .a(_00135_),
    .b(_00132_),
    .c(_00131_),
    .y(_00136_)
  );
  al_ao21 _04598_ (
    .a(_00129_),
    .b(_00130_),
    .c(_00128_),
    .y(_00137_)
  );
  al_nand3 _04599_ (
    .a(_00129_),
    .b(_00130_),
    .c(_00128_),
    .y(_00138_)
  );
  al_nand3 _04600_ (
    .a(_00135_),
    .b(_00138_),
    .c(_00137_),
    .y(_00139_)
  );
  al_and2 _04601_ (
    .a(_00139_),
    .b(_00136_),
    .y(DATA_9_22)
  );
  al_and2ft _04602_ (
    .a(\DFF_74.Q ),
    .b(\DFF_106.Q ),
    .y(_00140_)
  );
  al_and2ft _04603_ (
    .a(\DFF_106.Q ),
    .b(\DFF_74.Q ),
    .y(_00141_)
  );
  al_or2 _04604_ (
    .a(_00140_),
    .b(_00141_),
    .y(_00142_)
  );
  al_nand2ft _04605_ (
    .a(\DFF_42.Q ),
    .b(TM1),
    .y(_00143_)
  );
  al_nand2ft _04606_ (
    .a(TM1),
    .b(\DFF_42.Q ),
    .y(_00144_)
  );
  al_or3fft _04607_ (
    .a(_00143_),
    .b(_00144_),
    .c(_00142_),
    .y(_00145_)
  );
  al_ao21ttf _04608_ (
    .a(_00143_),
    .b(_00144_),
    .c(_00142_),
    .y(_00146_)
  );
  al_ao21ttf _04609_ (
    .a(TM0),
    .b(\DFF_10.Q ),
    .c(\DFF_138.Q ),
    .y(_00147_)
  );
  al_and3ftt _04610_ (
    .a(\DFF_138.Q ),
    .b(TM0),
    .c(\DFF_10.Q ),
    .y(_00148_)
  );
  al_and2ft _04611_ (
    .a(_00148_),
    .b(_00147_),
    .y(_00149_)
  );
  al_nand3ftt _04612_ (
    .a(_00149_),
    .b(_00146_),
    .c(_00145_),
    .y(_00150_)
  );
  al_ao21 _04613_ (
    .a(_00143_),
    .b(_00144_),
    .c(_00142_),
    .y(_00151_)
  );
  al_nand3 _04614_ (
    .a(_00143_),
    .b(_00144_),
    .c(_00142_),
    .y(_00152_)
  );
  al_nand3 _04615_ (
    .a(_00149_),
    .b(_00152_),
    .c(_00151_),
    .y(_00153_)
  );
  al_and2 _04616_ (
    .a(_00153_),
    .b(_00150_),
    .y(DATA_9_21)
  );
  al_and2ft _04617_ (
    .a(\DFF_75.Q ),
    .b(\DFF_107.Q ),
    .y(_00154_)
  );
  al_and2ft _04618_ (
    .a(\DFF_107.Q ),
    .b(\DFF_75.Q ),
    .y(_00155_)
  );
  al_or2 _04619_ (
    .a(_00154_),
    .b(_00155_),
    .y(_00156_)
  );
  al_nand2ft _04620_ (
    .a(\DFF_43.Q ),
    .b(TM1),
    .y(_00157_)
  );
  al_nand2ft _04621_ (
    .a(TM1),
    .b(\DFF_43.Q ),
    .y(_00158_)
  );
  al_or3fft _04622_ (
    .a(_00157_),
    .b(_00158_),
    .c(_00156_),
    .y(_00159_)
  );
  al_ao21ttf _04623_ (
    .a(_00157_),
    .b(_00158_),
    .c(_00156_),
    .y(_00160_)
  );
  al_ao21ttf _04624_ (
    .a(TM0),
    .b(\DFF_11.Q ),
    .c(\DFF_139.Q ),
    .y(_00161_)
  );
  al_and3ftt _04625_ (
    .a(\DFF_139.Q ),
    .b(TM0),
    .c(\DFF_11.Q ),
    .y(_00162_)
  );
  al_and2ft _04626_ (
    .a(_00162_),
    .b(_00161_),
    .y(_00163_)
  );
  al_nand3ftt _04627_ (
    .a(_00163_),
    .b(_00160_),
    .c(_00159_),
    .y(_00164_)
  );
  al_ao21 _04628_ (
    .a(_00157_),
    .b(_00158_),
    .c(_00156_),
    .y(_00165_)
  );
  al_nand3 _04629_ (
    .a(_00157_),
    .b(_00158_),
    .c(_00156_),
    .y(_00166_)
  );
  al_nand3 _04630_ (
    .a(_00163_),
    .b(_00166_),
    .c(_00165_),
    .y(_00167_)
  );
  al_and2 _04631_ (
    .a(_00167_),
    .b(_00164_),
    .y(DATA_9_20)
  );
  al_and2ft _04632_ (
    .a(\DFF_76.Q ),
    .b(\DFF_108.Q ),
    .y(_00168_)
  );
  al_and2ft _04633_ (
    .a(\DFF_108.Q ),
    .b(\DFF_76.Q ),
    .y(_00169_)
  );
  al_or2 _04634_ (
    .a(_00168_),
    .b(_00169_),
    .y(_00170_)
  );
  al_nand2ft _04635_ (
    .a(\DFF_44.Q ),
    .b(TM1),
    .y(_00171_)
  );
  al_nand2ft _04636_ (
    .a(TM1),
    .b(\DFF_44.Q ),
    .y(_00172_)
  );
  al_or3fft _04637_ (
    .a(_00171_),
    .b(_00172_),
    .c(_00170_),
    .y(_00173_)
  );
  al_ao21ttf _04638_ (
    .a(_00171_),
    .b(_00172_),
    .c(_00170_),
    .y(_00174_)
  );
  al_ao21ttf _04639_ (
    .a(TM0),
    .b(\DFF_12.Q ),
    .c(\DFF_140.Q ),
    .y(_00175_)
  );
  al_and3ftt _04640_ (
    .a(\DFF_140.Q ),
    .b(TM0),
    .c(\DFF_12.Q ),
    .y(_00176_)
  );
  al_and2ft _04641_ (
    .a(_00176_),
    .b(_00175_),
    .y(_00177_)
  );
  al_nand3ftt _04642_ (
    .a(_00177_),
    .b(_00174_),
    .c(_00173_),
    .y(_00178_)
  );
  al_ao21 _04643_ (
    .a(_00171_),
    .b(_00172_),
    .c(_00170_),
    .y(_00179_)
  );
  al_nand3 _04644_ (
    .a(_00171_),
    .b(_00172_),
    .c(_00170_),
    .y(_00180_)
  );
  al_nand3 _04645_ (
    .a(_00177_),
    .b(_00180_),
    .c(_00179_),
    .y(_00181_)
  );
  al_and2 _04646_ (
    .a(_00181_),
    .b(_00178_),
    .y(DATA_9_19)
  );
  al_and2ft _04647_ (
    .a(\DFF_77.Q ),
    .b(\DFF_109.Q ),
    .y(_00182_)
  );
  al_and2ft _04648_ (
    .a(\DFF_109.Q ),
    .b(\DFF_77.Q ),
    .y(_00183_)
  );
  al_or2 _04649_ (
    .a(_00182_),
    .b(_00183_),
    .y(_00184_)
  );
  al_nand2ft _04650_ (
    .a(\DFF_45.Q ),
    .b(TM1),
    .y(_00185_)
  );
  al_nand2ft _04651_ (
    .a(TM1),
    .b(\DFF_45.Q ),
    .y(_00186_)
  );
  al_or3fft _04652_ (
    .a(_00185_),
    .b(_00186_),
    .c(_00184_),
    .y(_00187_)
  );
  al_ao21ttf _04653_ (
    .a(_00185_),
    .b(_00186_),
    .c(_00184_),
    .y(_00188_)
  );
  al_ao21ttf _04654_ (
    .a(TM0),
    .b(\DFF_13.Q ),
    .c(\DFF_141.Q ),
    .y(_00189_)
  );
  al_and3ftt _04655_ (
    .a(\DFF_141.Q ),
    .b(TM0),
    .c(\DFF_13.Q ),
    .y(_00190_)
  );
  al_and2ft _04656_ (
    .a(_00190_),
    .b(_00189_),
    .y(_00191_)
  );
  al_nand3ftt _04657_ (
    .a(_00191_),
    .b(_00188_),
    .c(_00187_),
    .y(_00192_)
  );
  al_ao21 _04658_ (
    .a(_00185_),
    .b(_00186_),
    .c(_00184_),
    .y(_00193_)
  );
  al_nand3 _04659_ (
    .a(_00185_),
    .b(_00186_),
    .c(_00184_),
    .y(_00194_)
  );
  al_nand3 _04660_ (
    .a(_00191_),
    .b(_00194_),
    .c(_00193_),
    .y(_00195_)
  );
  al_and2 _04661_ (
    .a(_00195_),
    .b(_00192_),
    .y(DATA_9_18)
  );
  al_and2ft _04662_ (
    .a(\DFF_78.Q ),
    .b(\DFF_110.Q ),
    .y(_00196_)
  );
  al_and2ft _04663_ (
    .a(\DFF_110.Q ),
    .b(\DFF_78.Q ),
    .y(_00197_)
  );
  al_or2 _04664_ (
    .a(_00196_),
    .b(_00197_),
    .y(_00198_)
  );
  al_nand2ft _04665_ (
    .a(\DFF_46.Q ),
    .b(TM1),
    .y(_00199_)
  );
  al_nand2ft _04666_ (
    .a(TM1),
    .b(\DFF_46.Q ),
    .y(_00200_)
  );
  al_or3fft _04667_ (
    .a(_00199_),
    .b(_00200_),
    .c(_00198_),
    .y(_00201_)
  );
  al_ao21ttf _04668_ (
    .a(_00199_),
    .b(_00200_),
    .c(_00198_),
    .y(_00202_)
  );
  al_ao21ttf _04669_ (
    .a(TM0),
    .b(\DFF_14.Q ),
    .c(\DFF_142.Q ),
    .y(_00203_)
  );
  al_and3ftt _04670_ (
    .a(\DFF_142.Q ),
    .b(TM0),
    .c(\DFF_14.Q ),
    .y(_00204_)
  );
  al_and2ft _04671_ (
    .a(_00204_),
    .b(_00203_),
    .y(_00205_)
  );
  al_nand3ftt _04672_ (
    .a(_00205_),
    .b(_00202_),
    .c(_00201_),
    .y(_00206_)
  );
  al_ao21 _04673_ (
    .a(_00199_),
    .b(_00200_),
    .c(_00198_),
    .y(_00207_)
  );
  al_nand3 _04674_ (
    .a(_00199_),
    .b(_00200_),
    .c(_00198_),
    .y(_00208_)
  );
  al_nand3 _04675_ (
    .a(_00205_),
    .b(_00208_),
    .c(_00207_),
    .y(_00209_)
  );
  al_and2 _04676_ (
    .a(_00209_),
    .b(_00206_),
    .y(DATA_9_17)
  );
  al_and2ft _04677_ (
    .a(\DFF_79.Q ),
    .b(\DFF_111.Q ),
    .y(_00210_)
  );
  al_and2ft _04678_ (
    .a(\DFF_111.Q ),
    .b(\DFF_79.Q ),
    .y(_00211_)
  );
  al_or2 _04679_ (
    .a(_00210_),
    .b(_00211_),
    .y(_00212_)
  );
  al_nand2ft _04680_ (
    .a(\DFF_47.Q ),
    .b(TM1),
    .y(_00213_)
  );
  al_nand2ft _04681_ (
    .a(TM1),
    .b(\DFF_47.Q ),
    .y(_00214_)
  );
  al_or3fft _04682_ (
    .a(_00213_),
    .b(_00214_),
    .c(_00212_),
    .y(_00215_)
  );
  al_ao21ttf _04683_ (
    .a(_00213_),
    .b(_00214_),
    .c(_00212_),
    .y(_00216_)
  );
  al_ao21ttf _04684_ (
    .a(TM0),
    .b(\DFF_15.Q ),
    .c(\DFF_143.Q ),
    .y(_00217_)
  );
  al_and3ftt _04685_ (
    .a(\DFF_143.Q ),
    .b(TM0),
    .c(\DFF_15.Q ),
    .y(_00218_)
  );
  al_and2ft _04686_ (
    .a(_00218_),
    .b(_00217_),
    .y(_00219_)
  );
  al_nand3ftt _04687_ (
    .a(_00219_),
    .b(_00216_),
    .c(_00215_),
    .y(_00220_)
  );
  al_ao21 _04688_ (
    .a(_00213_),
    .b(_00214_),
    .c(_00212_),
    .y(_00221_)
  );
  al_nand3 _04689_ (
    .a(_00213_),
    .b(_00214_),
    .c(_00212_),
    .y(_00222_)
  );
  al_nand3 _04690_ (
    .a(_00219_),
    .b(_00222_),
    .c(_00221_),
    .y(_00223_)
  );
  al_and2 _04691_ (
    .a(_00223_),
    .b(_00220_),
    .y(DATA_9_16)
  );
  al_and2ft _04692_ (
    .a(\DFF_80.Q ),
    .b(\DFF_112.Q ),
    .y(_00224_)
  );
  al_and2ft _04693_ (
    .a(\DFF_112.Q ),
    .b(\DFF_80.Q ),
    .y(_00225_)
  );
  al_or2 _04694_ (
    .a(_00224_),
    .b(_00225_),
    .y(_00226_)
  );
  al_nand2ft _04695_ (
    .a(\DFF_48.Q ),
    .b(TM0),
    .y(_00227_)
  );
  al_nand2ft _04696_ (
    .a(TM0),
    .b(\DFF_48.Q ),
    .y(_00228_)
  );
  al_or3fft _04697_ (
    .a(_00227_),
    .b(_00228_),
    .c(_00226_),
    .y(_00229_)
  );
  al_ao21ttf _04698_ (
    .a(_00227_),
    .b(_00228_),
    .c(_00226_),
    .y(_00230_)
  );
  al_ao21ttf _04699_ (
    .a(TM0),
    .b(\DFF_16.Q ),
    .c(\DFF_144.Q ),
    .y(_00231_)
  );
  al_and3ftt _04700_ (
    .a(\DFF_144.Q ),
    .b(TM0),
    .c(\DFF_16.Q ),
    .y(_00232_)
  );
  al_and2ft _04701_ (
    .a(_00232_),
    .b(_00231_),
    .y(_00233_)
  );
  al_nand3ftt _04702_ (
    .a(_00233_),
    .b(_00230_),
    .c(_00229_),
    .y(_00234_)
  );
  al_ao21 _04703_ (
    .a(_00227_),
    .b(_00228_),
    .c(_00226_),
    .y(_00235_)
  );
  al_nand3 _04704_ (
    .a(_00227_),
    .b(_00228_),
    .c(_00226_),
    .y(_00236_)
  );
  al_nand3 _04705_ (
    .a(_00233_),
    .b(_00236_),
    .c(_00235_),
    .y(_00237_)
  );
  al_and2 _04706_ (
    .a(_00237_),
    .b(_00234_),
    .y(DATA_9_15)
  );
  al_and2ft _04707_ (
    .a(\DFF_81.Q ),
    .b(\DFF_113.Q ),
    .y(_00238_)
  );
  al_and2ft _04708_ (
    .a(\DFF_113.Q ),
    .b(\DFF_81.Q ),
    .y(_00239_)
  );
  al_or2 _04709_ (
    .a(_00238_),
    .b(_00239_),
    .y(_00240_)
  );
  al_nand2ft _04710_ (
    .a(\DFF_49.Q ),
    .b(TM0),
    .y(_00241_)
  );
  al_nand2ft _04711_ (
    .a(TM0),
    .b(\DFF_49.Q ),
    .y(_00242_)
  );
  al_or3fft _04712_ (
    .a(_00241_),
    .b(_00242_),
    .c(_00240_),
    .y(_00243_)
  );
  al_ao21ttf _04713_ (
    .a(_00241_),
    .b(_00242_),
    .c(_00240_),
    .y(_00244_)
  );
  al_ao21ttf _04714_ (
    .a(TM0),
    .b(\DFF_17.Q ),
    .c(\DFF_145.Q ),
    .y(_00245_)
  );
  al_and3ftt _04715_ (
    .a(\DFF_145.Q ),
    .b(TM0),
    .c(\DFF_17.Q ),
    .y(_00246_)
  );
  al_and2ft _04716_ (
    .a(_00246_),
    .b(_00245_),
    .y(_00247_)
  );
  al_nand3ftt _04717_ (
    .a(_00247_),
    .b(_00244_),
    .c(_00243_),
    .y(_00248_)
  );
  al_ao21 _04718_ (
    .a(_00241_),
    .b(_00242_),
    .c(_00240_),
    .y(_00249_)
  );
  al_nand3 _04719_ (
    .a(_00241_),
    .b(_00242_),
    .c(_00240_),
    .y(_00250_)
  );
  al_nand3 _04720_ (
    .a(_00247_),
    .b(_00250_),
    .c(_00249_),
    .y(_00251_)
  );
  al_and2 _04721_ (
    .a(_00251_),
    .b(_00248_),
    .y(DATA_9_14)
  );
  al_and2ft _04722_ (
    .a(\DFF_82.Q ),
    .b(\DFF_114.Q ),
    .y(_00252_)
  );
  al_and2ft _04723_ (
    .a(\DFF_114.Q ),
    .b(\DFF_82.Q ),
    .y(_00253_)
  );
  al_or2 _04724_ (
    .a(_00252_),
    .b(_00253_),
    .y(_00254_)
  );
  al_nand2ft _04725_ (
    .a(\DFF_50.Q ),
    .b(TM0),
    .y(_00255_)
  );
  al_nand2ft _04726_ (
    .a(TM0),
    .b(\DFF_50.Q ),
    .y(_00256_)
  );
  al_or3fft _04727_ (
    .a(_00255_),
    .b(_00256_),
    .c(_00254_),
    .y(_00257_)
  );
  al_ao21ttf _04728_ (
    .a(_00255_),
    .b(_00256_),
    .c(_00254_),
    .y(_00258_)
  );
  al_ao21ttf _04729_ (
    .a(TM0),
    .b(\DFF_18.Q ),
    .c(\DFF_146.Q ),
    .y(_00259_)
  );
  al_and3ftt _04730_ (
    .a(\DFF_146.Q ),
    .b(TM0),
    .c(\DFF_18.Q ),
    .y(_00260_)
  );
  al_and2ft _04731_ (
    .a(_00260_),
    .b(_00259_),
    .y(_00261_)
  );
  al_nand3ftt _04732_ (
    .a(_00261_),
    .b(_00258_),
    .c(_00257_),
    .y(_00262_)
  );
  al_ao21 _04733_ (
    .a(_00255_),
    .b(_00256_),
    .c(_00254_),
    .y(_00263_)
  );
  al_nand3 _04734_ (
    .a(_00255_),
    .b(_00256_),
    .c(_00254_),
    .y(_00264_)
  );
  al_nand3 _04735_ (
    .a(_00261_),
    .b(_00264_),
    .c(_00263_),
    .y(_00265_)
  );
  al_and2 _04736_ (
    .a(_00265_),
    .b(_00262_),
    .y(DATA_9_13)
  );
  al_and2ft _04737_ (
    .a(\DFF_83.Q ),
    .b(\DFF_115.Q ),
    .y(_00266_)
  );
  al_and2ft _04738_ (
    .a(\DFF_115.Q ),
    .b(\DFF_83.Q ),
    .y(_00267_)
  );
  al_or2 _04739_ (
    .a(_00266_),
    .b(_00267_),
    .y(_00268_)
  );
  al_nand2ft _04740_ (
    .a(\DFF_51.Q ),
    .b(TM0),
    .y(_00269_)
  );
  al_nand2ft _04741_ (
    .a(TM0),
    .b(\DFF_51.Q ),
    .y(_00270_)
  );
  al_or3fft _04742_ (
    .a(_00269_),
    .b(_00270_),
    .c(_00268_),
    .y(_00271_)
  );
  al_ao21ttf _04743_ (
    .a(_00269_),
    .b(_00270_),
    .c(_00268_),
    .y(_00272_)
  );
  al_ao21ttf _04744_ (
    .a(TM0),
    .b(\DFF_19.Q ),
    .c(\DFF_147.Q ),
    .y(_00273_)
  );
  al_and3ftt _04745_ (
    .a(\DFF_147.Q ),
    .b(TM0),
    .c(\DFF_19.Q ),
    .y(_00274_)
  );
  al_and2ft _04746_ (
    .a(_00274_),
    .b(_00273_),
    .y(_00275_)
  );
  al_nand3ftt _04747_ (
    .a(_00275_),
    .b(_00272_),
    .c(_00271_),
    .y(_00276_)
  );
  al_ao21 _04748_ (
    .a(_00269_),
    .b(_00270_),
    .c(_00268_),
    .y(_00277_)
  );
  al_nand3 _04749_ (
    .a(_00269_),
    .b(_00270_),
    .c(_00268_),
    .y(_00278_)
  );
  al_nand3 _04750_ (
    .a(_00275_),
    .b(_00278_),
    .c(_00277_),
    .y(_00279_)
  );
  al_and2 _04751_ (
    .a(_00279_),
    .b(_00276_),
    .y(DATA_9_12)
  );
  al_and2ft _04752_ (
    .a(\DFF_84.Q ),
    .b(\DFF_116.Q ),
    .y(_00280_)
  );
  al_and2ft _04753_ (
    .a(\DFF_116.Q ),
    .b(\DFF_84.Q ),
    .y(_00281_)
  );
  al_or2 _04754_ (
    .a(_00280_),
    .b(_00281_),
    .y(_00282_)
  );
  al_nand2ft _04755_ (
    .a(\DFF_52.Q ),
    .b(TM0),
    .y(_00283_)
  );
  al_nand2ft _04756_ (
    .a(TM0),
    .b(\DFF_52.Q ),
    .y(_00284_)
  );
  al_or3fft _04757_ (
    .a(_00283_),
    .b(_00284_),
    .c(_00282_),
    .y(_00285_)
  );
  al_ao21ttf _04758_ (
    .a(_00283_),
    .b(_00284_),
    .c(_00282_),
    .y(_00286_)
  );
  al_ao21ttf _04759_ (
    .a(TM0),
    .b(\DFF_20.Q ),
    .c(\DFF_148.Q ),
    .y(_00287_)
  );
  al_and3ftt _04760_ (
    .a(\DFF_148.Q ),
    .b(TM0),
    .c(\DFF_20.Q ),
    .y(_00288_)
  );
  al_and2ft _04761_ (
    .a(_00288_),
    .b(_00287_),
    .y(_00289_)
  );
  al_nand3ftt _04762_ (
    .a(_00289_),
    .b(_00286_),
    .c(_00285_),
    .y(_00290_)
  );
  al_ao21 _04763_ (
    .a(_00283_),
    .b(_00284_),
    .c(_00282_),
    .y(_00291_)
  );
  al_nand3 _04764_ (
    .a(_00283_),
    .b(_00284_),
    .c(_00282_),
    .y(_00292_)
  );
  al_nand3 _04765_ (
    .a(_00289_),
    .b(_00292_),
    .c(_00291_),
    .y(_00293_)
  );
  al_and2 _04766_ (
    .a(_00293_),
    .b(_00290_),
    .y(DATA_9_11)
  );
  al_and2ft _04767_ (
    .a(\DFF_85.Q ),
    .b(\DFF_117.Q ),
    .y(_00294_)
  );
  al_and2ft _04768_ (
    .a(\DFF_117.Q ),
    .b(\DFF_85.Q ),
    .y(_00295_)
  );
  al_or2 _04769_ (
    .a(_00294_),
    .b(_00295_),
    .y(_00296_)
  );
  al_nand2ft _04770_ (
    .a(\DFF_53.Q ),
    .b(TM0),
    .y(_00297_)
  );
  al_nand2ft _04771_ (
    .a(TM0),
    .b(\DFF_53.Q ),
    .y(_00298_)
  );
  al_or3fft _04772_ (
    .a(_00297_),
    .b(_00298_),
    .c(_00296_),
    .y(_00299_)
  );
  al_ao21ttf _04773_ (
    .a(_00297_),
    .b(_00298_),
    .c(_00296_),
    .y(_00300_)
  );
  al_ao21ttf _04774_ (
    .a(TM0),
    .b(\DFF_21.Q ),
    .c(\DFF_149.Q ),
    .y(_00301_)
  );
  al_and3ftt _04775_ (
    .a(\DFF_149.Q ),
    .b(TM0),
    .c(\DFF_21.Q ),
    .y(_00302_)
  );
  al_and2ft _04776_ (
    .a(_00302_),
    .b(_00301_),
    .y(_00303_)
  );
  al_nand3ftt _04777_ (
    .a(_00303_),
    .b(_00300_),
    .c(_00299_),
    .y(_00304_)
  );
  al_ao21 _04778_ (
    .a(_00297_),
    .b(_00298_),
    .c(_00296_),
    .y(_00305_)
  );
  al_nand3 _04779_ (
    .a(_00297_),
    .b(_00298_),
    .c(_00296_),
    .y(_00306_)
  );
  al_nand3 _04780_ (
    .a(_00303_),
    .b(_00306_),
    .c(_00305_),
    .y(_00307_)
  );
  al_and2 _04781_ (
    .a(_00307_),
    .b(_00304_),
    .y(DATA_9_10)
  );
  al_and2ft _04782_ (
    .a(\DFF_86.Q ),
    .b(\DFF_118.Q ),
    .y(_00308_)
  );
  al_and2ft _04783_ (
    .a(\DFF_118.Q ),
    .b(\DFF_86.Q ),
    .y(_00309_)
  );
  al_or2 _04784_ (
    .a(_00308_),
    .b(_00309_),
    .y(_00310_)
  );
  al_nand2ft _04785_ (
    .a(\DFF_54.Q ),
    .b(TM0),
    .y(_00311_)
  );
  al_nand2ft _04786_ (
    .a(TM0),
    .b(\DFF_54.Q ),
    .y(_00312_)
  );
  al_or3fft _04787_ (
    .a(_00311_),
    .b(_00312_),
    .c(_00310_),
    .y(_00313_)
  );
  al_ao21ttf _04788_ (
    .a(_00311_),
    .b(_00312_),
    .c(_00310_),
    .y(_00314_)
  );
  al_ao21ttf _04789_ (
    .a(TM0),
    .b(\DFF_22.Q ),
    .c(\DFF_150.Q ),
    .y(_00315_)
  );
  al_and3ftt _04790_ (
    .a(\DFF_150.Q ),
    .b(TM0),
    .c(\DFF_22.Q ),
    .y(_00316_)
  );
  al_and2ft _04791_ (
    .a(_00316_),
    .b(_00315_),
    .y(_00317_)
  );
  al_nand3ftt _04792_ (
    .a(_00317_),
    .b(_00314_),
    .c(_00313_),
    .y(_00318_)
  );
  al_ao21 _04793_ (
    .a(_00311_),
    .b(_00312_),
    .c(_00310_),
    .y(_00319_)
  );
  al_nand3 _04794_ (
    .a(_00311_),
    .b(_00312_),
    .c(_00310_),
    .y(_00320_)
  );
  al_nand3 _04795_ (
    .a(_00317_),
    .b(_00320_),
    .c(_00319_),
    .y(_00321_)
  );
  al_and2 _04796_ (
    .a(_00321_),
    .b(_00318_),
    .y(DATA_9_9)
  );
  al_and2ft _04797_ (
    .a(\DFF_87.Q ),
    .b(\DFF_119.Q ),
    .y(_00322_)
  );
  al_and2ft _04798_ (
    .a(\DFF_119.Q ),
    .b(\DFF_87.Q ),
    .y(_00323_)
  );
  al_or2 _04799_ (
    .a(_00322_),
    .b(_00323_),
    .y(_00324_)
  );
  al_nand2ft _04800_ (
    .a(\DFF_55.Q ),
    .b(TM0),
    .y(_00325_)
  );
  al_nand2ft _04801_ (
    .a(TM0),
    .b(\DFF_55.Q ),
    .y(_00326_)
  );
  al_or3fft _04802_ (
    .a(_00325_),
    .b(_00326_),
    .c(_00324_),
    .y(_00327_)
  );
  al_ao21ttf _04803_ (
    .a(_00325_),
    .b(_00326_),
    .c(_00324_),
    .y(_00328_)
  );
  al_ao21ttf _04804_ (
    .a(TM0),
    .b(\DFF_23.Q ),
    .c(\DFF_151.Q ),
    .y(_00329_)
  );
  al_and3ftt _04805_ (
    .a(\DFF_151.Q ),
    .b(TM0),
    .c(\DFF_23.Q ),
    .y(_00330_)
  );
  al_and2ft _04806_ (
    .a(_00330_),
    .b(_00329_),
    .y(_00331_)
  );
  al_nand3ftt _04807_ (
    .a(_00331_),
    .b(_00328_),
    .c(_00327_),
    .y(_00332_)
  );
  al_ao21 _04808_ (
    .a(_00325_),
    .b(_00326_),
    .c(_00324_),
    .y(_00333_)
  );
  al_nand3 _04809_ (
    .a(_00325_),
    .b(_00326_),
    .c(_00324_),
    .y(_00334_)
  );
  al_nand3 _04810_ (
    .a(_00331_),
    .b(_00334_),
    .c(_00333_),
    .y(_00335_)
  );
  al_and2 _04811_ (
    .a(_00335_),
    .b(_00332_),
    .y(DATA_9_8)
  );
  al_and2ft _04812_ (
    .a(\DFF_88.Q ),
    .b(\DFF_120.Q ),
    .y(_00336_)
  );
  al_and2ft _04813_ (
    .a(\DFF_120.Q ),
    .b(\DFF_88.Q ),
    .y(_00337_)
  );
  al_or2 _04814_ (
    .a(_00336_),
    .b(_00337_),
    .y(_00338_)
  );
  al_nand2ft _04815_ (
    .a(\DFF_56.Q ),
    .b(TM0),
    .y(_00339_)
  );
  al_nand2ft _04816_ (
    .a(TM0),
    .b(\DFF_56.Q ),
    .y(_00340_)
  );
  al_or3fft _04817_ (
    .a(_00339_),
    .b(_00340_),
    .c(_00338_),
    .y(_00341_)
  );
  al_ao21ttf _04818_ (
    .a(_00339_),
    .b(_00340_),
    .c(_00338_),
    .y(_00342_)
  );
  al_ao21ttf _04819_ (
    .a(TM0),
    .b(\DFF_24.Q ),
    .c(\DFF_152.Q ),
    .y(_00343_)
  );
  al_and3ftt _04820_ (
    .a(\DFF_152.Q ),
    .b(TM0),
    .c(\DFF_24.Q ),
    .y(_00344_)
  );
  al_and2ft _04821_ (
    .a(_00344_),
    .b(_00343_),
    .y(_00345_)
  );
  al_nand3ftt _04822_ (
    .a(_00345_),
    .b(_00342_),
    .c(_00341_),
    .y(_00346_)
  );
  al_ao21 _04823_ (
    .a(_00339_),
    .b(_00340_),
    .c(_00338_),
    .y(_00347_)
  );
  al_nand3 _04824_ (
    .a(_00339_),
    .b(_00340_),
    .c(_00338_),
    .y(_00348_)
  );
  al_nand3 _04825_ (
    .a(_00345_),
    .b(_00348_),
    .c(_00347_),
    .y(_00349_)
  );
  al_and2 _04826_ (
    .a(_00349_),
    .b(_00346_),
    .y(DATA_9_7)
  );
  al_and2ft _04827_ (
    .a(\DFF_89.Q ),
    .b(\DFF_121.Q ),
    .y(_00350_)
  );
  al_and2ft _04828_ (
    .a(\DFF_121.Q ),
    .b(\DFF_89.Q ),
    .y(_00351_)
  );
  al_or2 _04829_ (
    .a(_00350_),
    .b(_00351_),
    .y(_00352_)
  );
  al_nand2ft _04830_ (
    .a(\DFF_57.Q ),
    .b(TM0),
    .y(_00353_)
  );
  al_nand2ft _04831_ (
    .a(TM0),
    .b(\DFF_57.Q ),
    .y(_00354_)
  );
  al_or3fft _04832_ (
    .a(_00353_),
    .b(_00354_),
    .c(_00352_),
    .y(_00355_)
  );
  al_ao21ttf _04833_ (
    .a(_00353_),
    .b(_00354_),
    .c(_00352_),
    .y(_00356_)
  );
  al_ao21ttf _04834_ (
    .a(TM0),
    .b(\DFF_25.Q ),
    .c(\DFF_153.Q ),
    .y(_00357_)
  );
  al_and3ftt _04835_ (
    .a(\DFF_153.Q ),
    .b(TM0),
    .c(\DFF_25.Q ),
    .y(_00358_)
  );
  al_and2ft _04836_ (
    .a(_00358_),
    .b(_00357_),
    .y(_00359_)
  );
  al_nand3ftt _04837_ (
    .a(_00359_),
    .b(_00356_),
    .c(_00355_),
    .y(_00360_)
  );
  al_ao21 _04838_ (
    .a(_00353_),
    .b(_00354_),
    .c(_00352_),
    .y(_00361_)
  );
  al_nand3 _04839_ (
    .a(_00353_),
    .b(_00354_),
    .c(_00352_),
    .y(_00362_)
  );
  al_nand3 _04840_ (
    .a(_00359_),
    .b(_00362_),
    .c(_00361_),
    .y(_00363_)
  );
  al_and2 _04841_ (
    .a(_00363_),
    .b(_00360_),
    .y(DATA_9_6)
  );
  al_and2ft _04842_ (
    .a(\DFF_90.Q ),
    .b(\DFF_122.Q ),
    .y(_00364_)
  );
  al_and2ft _04843_ (
    .a(\DFF_122.Q ),
    .b(\DFF_90.Q ),
    .y(_00365_)
  );
  al_or2 _04844_ (
    .a(_00364_),
    .b(_00365_),
    .y(_00366_)
  );
  al_nand2ft _04845_ (
    .a(\DFF_58.Q ),
    .b(TM0),
    .y(_00367_)
  );
  al_nand2ft _04846_ (
    .a(TM0),
    .b(\DFF_58.Q ),
    .y(_00368_)
  );
  al_or3fft _04847_ (
    .a(_00367_),
    .b(_00368_),
    .c(_00366_),
    .y(_00369_)
  );
  al_ao21ttf _04848_ (
    .a(_00367_),
    .b(_00368_),
    .c(_00366_),
    .y(_00370_)
  );
  al_ao21ttf _04849_ (
    .a(TM0),
    .b(\DFF_26.Q ),
    .c(\DFF_154.Q ),
    .y(_00371_)
  );
  al_and3ftt _04850_ (
    .a(\DFF_154.Q ),
    .b(TM0),
    .c(\DFF_26.Q ),
    .y(_00372_)
  );
  al_and2ft _04851_ (
    .a(_00372_),
    .b(_00371_),
    .y(_00373_)
  );
  al_nand3ftt _04852_ (
    .a(_00373_),
    .b(_00370_),
    .c(_00369_),
    .y(_00374_)
  );
  al_ao21 _04853_ (
    .a(_00367_),
    .b(_00368_),
    .c(_00366_),
    .y(_00375_)
  );
  al_nand3 _04854_ (
    .a(_00367_),
    .b(_00368_),
    .c(_00366_),
    .y(_00376_)
  );
  al_nand3 _04855_ (
    .a(_00373_),
    .b(_00376_),
    .c(_00375_),
    .y(_00377_)
  );
  al_and2 _04856_ (
    .a(_00377_),
    .b(_00374_),
    .y(DATA_9_5)
  );
  al_and2ft _04857_ (
    .a(\DFF_91.Q ),
    .b(\DFF_123.Q ),
    .y(_00378_)
  );
  al_and2ft _04858_ (
    .a(\DFF_123.Q ),
    .b(\DFF_91.Q ),
    .y(_00379_)
  );
  al_or2 _04859_ (
    .a(_00378_),
    .b(_00379_),
    .y(_00380_)
  );
  al_nand2ft _04860_ (
    .a(\DFF_59.Q ),
    .b(TM0),
    .y(_00381_)
  );
  al_nand2ft _04861_ (
    .a(TM0),
    .b(\DFF_59.Q ),
    .y(_00382_)
  );
  al_or3fft _04862_ (
    .a(_00381_),
    .b(_00382_),
    .c(_00380_),
    .y(_00383_)
  );
  al_ao21ttf _04863_ (
    .a(_00381_),
    .b(_00382_),
    .c(_00380_),
    .y(_00384_)
  );
  al_ao21ttf _04864_ (
    .a(TM0),
    .b(\DFF_27.Q ),
    .c(\DFF_155.Q ),
    .y(_00385_)
  );
  al_and3ftt _04865_ (
    .a(\DFF_155.Q ),
    .b(TM0),
    .c(\DFF_27.Q ),
    .y(_00386_)
  );
  al_and2ft _04866_ (
    .a(_00386_),
    .b(_00385_),
    .y(_00387_)
  );
  al_nand3ftt _04867_ (
    .a(_00387_),
    .b(_00384_),
    .c(_00383_),
    .y(_00388_)
  );
  al_ao21 _04868_ (
    .a(_00381_),
    .b(_00382_),
    .c(_00380_),
    .y(_00389_)
  );
  al_nand3 _04869_ (
    .a(_00381_),
    .b(_00382_),
    .c(_00380_),
    .y(_00390_)
  );
  al_nand3 _04870_ (
    .a(_00387_),
    .b(_00390_),
    .c(_00389_),
    .y(_00391_)
  );
  al_and2 _04871_ (
    .a(_00391_),
    .b(_00388_),
    .y(DATA_9_4)
  );
  al_and2ft _04872_ (
    .a(\DFF_92.Q ),
    .b(\DFF_124.Q ),
    .y(_00392_)
  );
  al_and2ft _04873_ (
    .a(\DFF_124.Q ),
    .b(\DFF_92.Q ),
    .y(_00393_)
  );
  al_or2 _04874_ (
    .a(_00392_),
    .b(_00393_),
    .y(_00394_)
  );
  al_nand2ft _04875_ (
    .a(\DFF_60.Q ),
    .b(TM0),
    .y(_00395_)
  );
  al_nand2ft _04876_ (
    .a(TM0),
    .b(\DFF_60.Q ),
    .y(_00396_)
  );
  al_or3fft _04877_ (
    .a(_00395_),
    .b(_00396_),
    .c(_00394_),
    .y(_00397_)
  );
  al_ao21ttf _04878_ (
    .a(_00395_),
    .b(_00396_),
    .c(_00394_),
    .y(_00398_)
  );
  al_ao21ttf _04879_ (
    .a(TM0),
    .b(\DFF_28.Q ),
    .c(\DFF_156.Q ),
    .y(_00399_)
  );
  al_and3ftt _04880_ (
    .a(\DFF_156.Q ),
    .b(TM0),
    .c(\DFF_28.Q ),
    .y(_00400_)
  );
  al_and2ft _04881_ (
    .a(_00400_),
    .b(_00399_),
    .y(_00401_)
  );
  al_nand3ftt _04882_ (
    .a(_00401_),
    .b(_00398_),
    .c(_00397_),
    .y(_00402_)
  );
  al_ao21 _04883_ (
    .a(_00395_),
    .b(_00396_),
    .c(_00394_),
    .y(_00403_)
  );
  al_nand3 _04884_ (
    .a(_00395_),
    .b(_00396_),
    .c(_00394_),
    .y(_00404_)
  );
  al_nand3 _04885_ (
    .a(_00401_),
    .b(_00404_),
    .c(_00403_),
    .y(_00405_)
  );
  al_and2 _04886_ (
    .a(_00405_),
    .b(_00402_),
    .y(DATA_9_3)
  );
  al_and2ft _04887_ (
    .a(\DFF_93.Q ),
    .b(\DFF_125.Q ),
    .y(_00406_)
  );
  al_and2ft _04888_ (
    .a(\DFF_125.Q ),
    .b(\DFF_93.Q ),
    .y(_00407_)
  );
  al_or2 _04889_ (
    .a(_00406_),
    .b(_00407_),
    .y(_00408_)
  );
  al_nand2ft _04890_ (
    .a(\DFF_61.Q ),
    .b(TM0),
    .y(_00409_)
  );
  al_nand2ft _04891_ (
    .a(TM0),
    .b(\DFF_61.Q ),
    .y(_00410_)
  );
  al_or3fft _04892_ (
    .a(_00409_),
    .b(_00410_),
    .c(_00408_),
    .y(_00411_)
  );
  al_ao21ttf _04893_ (
    .a(_00409_),
    .b(_00410_),
    .c(_00408_),
    .y(_00412_)
  );
  al_ao21ttf _04894_ (
    .a(TM0),
    .b(\DFF_29.Q ),
    .c(\DFF_157.Q ),
    .y(_00413_)
  );
  al_and3ftt _04895_ (
    .a(\DFF_157.Q ),
    .b(TM0),
    .c(\DFF_29.Q ),
    .y(_00414_)
  );
  al_and2ft _04896_ (
    .a(_00414_),
    .b(_00413_),
    .y(_00415_)
  );
  al_nand3ftt _04897_ (
    .a(_00415_),
    .b(_00412_),
    .c(_00411_),
    .y(_00416_)
  );
  al_ao21 _04898_ (
    .a(_00409_),
    .b(_00410_),
    .c(_00408_),
    .y(_00417_)
  );
  al_nand3 _04899_ (
    .a(_00409_),
    .b(_00410_),
    .c(_00408_),
    .y(_00418_)
  );
  al_nand3 _04900_ (
    .a(_00415_),
    .b(_00418_),
    .c(_00417_),
    .y(_00419_)
  );
  al_and2 _04901_ (
    .a(_00419_),
    .b(_00416_),
    .y(DATA_9_2)
  );
  al_and2ft _04902_ (
    .a(\DFF_94.Q ),
    .b(\DFF_126.Q ),
    .y(_00420_)
  );
  al_and2ft _04903_ (
    .a(\DFF_126.Q ),
    .b(\DFF_94.Q ),
    .y(_00421_)
  );
  al_or2 _04904_ (
    .a(_00420_),
    .b(_00421_),
    .y(_00422_)
  );
  al_nand2ft _04905_ (
    .a(\DFF_62.Q ),
    .b(TM0),
    .y(_00423_)
  );
  al_nand2ft _04906_ (
    .a(TM0),
    .b(\DFF_62.Q ),
    .y(_00424_)
  );
  al_or3fft _04907_ (
    .a(_00423_),
    .b(_00424_),
    .c(_00422_),
    .y(_00425_)
  );
  al_ao21ttf _04908_ (
    .a(_00423_),
    .b(_00424_),
    .c(_00422_),
    .y(_00426_)
  );
  al_ao21ttf _04909_ (
    .a(TM0),
    .b(\DFF_30.Q ),
    .c(\DFF_158.Q ),
    .y(_00427_)
  );
  al_and3ftt _04910_ (
    .a(\DFF_158.Q ),
    .b(TM0),
    .c(\DFF_30.Q ),
    .y(_00428_)
  );
  al_and2ft _04911_ (
    .a(_00428_),
    .b(_00427_),
    .y(_00429_)
  );
  al_nand3ftt _04912_ (
    .a(_00429_),
    .b(_00426_),
    .c(_00425_),
    .y(_00430_)
  );
  al_ao21 _04913_ (
    .a(_00423_),
    .b(_00424_),
    .c(_00422_),
    .y(_00431_)
  );
  al_nand3 _04914_ (
    .a(_00423_),
    .b(_00424_),
    .c(_00422_),
    .y(_00432_)
  );
  al_nand3 _04915_ (
    .a(_00429_),
    .b(_00432_),
    .c(_00431_),
    .y(_00433_)
  );
  al_and2 _04916_ (
    .a(_00433_),
    .b(_00430_),
    .y(DATA_9_1)
  );
  al_and2ft _04917_ (
    .a(\DFF_95.Q ),
    .b(\DFF_127.Q ),
    .y(_00434_)
  );
  al_and2ft _04918_ (
    .a(\DFF_127.Q ),
    .b(\DFF_95.Q ),
    .y(_00435_)
  );
  al_or2 _04919_ (
    .a(_00434_),
    .b(_00435_),
    .y(_00436_)
  );
  al_nand2ft _04920_ (
    .a(\DFF_63.Q ),
    .b(TM0),
    .y(_00437_)
  );
  al_nand2ft _04921_ (
    .a(TM0),
    .b(\DFF_63.Q ),
    .y(_00438_)
  );
  al_or3fft _04922_ (
    .a(_00437_),
    .b(_00438_),
    .c(_00436_),
    .y(_00439_)
  );
  al_ao21ttf _04923_ (
    .a(_00437_),
    .b(_00438_),
    .c(_00436_),
    .y(_00440_)
  );
  al_ao21ttf _04924_ (
    .a(TM0),
    .b(\DFF_31.Q ),
    .c(\DFF_159.Q ),
    .y(_00441_)
  );
  al_and3ftt _04925_ (
    .a(\DFF_159.Q ),
    .b(TM0),
    .c(\DFF_31.Q ),
    .y(_00442_)
  );
  al_and2ft _04926_ (
    .a(_00442_),
    .b(_00441_),
    .y(_00443_)
  );
  al_nand3ftt _04927_ (
    .a(_00443_),
    .b(_00440_),
    .c(_00439_),
    .y(_00444_)
  );
  al_ao21 _04928_ (
    .a(_00437_),
    .b(_00438_),
    .c(_00436_),
    .y(_00445_)
  );
  al_nand3 _04929_ (
    .a(_00437_),
    .b(_00438_),
    .c(_00436_),
    .y(_00446_)
  );
  al_nand3 _04930_ (
    .a(_00443_),
    .b(_00446_),
    .c(_00445_),
    .y(_00447_)
  );
  al_and2 _04931_ (
    .a(_00447_),
    .b(_00444_),
    .y(DATA_9_0)
  );
  al_and2 _04932_ (
    .a(\DFF_1.Q ),
    .b(RESET),
    .y(\DFF_0.D )
  );
  al_and2 _04933_ (
    .a(\DFF_2.Q ),
    .b(RESET),
    .y(\DFF_1.D )
  );
  al_and2 _04934_ (
    .a(\DFF_3.Q ),
    .b(RESET),
    .y(\DFF_2.D )
  );
  al_and2 _04935_ (
    .a(\DFF_4.Q ),
    .b(RESET),
    .y(\DFF_3.D )
  );
  al_and2 _04936_ (
    .a(\DFF_5.Q ),
    .b(RESET),
    .y(\DFF_4.D )
  );
  al_and2 _04937_ (
    .a(\DFF_6.Q ),
    .b(RESET),
    .y(\DFF_5.D )
  );
  al_and2 _04938_ (
    .a(\DFF_7.Q ),
    .b(RESET),
    .y(\DFF_6.D )
  );
  al_and2 _04939_ (
    .a(\DFF_8.Q ),
    .b(RESET),
    .y(\DFF_7.D )
  );
  al_and2 _04940_ (
    .a(\DFF_9.Q ),
    .b(RESET),
    .y(\DFF_8.D )
  );
  al_and2 _04941_ (
    .a(\DFF_10.Q ),
    .b(RESET),
    .y(\DFF_9.D )
  );
  al_and2 _04942_ (
    .a(\DFF_11.Q ),
    .b(RESET),
    .y(\DFF_10.D )
  );
  al_and2 _04943_ (
    .a(\DFF_12.Q ),
    .b(RESET),
    .y(\DFF_11.D )
  );
  al_and2 _04944_ (
    .a(\DFF_13.Q ),
    .b(RESET),
    .y(\DFF_12.D )
  );
  al_and2 _04945_ (
    .a(\DFF_14.Q ),
    .b(RESET),
    .y(\DFF_13.D )
  );
  al_and2 _04946_ (
    .a(\DFF_15.Q ),
    .b(RESET),
    .y(\DFF_14.D )
  );
  al_and2 _04947_ (
    .a(\DFF_16.Q ),
    .b(RESET),
    .y(\DFF_15.D )
  );
  al_and2 _04948_ (
    .a(\DFF_17.Q ),
    .b(RESET),
    .y(\DFF_16.D )
  );
  al_and2 _04949_ (
    .a(\DFF_18.Q ),
    .b(RESET),
    .y(\DFF_17.D )
  );
  al_and2 _04950_ (
    .a(\DFF_19.Q ),
    .b(RESET),
    .y(\DFF_18.D )
  );
  al_and2 _04951_ (
    .a(\DFF_20.Q ),
    .b(RESET),
    .y(\DFF_19.D )
  );
  al_and2 _04952_ (
    .a(\DFF_21.Q ),
    .b(RESET),
    .y(\DFF_20.D )
  );
  al_and2 _04953_ (
    .a(\DFF_22.Q ),
    .b(RESET),
    .y(\DFF_21.D )
  );
  al_and2 _04954_ (
    .a(\DFF_23.Q ),
    .b(RESET),
    .y(\DFF_22.D )
  );
  al_and2 _04955_ (
    .a(\DFF_24.Q ),
    .b(RESET),
    .y(\DFF_23.D )
  );
  al_and2 _04956_ (
    .a(\DFF_25.Q ),
    .b(RESET),
    .y(\DFF_24.D )
  );
  al_and2 _04957_ (
    .a(\DFF_26.Q ),
    .b(RESET),
    .y(\DFF_25.D )
  );
  al_and2 _04958_ (
    .a(\DFF_27.Q ),
    .b(RESET),
    .y(\DFF_26.D )
  );
  al_and2 _04959_ (
    .a(\DFF_28.Q ),
    .b(RESET),
    .y(\DFF_27.D )
  );
  al_and2 _04960_ (
    .a(\DFF_29.Q ),
    .b(RESET),
    .y(\DFF_28.D )
  );
  al_and2 _04961_ (
    .a(\DFF_30.Q ),
    .b(RESET),
    .y(\DFF_29.D )
  );
  al_and2 _04962_ (
    .a(\DFF_31.Q ),
    .b(RESET),
    .y(\DFF_30.D )
  );
  al_and2ft _04963_ (
    .a(\DFF_0.Q ),
    .b(RESET),
    .y(\DFF_31.D )
  );
  al_inv _04964_ (
    .a(TM0),
    .y(_00448_)
  );
  al_nand3 _04965_ (
    .a(_00448_),
    .b(_00013_),
    .c(_00010_),
    .y(_00449_)
  );
  al_ao21ttf _04966_ (
    .a(\DFF_0.Q ),
    .b(TM0),
    .c(TM1),
    .y(_00450_)
  );
  al_inv _04967_ (
    .a(RESET),
    .y(_00451_)
  );
  al_or2 _04968_ (
    .a(TM1),
    .b(\DFF_288.Q ),
    .y(_00452_)
  );
  al_nand2 _04969_ (
    .a(TM1),
    .b(\DFF_288.Q ),
    .y(_00453_)
  );
  al_nand3 _04970_ (
    .a(\DFF_320.Q ),
    .b(_00452_),
    .c(_00453_),
    .y(_00454_)
  );
  al_nand2ft _04971_ (
    .a(TM1),
    .b(\DFF_288.Q ),
    .y(_00455_)
  );
  al_nand2ft _04972_ (
    .a(\DFF_288.Q ),
    .b(TM1),
    .y(_00456_)
  );
  al_nand3ftt _04973_ (
    .a(\DFF_320.Q ),
    .b(_00455_),
    .c(_00456_),
    .y(_00457_)
  );
  al_and2ft _04974_ (
    .a(\DFF_256.Q ),
    .b(\DFF_224.Q ),
    .y(_00458_)
  );
  al_nand2ft _04975_ (
    .a(\DFF_224.Q ),
    .b(\DFF_256.Q ),
    .y(_00459_)
  );
  al_nand2ft _04976_ (
    .a(_00458_),
    .b(_00459_),
    .y(_00460_)
  );
  al_ao21 _04977_ (
    .a(_00457_),
    .b(_00454_),
    .c(_00460_),
    .y(_00461_)
  );
  al_nand3 _04978_ (
    .a(_00457_),
    .b(_00454_),
    .c(_00460_),
    .y(_00462_)
  );
  al_nand3 _04979_ (
    .a(_00448_),
    .b(_00461_),
    .c(_00462_),
    .y(_00463_)
  );
  al_aoi21 _04980_ (
    .a(TM0),
    .b(\DFF_191.Q ),
    .c(TM1),
    .y(_00464_)
  );
  al_aoi21 _04981_ (
    .a(_00464_),
    .b(_00463_),
    .c(_00451_),
    .y(_00465_)
  );
  al_aoi21ftf _04982_ (
    .a(_00450_),
    .b(_00449_),
    .c(_00465_),
    .y(\DFF_32.D )
  );
  al_nand3 _04983_ (
    .a(_00448_),
    .b(_00027_),
    .c(_00024_),
    .y(_00466_)
  );
  al_ao21ttf _04984_ (
    .a(TM0),
    .b(\DFF_1.Q ),
    .c(TM1),
    .y(_00467_)
  );
  al_or2 _04985_ (
    .a(TM1),
    .b(\DFF_289.Q ),
    .y(_00468_)
  );
  al_nand2 _04986_ (
    .a(TM1),
    .b(\DFF_289.Q ),
    .y(_00469_)
  );
  al_nand3 _04987_ (
    .a(\DFF_321.Q ),
    .b(_00468_),
    .c(_00469_),
    .y(_00470_)
  );
  al_nand2ft _04988_ (
    .a(TM1),
    .b(\DFF_289.Q ),
    .y(_00471_)
  );
  al_nand2ft _04989_ (
    .a(\DFF_289.Q ),
    .b(TM1),
    .y(_00472_)
  );
  al_nand3ftt _04990_ (
    .a(\DFF_321.Q ),
    .b(_00471_),
    .c(_00472_),
    .y(_00473_)
  );
  al_and2ft _04991_ (
    .a(\DFF_257.Q ),
    .b(\DFF_225.Q ),
    .y(_00474_)
  );
  al_nand2ft _04992_ (
    .a(\DFF_225.Q ),
    .b(\DFF_257.Q ),
    .y(_00475_)
  );
  al_nand2ft _04993_ (
    .a(_00474_),
    .b(_00475_),
    .y(_00476_)
  );
  al_ao21 _04994_ (
    .a(_00473_),
    .b(_00470_),
    .c(_00476_),
    .y(_00477_)
  );
  al_nand3 _04995_ (
    .a(_00473_),
    .b(_00470_),
    .c(_00476_),
    .y(_00478_)
  );
  al_nand3 _04996_ (
    .a(_00448_),
    .b(_00477_),
    .c(_00478_),
    .y(_00479_)
  );
  al_aoi21 _04997_ (
    .a(TM0),
    .b(\DFF_190.Q ),
    .c(TM1),
    .y(_00480_)
  );
  al_aoi21 _04998_ (
    .a(_00480_),
    .b(_00479_),
    .c(_00451_),
    .y(_00481_)
  );
  al_aoi21ftf _04999_ (
    .a(_00467_),
    .b(_00466_),
    .c(_00481_),
    .y(\DFF_33.D )
  );
  al_nand3 _05000_ (
    .a(_00448_),
    .b(_00041_),
    .c(_00038_),
    .y(_00482_)
  );
  al_ao21ttf _05001_ (
    .a(TM0),
    .b(\DFF_2.Q ),
    .c(TM1),
    .y(_00483_)
  );
  al_or2 _05002_ (
    .a(TM1),
    .b(\DFF_290.Q ),
    .y(_00484_)
  );
  al_nand2 _05003_ (
    .a(TM1),
    .b(\DFF_290.Q ),
    .y(_00485_)
  );
  al_nand3 _05004_ (
    .a(\DFF_322.Q ),
    .b(_00484_),
    .c(_00485_),
    .y(_00486_)
  );
  al_nand2ft _05005_ (
    .a(TM1),
    .b(\DFF_290.Q ),
    .y(_00487_)
  );
  al_nand2ft _05006_ (
    .a(\DFF_290.Q ),
    .b(TM1),
    .y(_00488_)
  );
  al_nand3ftt _05007_ (
    .a(\DFF_322.Q ),
    .b(_00487_),
    .c(_00488_),
    .y(_00489_)
  );
  al_and2ft _05008_ (
    .a(\DFF_258.Q ),
    .b(\DFF_226.Q ),
    .y(_00490_)
  );
  al_nand2ft _05009_ (
    .a(\DFF_226.Q ),
    .b(\DFF_258.Q ),
    .y(_00491_)
  );
  al_nand2ft _05010_ (
    .a(_00490_),
    .b(_00491_),
    .y(_00492_)
  );
  al_ao21 _05011_ (
    .a(_00489_),
    .b(_00486_),
    .c(_00492_),
    .y(_00493_)
  );
  al_nand3 _05012_ (
    .a(_00489_),
    .b(_00486_),
    .c(_00492_),
    .y(_00494_)
  );
  al_nand3 _05013_ (
    .a(_00448_),
    .b(_00493_),
    .c(_00494_),
    .y(_00495_)
  );
  al_aoi21 _05014_ (
    .a(TM0),
    .b(\DFF_189.Q ),
    .c(TM1),
    .y(_00496_)
  );
  al_aoi21 _05015_ (
    .a(_00496_),
    .b(_00495_),
    .c(_00451_),
    .y(_00497_)
  );
  al_aoi21ftf _05016_ (
    .a(_00483_),
    .b(_00482_),
    .c(_00497_),
    .y(\DFF_34.D )
  );
  al_nand3 _05017_ (
    .a(_00448_),
    .b(_00055_),
    .c(_00052_),
    .y(_00498_)
  );
  al_ao21ttf _05018_ (
    .a(TM0),
    .b(\DFF_3.Q ),
    .c(TM1),
    .y(_00499_)
  );
  al_or2 _05019_ (
    .a(TM1),
    .b(\DFF_291.Q ),
    .y(_00500_)
  );
  al_nand2 _05020_ (
    .a(TM1),
    .b(\DFF_291.Q ),
    .y(_00501_)
  );
  al_nand3 _05021_ (
    .a(\DFF_323.Q ),
    .b(_00500_),
    .c(_00501_),
    .y(_00502_)
  );
  al_nand2ft _05022_ (
    .a(TM1),
    .b(\DFF_291.Q ),
    .y(_00503_)
  );
  al_nand2ft _05023_ (
    .a(\DFF_291.Q ),
    .b(TM1),
    .y(_00504_)
  );
  al_nand3ftt _05024_ (
    .a(\DFF_323.Q ),
    .b(_00503_),
    .c(_00504_),
    .y(_00505_)
  );
  al_and2ft _05025_ (
    .a(\DFF_259.Q ),
    .b(\DFF_227.Q ),
    .y(_00506_)
  );
  al_nand2ft _05026_ (
    .a(\DFF_227.Q ),
    .b(\DFF_259.Q ),
    .y(_00507_)
  );
  al_nand2ft _05027_ (
    .a(_00506_),
    .b(_00507_),
    .y(_00508_)
  );
  al_ao21 _05028_ (
    .a(_00505_),
    .b(_00502_),
    .c(_00508_),
    .y(_00509_)
  );
  al_nand3 _05029_ (
    .a(_00505_),
    .b(_00502_),
    .c(_00508_),
    .y(_00510_)
  );
  al_nand3 _05030_ (
    .a(_00448_),
    .b(_00509_),
    .c(_00510_),
    .y(_00511_)
  );
  al_aoi21 _05031_ (
    .a(TM0),
    .b(\DFF_188.Q ),
    .c(TM1),
    .y(_00512_)
  );
  al_aoi21 _05032_ (
    .a(_00512_),
    .b(_00511_),
    .c(_00451_),
    .y(_00513_)
  );
  al_aoi21ftf _05033_ (
    .a(_00499_),
    .b(_00498_),
    .c(_00513_),
    .y(\DFF_35.D )
  );
  al_nand3 _05034_ (
    .a(_00448_),
    .b(_00069_),
    .c(_00066_),
    .y(_00514_)
  );
  al_ao21ttf _05035_ (
    .a(TM0),
    .b(\DFF_4.Q ),
    .c(TM1),
    .y(_00515_)
  );
  al_or2 _05036_ (
    .a(TM1),
    .b(\DFF_292.Q ),
    .y(_00516_)
  );
  al_nand2 _05037_ (
    .a(TM1),
    .b(\DFF_292.Q ),
    .y(_00517_)
  );
  al_nand3 _05038_ (
    .a(\DFF_324.Q ),
    .b(_00516_),
    .c(_00517_),
    .y(_00518_)
  );
  al_nand2ft _05039_ (
    .a(TM1),
    .b(\DFF_292.Q ),
    .y(_00519_)
  );
  al_nand2ft _05040_ (
    .a(\DFF_292.Q ),
    .b(TM1),
    .y(_00520_)
  );
  al_nand3ftt _05041_ (
    .a(\DFF_324.Q ),
    .b(_00519_),
    .c(_00520_),
    .y(_00521_)
  );
  al_and2ft _05042_ (
    .a(\DFF_260.Q ),
    .b(\DFF_228.Q ),
    .y(_00522_)
  );
  al_nand2ft _05043_ (
    .a(\DFF_228.Q ),
    .b(\DFF_260.Q ),
    .y(_00523_)
  );
  al_nand2ft _05044_ (
    .a(_00522_),
    .b(_00523_),
    .y(_00524_)
  );
  al_ao21 _05045_ (
    .a(_00521_),
    .b(_00518_),
    .c(_00524_),
    .y(_00525_)
  );
  al_nand3 _05046_ (
    .a(_00521_),
    .b(_00518_),
    .c(_00524_),
    .y(_00526_)
  );
  al_nand3 _05047_ (
    .a(_00448_),
    .b(_00525_),
    .c(_00526_),
    .y(_00527_)
  );
  al_aoi21 _05048_ (
    .a(TM0),
    .b(\DFF_187.Q ),
    .c(TM1),
    .y(_00528_)
  );
  al_aoi21 _05049_ (
    .a(_00528_),
    .b(_00527_),
    .c(_00451_),
    .y(_00529_)
  );
  al_aoi21ftf _05050_ (
    .a(_00515_),
    .b(_00514_),
    .c(_00529_),
    .y(\DFF_36.D )
  );
  al_nand3 _05051_ (
    .a(_00448_),
    .b(_00083_),
    .c(_00080_),
    .y(_00530_)
  );
  al_ao21ttf _05052_ (
    .a(TM0),
    .b(\DFF_5.Q ),
    .c(TM1),
    .y(_00531_)
  );
  al_or2 _05053_ (
    .a(TM1),
    .b(\DFF_293.Q ),
    .y(_00532_)
  );
  al_nand2 _05054_ (
    .a(TM1),
    .b(\DFF_293.Q ),
    .y(_00533_)
  );
  al_nand3 _05055_ (
    .a(\DFF_325.Q ),
    .b(_00532_),
    .c(_00533_),
    .y(_00534_)
  );
  al_nand2ft _05056_ (
    .a(TM1),
    .b(\DFF_293.Q ),
    .y(_00535_)
  );
  al_nand2ft _05057_ (
    .a(\DFF_293.Q ),
    .b(TM1),
    .y(_00536_)
  );
  al_nand3ftt _05058_ (
    .a(\DFF_325.Q ),
    .b(_00535_),
    .c(_00536_),
    .y(_00537_)
  );
  al_and2ft _05059_ (
    .a(\DFF_261.Q ),
    .b(\DFF_229.Q ),
    .y(_00538_)
  );
  al_nand2ft _05060_ (
    .a(\DFF_229.Q ),
    .b(\DFF_261.Q ),
    .y(_00539_)
  );
  al_nand2ft _05061_ (
    .a(_00538_),
    .b(_00539_),
    .y(_00540_)
  );
  al_ao21 _05062_ (
    .a(_00537_),
    .b(_00534_),
    .c(_00540_),
    .y(_00541_)
  );
  al_nand3 _05063_ (
    .a(_00537_),
    .b(_00534_),
    .c(_00540_),
    .y(_00542_)
  );
  al_nand3 _05064_ (
    .a(_00448_),
    .b(_00541_),
    .c(_00542_),
    .y(_00543_)
  );
  al_aoi21 _05065_ (
    .a(TM0),
    .b(\DFF_186.Q ),
    .c(TM1),
    .y(_00544_)
  );
  al_aoi21 _05066_ (
    .a(_00544_),
    .b(_00543_),
    .c(_00451_),
    .y(_00545_)
  );
  al_aoi21ftf _05067_ (
    .a(_00531_),
    .b(_00530_),
    .c(_00545_),
    .y(\DFF_37.D )
  );
  al_nand3 _05068_ (
    .a(_00448_),
    .b(_00097_),
    .c(_00094_),
    .y(_00546_)
  );
  al_ao21ttf _05069_ (
    .a(TM0),
    .b(\DFF_6.Q ),
    .c(TM1),
    .y(_00547_)
  );
  al_or2 _05070_ (
    .a(TM1),
    .b(\DFF_294.Q ),
    .y(_00548_)
  );
  al_nand2 _05071_ (
    .a(TM1),
    .b(\DFF_294.Q ),
    .y(_00549_)
  );
  al_nand3 _05072_ (
    .a(\DFF_326.Q ),
    .b(_00548_),
    .c(_00549_),
    .y(_00550_)
  );
  al_nand2ft _05073_ (
    .a(TM1),
    .b(\DFF_294.Q ),
    .y(_00551_)
  );
  al_nand2ft _05074_ (
    .a(\DFF_294.Q ),
    .b(TM1),
    .y(_00552_)
  );
  al_nand3ftt _05075_ (
    .a(\DFF_326.Q ),
    .b(_00551_),
    .c(_00552_),
    .y(_00553_)
  );
  al_and2ft _05076_ (
    .a(\DFF_262.Q ),
    .b(\DFF_230.Q ),
    .y(_00554_)
  );
  al_nand2ft _05077_ (
    .a(\DFF_230.Q ),
    .b(\DFF_262.Q ),
    .y(_00555_)
  );
  al_nand2ft _05078_ (
    .a(_00554_),
    .b(_00555_),
    .y(_00556_)
  );
  al_ao21 _05079_ (
    .a(_00553_),
    .b(_00550_),
    .c(_00556_),
    .y(_00557_)
  );
  al_nand3 _05080_ (
    .a(_00553_),
    .b(_00550_),
    .c(_00556_),
    .y(_00558_)
  );
  al_nand3 _05081_ (
    .a(_00448_),
    .b(_00557_),
    .c(_00558_),
    .y(_00559_)
  );
  al_aoi21 _05082_ (
    .a(TM0),
    .b(\DFF_185.Q ),
    .c(TM1),
    .y(_00560_)
  );
  al_aoi21 _05083_ (
    .a(_00560_),
    .b(_00559_),
    .c(_00451_),
    .y(_00561_)
  );
  al_aoi21ftf _05084_ (
    .a(_00547_),
    .b(_00546_),
    .c(_00561_),
    .y(\DFF_38.D )
  );
  al_nand3 _05085_ (
    .a(_00448_),
    .b(_00111_),
    .c(_00108_),
    .y(_00562_)
  );
  al_ao21ttf _05086_ (
    .a(TM0),
    .b(\DFF_7.Q ),
    .c(TM1),
    .y(_00563_)
  );
  al_or2 _05087_ (
    .a(TM1),
    .b(\DFF_295.Q ),
    .y(_00564_)
  );
  al_nand2 _05088_ (
    .a(TM1),
    .b(\DFF_295.Q ),
    .y(_00565_)
  );
  al_nand3 _05089_ (
    .a(\DFF_327.Q ),
    .b(_00564_),
    .c(_00565_),
    .y(_00566_)
  );
  al_nand2ft _05090_ (
    .a(TM1),
    .b(\DFF_295.Q ),
    .y(_00567_)
  );
  al_nand2ft _05091_ (
    .a(\DFF_295.Q ),
    .b(TM1),
    .y(_00568_)
  );
  al_nand3ftt _05092_ (
    .a(\DFF_327.Q ),
    .b(_00567_),
    .c(_00568_),
    .y(_00569_)
  );
  al_and2ft _05093_ (
    .a(\DFF_263.Q ),
    .b(\DFF_231.Q ),
    .y(_00570_)
  );
  al_nand2ft _05094_ (
    .a(\DFF_231.Q ),
    .b(\DFF_263.Q ),
    .y(_00571_)
  );
  al_nand2ft _05095_ (
    .a(_00570_),
    .b(_00571_),
    .y(_00572_)
  );
  al_ao21 _05096_ (
    .a(_00569_),
    .b(_00566_),
    .c(_00572_),
    .y(_00573_)
  );
  al_nand3 _05097_ (
    .a(_00569_),
    .b(_00566_),
    .c(_00572_),
    .y(_00574_)
  );
  al_nand3 _05098_ (
    .a(_00448_),
    .b(_00573_),
    .c(_00574_),
    .y(_00575_)
  );
  al_aoi21 _05099_ (
    .a(TM0),
    .b(\DFF_184.Q ),
    .c(TM1),
    .y(_00576_)
  );
  al_aoi21 _05100_ (
    .a(_00576_),
    .b(_00575_),
    .c(_00451_),
    .y(_00577_)
  );
  al_aoi21ftf _05101_ (
    .a(_00563_),
    .b(_00562_),
    .c(_00577_),
    .y(\DFF_39.D )
  );
  al_nand3 _05102_ (
    .a(_00448_),
    .b(_00125_),
    .c(_00122_),
    .y(_00578_)
  );
  al_ao21ttf _05103_ (
    .a(TM0),
    .b(\DFF_8.Q ),
    .c(TM1),
    .y(_00579_)
  );
  al_or2 _05104_ (
    .a(TM1),
    .b(\DFF_296.Q ),
    .y(_00580_)
  );
  al_nand2 _05105_ (
    .a(TM1),
    .b(\DFF_296.Q ),
    .y(_00581_)
  );
  al_nand3 _05106_ (
    .a(\DFF_328.Q ),
    .b(_00580_),
    .c(_00581_),
    .y(_00582_)
  );
  al_nand2ft _05107_ (
    .a(TM1),
    .b(\DFF_296.Q ),
    .y(_00583_)
  );
  al_nand2ft _05108_ (
    .a(\DFF_296.Q ),
    .b(TM1),
    .y(_00584_)
  );
  al_nand3ftt _05109_ (
    .a(\DFF_328.Q ),
    .b(_00583_),
    .c(_00584_),
    .y(_00585_)
  );
  al_and2ft _05110_ (
    .a(\DFF_264.Q ),
    .b(\DFF_232.Q ),
    .y(_00586_)
  );
  al_nand2ft _05111_ (
    .a(\DFF_232.Q ),
    .b(\DFF_264.Q ),
    .y(_00587_)
  );
  al_nand2ft _05112_ (
    .a(_00586_),
    .b(_00587_),
    .y(_00588_)
  );
  al_ao21 _05113_ (
    .a(_00585_),
    .b(_00582_),
    .c(_00588_),
    .y(_00589_)
  );
  al_nand3 _05114_ (
    .a(_00585_),
    .b(_00582_),
    .c(_00588_),
    .y(_00590_)
  );
  al_nand3 _05115_ (
    .a(_00448_),
    .b(_00589_),
    .c(_00590_),
    .y(_00591_)
  );
  al_aoi21 _05116_ (
    .a(TM0),
    .b(\DFF_183.Q ),
    .c(TM1),
    .y(_00592_)
  );
  al_aoi21 _05117_ (
    .a(_00592_),
    .b(_00591_),
    .c(_00451_),
    .y(_00593_)
  );
  al_aoi21ftf _05118_ (
    .a(_00579_),
    .b(_00578_),
    .c(_00593_),
    .y(\DFF_40.D )
  );
  al_nand3 _05119_ (
    .a(_00448_),
    .b(_00139_),
    .c(_00136_),
    .y(_00594_)
  );
  al_ao21ttf _05120_ (
    .a(TM0),
    .b(\DFF_9.Q ),
    .c(TM1),
    .y(_00595_)
  );
  al_or2 _05121_ (
    .a(TM1),
    .b(\DFF_297.Q ),
    .y(_00596_)
  );
  al_nand2 _05122_ (
    .a(TM1),
    .b(\DFF_297.Q ),
    .y(_00597_)
  );
  al_nand3 _05123_ (
    .a(\DFF_329.Q ),
    .b(_00596_),
    .c(_00597_),
    .y(_00598_)
  );
  al_nand2ft _05124_ (
    .a(TM1),
    .b(\DFF_297.Q ),
    .y(_00599_)
  );
  al_nand2ft _05125_ (
    .a(\DFF_297.Q ),
    .b(TM1),
    .y(_00600_)
  );
  al_nand3ftt _05126_ (
    .a(\DFF_329.Q ),
    .b(_00599_),
    .c(_00600_),
    .y(_00601_)
  );
  al_and2ft _05127_ (
    .a(\DFF_265.Q ),
    .b(\DFF_233.Q ),
    .y(_00602_)
  );
  al_nand2ft _05128_ (
    .a(\DFF_233.Q ),
    .b(\DFF_265.Q ),
    .y(_00603_)
  );
  al_nand2ft _05129_ (
    .a(_00602_),
    .b(_00603_),
    .y(_00604_)
  );
  al_ao21 _05130_ (
    .a(_00601_),
    .b(_00598_),
    .c(_00604_),
    .y(_00605_)
  );
  al_nand3 _05131_ (
    .a(_00601_),
    .b(_00598_),
    .c(_00604_),
    .y(_00606_)
  );
  al_nand3 _05132_ (
    .a(_00448_),
    .b(_00605_),
    .c(_00606_),
    .y(_00607_)
  );
  al_aoi21 _05133_ (
    .a(TM0),
    .b(\DFF_182.Q ),
    .c(TM1),
    .y(_00608_)
  );
  al_aoi21 _05134_ (
    .a(_00608_),
    .b(_00607_),
    .c(_00451_),
    .y(_00609_)
  );
  al_aoi21ftf _05135_ (
    .a(_00595_),
    .b(_00594_),
    .c(_00609_),
    .y(\DFF_41.D )
  );
  al_nand3 _05136_ (
    .a(_00448_),
    .b(_00153_),
    .c(_00150_),
    .y(_00610_)
  );
  al_ao21ttf _05137_ (
    .a(TM0),
    .b(\DFF_10.Q ),
    .c(TM1),
    .y(_00611_)
  );
  al_or2 _05138_ (
    .a(TM1),
    .b(\DFF_298.Q ),
    .y(_00612_)
  );
  al_nand2 _05139_ (
    .a(TM1),
    .b(\DFF_298.Q ),
    .y(_00613_)
  );
  al_nand3 _05140_ (
    .a(\DFF_330.Q ),
    .b(_00612_),
    .c(_00613_),
    .y(_00614_)
  );
  al_nand2ft _05141_ (
    .a(TM1),
    .b(\DFF_298.Q ),
    .y(_00615_)
  );
  al_nand2ft _05142_ (
    .a(\DFF_298.Q ),
    .b(TM1),
    .y(_00616_)
  );
  al_nand3ftt _05143_ (
    .a(\DFF_330.Q ),
    .b(_00615_),
    .c(_00616_),
    .y(_00617_)
  );
  al_and2ft _05144_ (
    .a(\DFF_266.Q ),
    .b(\DFF_234.Q ),
    .y(_00618_)
  );
  al_nand2ft _05145_ (
    .a(\DFF_234.Q ),
    .b(\DFF_266.Q ),
    .y(_00619_)
  );
  al_nand2ft _05146_ (
    .a(_00618_),
    .b(_00619_),
    .y(_00620_)
  );
  al_ao21 _05147_ (
    .a(_00617_),
    .b(_00614_),
    .c(_00620_),
    .y(_00621_)
  );
  al_nand3 _05148_ (
    .a(_00617_),
    .b(_00614_),
    .c(_00620_),
    .y(_00622_)
  );
  al_nand3 _05149_ (
    .a(_00448_),
    .b(_00621_),
    .c(_00622_),
    .y(_00623_)
  );
  al_aoi21 _05150_ (
    .a(TM0),
    .b(\DFF_181.Q ),
    .c(TM1),
    .y(_00624_)
  );
  al_aoi21 _05151_ (
    .a(_00624_),
    .b(_00623_),
    .c(_00451_),
    .y(_00625_)
  );
  al_aoi21ftf _05152_ (
    .a(_00611_),
    .b(_00610_),
    .c(_00625_),
    .y(\DFF_42.D )
  );
  al_nand3 _05153_ (
    .a(_00448_),
    .b(_00167_),
    .c(_00164_),
    .y(_00626_)
  );
  al_ao21ttf _05154_ (
    .a(TM0),
    .b(\DFF_11.Q ),
    .c(TM1),
    .y(_00627_)
  );
  al_or2 _05155_ (
    .a(TM1),
    .b(\DFF_299.Q ),
    .y(_00628_)
  );
  al_nand2 _05156_ (
    .a(TM1),
    .b(\DFF_299.Q ),
    .y(_00629_)
  );
  al_nand3 _05157_ (
    .a(\DFF_331.Q ),
    .b(_00628_),
    .c(_00629_),
    .y(_00630_)
  );
  al_nand2ft _05158_ (
    .a(TM1),
    .b(\DFF_299.Q ),
    .y(_00631_)
  );
  al_nand2ft _05159_ (
    .a(\DFF_299.Q ),
    .b(TM1),
    .y(_00632_)
  );
  al_nand3ftt _05160_ (
    .a(\DFF_331.Q ),
    .b(_00631_),
    .c(_00632_),
    .y(_00633_)
  );
  al_and2ft _05161_ (
    .a(\DFF_267.Q ),
    .b(\DFF_235.Q ),
    .y(_00634_)
  );
  al_nand2ft _05162_ (
    .a(\DFF_235.Q ),
    .b(\DFF_267.Q ),
    .y(_00635_)
  );
  al_nand2ft _05163_ (
    .a(_00634_),
    .b(_00635_),
    .y(_00636_)
  );
  al_ao21 _05164_ (
    .a(_00633_),
    .b(_00630_),
    .c(_00636_),
    .y(_00637_)
  );
  al_nand3 _05165_ (
    .a(_00633_),
    .b(_00630_),
    .c(_00636_),
    .y(_00638_)
  );
  al_nand3 _05166_ (
    .a(_00448_),
    .b(_00637_),
    .c(_00638_),
    .y(_00639_)
  );
  al_aoi21 _05167_ (
    .a(TM0),
    .b(\DFF_180.Q ),
    .c(TM1),
    .y(_00640_)
  );
  al_aoi21 _05168_ (
    .a(_00640_),
    .b(_00639_),
    .c(_00451_),
    .y(_00641_)
  );
  al_aoi21ftf _05169_ (
    .a(_00627_),
    .b(_00626_),
    .c(_00641_),
    .y(\DFF_43.D )
  );
  al_nand3 _05170_ (
    .a(_00448_),
    .b(_00181_),
    .c(_00178_),
    .y(_00642_)
  );
  al_ao21ttf _05171_ (
    .a(TM0),
    .b(\DFF_12.Q ),
    .c(TM1),
    .y(_00643_)
  );
  al_or2 _05172_ (
    .a(TM1),
    .b(\DFF_300.Q ),
    .y(_00644_)
  );
  al_nand2 _05173_ (
    .a(TM1),
    .b(\DFF_300.Q ),
    .y(_00645_)
  );
  al_nand3 _05174_ (
    .a(\DFF_332.Q ),
    .b(_00644_),
    .c(_00645_),
    .y(_00646_)
  );
  al_nand2ft _05175_ (
    .a(TM1),
    .b(\DFF_300.Q ),
    .y(_00647_)
  );
  al_nand2ft _05176_ (
    .a(\DFF_300.Q ),
    .b(TM1),
    .y(_00648_)
  );
  al_nand3ftt _05177_ (
    .a(\DFF_332.Q ),
    .b(_00647_),
    .c(_00648_),
    .y(_00649_)
  );
  al_and2ft _05178_ (
    .a(\DFF_268.Q ),
    .b(\DFF_236.Q ),
    .y(_00650_)
  );
  al_nand2ft _05179_ (
    .a(\DFF_236.Q ),
    .b(\DFF_268.Q ),
    .y(_00651_)
  );
  al_nand2ft _05180_ (
    .a(_00650_),
    .b(_00651_),
    .y(_00652_)
  );
  al_ao21 _05181_ (
    .a(_00649_),
    .b(_00646_),
    .c(_00652_),
    .y(_00653_)
  );
  al_nand3 _05182_ (
    .a(_00649_),
    .b(_00646_),
    .c(_00652_),
    .y(_00654_)
  );
  al_nand3 _05183_ (
    .a(_00448_),
    .b(_00653_),
    .c(_00654_),
    .y(_00655_)
  );
  al_aoi21 _05184_ (
    .a(TM0),
    .b(\DFF_179.Q ),
    .c(TM1),
    .y(_00656_)
  );
  al_aoi21 _05185_ (
    .a(_00656_),
    .b(_00655_),
    .c(_00451_),
    .y(_00657_)
  );
  al_aoi21ftf _05186_ (
    .a(_00643_),
    .b(_00642_),
    .c(_00657_),
    .y(\DFF_44.D )
  );
  al_nand3 _05187_ (
    .a(_00448_),
    .b(_00195_),
    .c(_00192_),
    .y(_00658_)
  );
  al_ao21ttf _05188_ (
    .a(TM0),
    .b(\DFF_13.Q ),
    .c(TM1),
    .y(_00659_)
  );
  al_or2 _05189_ (
    .a(TM1),
    .b(\DFF_301.Q ),
    .y(_00660_)
  );
  al_nand2 _05190_ (
    .a(TM1),
    .b(\DFF_301.Q ),
    .y(_00661_)
  );
  al_nand3 _05191_ (
    .a(\DFF_333.Q ),
    .b(_00660_),
    .c(_00661_),
    .y(_00662_)
  );
  al_nand2ft _05192_ (
    .a(TM1),
    .b(\DFF_301.Q ),
    .y(_00663_)
  );
  al_nand2ft _05193_ (
    .a(\DFF_301.Q ),
    .b(TM1),
    .y(_00664_)
  );
  al_nand3ftt _05194_ (
    .a(\DFF_333.Q ),
    .b(_00663_),
    .c(_00664_),
    .y(_00665_)
  );
  al_and2ft _05195_ (
    .a(\DFF_269.Q ),
    .b(\DFF_237.Q ),
    .y(_00666_)
  );
  al_nand2ft _05196_ (
    .a(\DFF_237.Q ),
    .b(\DFF_269.Q ),
    .y(_00667_)
  );
  al_nand2ft _05197_ (
    .a(_00666_),
    .b(_00667_),
    .y(_00668_)
  );
  al_ao21 _05198_ (
    .a(_00665_),
    .b(_00662_),
    .c(_00668_),
    .y(_00669_)
  );
  al_nand3 _05199_ (
    .a(_00665_),
    .b(_00662_),
    .c(_00668_),
    .y(_00670_)
  );
  al_nand3 _05200_ (
    .a(_00448_),
    .b(_00669_),
    .c(_00670_),
    .y(_00671_)
  );
  al_aoi21 _05201_ (
    .a(TM0),
    .b(\DFF_178.Q ),
    .c(TM1),
    .y(_00672_)
  );
  al_aoi21 _05202_ (
    .a(_00672_),
    .b(_00671_),
    .c(_00451_),
    .y(_00673_)
  );
  al_aoi21ftf _05203_ (
    .a(_00659_),
    .b(_00658_),
    .c(_00673_),
    .y(\DFF_45.D )
  );
  al_nand3 _05204_ (
    .a(_00448_),
    .b(_00209_),
    .c(_00206_),
    .y(_00674_)
  );
  al_ao21ttf _05205_ (
    .a(TM0),
    .b(\DFF_14.Q ),
    .c(TM1),
    .y(_00675_)
  );
  al_or2 _05206_ (
    .a(TM1),
    .b(\DFF_302.Q ),
    .y(_00676_)
  );
  al_nand2 _05207_ (
    .a(TM1),
    .b(\DFF_302.Q ),
    .y(_00677_)
  );
  al_nand3 _05208_ (
    .a(\DFF_334.Q ),
    .b(_00676_),
    .c(_00677_),
    .y(_00678_)
  );
  al_nand2ft _05209_ (
    .a(TM1),
    .b(\DFF_302.Q ),
    .y(_00679_)
  );
  al_nand2ft _05210_ (
    .a(\DFF_302.Q ),
    .b(TM1),
    .y(_00680_)
  );
  al_nand3ftt _05211_ (
    .a(\DFF_334.Q ),
    .b(_00679_),
    .c(_00680_),
    .y(_00681_)
  );
  al_and2ft _05212_ (
    .a(\DFF_270.Q ),
    .b(\DFF_238.Q ),
    .y(_00682_)
  );
  al_nand2ft _05213_ (
    .a(\DFF_238.Q ),
    .b(\DFF_270.Q ),
    .y(_00683_)
  );
  al_nand2ft _05214_ (
    .a(_00682_),
    .b(_00683_),
    .y(_00684_)
  );
  al_ao21 _05215_ (
    .a(_00681_),
    .b(_00678_),
    .c(_00684_),
    .y(_00685_)
  );
  al_nand3 _05216_ (
    .a(_00681_),
    .b(_00678_),
    .c(_00684_),
    .y(_00686_)
  );
  al_nand3 _05217_ (
    .a(_00448_),
    .b(_00685_),
    .c(_00686_),
    .y(_00687_)
  );
  al_aoi21 _05218_ (
    .a(TM0),
    .b(\DFF_177.Q ),
    .c(TM1),
    .y(_00688_)
  );
  al_aoi21 _05219_ (
    .a(_00688_),
    .b(_00687_),
    .c(_00451_),
    .y(_00689_)
  );
  al_aoi21ftf _05220_ (
    .a(_00675_),
    .b(_00674_),
    .c(_00689_),
    .y(\DFF_46.D )
  );
  al_nand3 _05221_ (
    .a(_00448_),
    .b(_00223_),
    .c(_00220_),
    .y(_00690_)
  );
  al_ao21ttf _05222_ (
    .a(TM0),
    .b(\DFF_15.Q ),
    .c(TM1),
    .y(_00691_)
  );
  al_or2 _05223_ (
    .a(TM1),
    .b(\DFF_303.Q ),
    .y(_00692_)
  );
  al_nand2 _05224_ (
    .a(TM1),
    .b(\DFF_303.Q ),
    .y(_00693_)
  );
  al_nand3 _05225_ (
    .a(\DFF_335.Q ),
    .b(_00692_),
    .c(_00693_),
    .y(_00694_)
  );
  al_nand2ft _05226_ (
    .a(TM1),
    .b(\DFF_303.Q ),
    .y(_00695_)
  );
  al_nand2ft _05227_ (
    .a(\DFF_303.Q ),
    .b(TM1),
    .y(_00696_)
  );
  al_nand3ftt _05228_ (
    .a(\DFF_335.Q ),
    .b(_00695_),
    .c(_00696_),
    .y(_00697_)
  );
  al_and2ft _05229_ (
    .a(\DFF_271.Q ),
    .b(\DFF_239.Q ),
    .y(_00698_)
  );
  al_nand2ft _05230_ (
    .a(\DFF_239.Q ),
    .b(\DFF_271.Q ),
    .y(_00699_)
  );
  al_nand2ft _05231_ (
    .a(_00698_),
    .b(_00699_),
    .y(_00700_)
  );
  al_ao21 _05232_ (
    .a(_00697_),
    .b(_00694_),
    .c(_00700_),
    .y(_00701_)
  );
  al_nand3 _05233_ (
    .a(_00697_),
    .b(_00694_),
    .c(_00700_),
    .y(_00702_)
  );
  al_nand3 _05234_ (
    .a(_00448_),
    .b(_00701_),
    .c(_00702_),
    .y(_00703_)
  );
  al_aoi21 _05235_ (
    .a(TM0),
    .b(\DFF_176.Q ),
    .c(TM1),
    .y(_00704_)
  );
  al_aoi21 _05236_ (
    .a(_00704_),
    .b(_00703_),
    .c(_00451_),
    .y(_00705_)
  );
  al_aoi21ftf _05237_ (
    .a(_00691_),
    .b(_00690_),
    .c(_00705_),
    .y(\DFF_47.D )
  );
  al_nand3 _05238_ (
    .a(_00448_),
    .b(_00237_),
    .c(_00234_),
    .y(_00706_)
  );
  al_aoi21ttf _05239_ (
    .a(TM0),
    .b(\DFF_16.Q ),
    .c(TM1),
    .y(_00707_)
  );
  al_and2ft _05240_ (
    .a(\DFF_272.Q ),
    .b(\DFF_304.Q ),
    .y(_00708_)
  );
  al_nand2ft _05241_ (
    .a(\DFF_304.Q ),
    .b(\DFF_272.Q ),
    .y(_00709_)
  );
  al_and2ft _05242_ (
    .a(\DFF_240.Q ),
    .b(\DFF_336.Q ),
    .y(_00710_)
  );
  al_nand2ft _05243_ (
    .a(\DFF_336.Q ),
    .b(\DFF_240.Q ),
    .y(_00711_)
  );
  al_nand2ft _05244_ (
    .a(_00710_),
    .b(_00711_),
    .y(_00712_)
  );
  al_or3ftt _05245_ (
    .a(_00709_),
    .b(_00708_),
    .c(_00712_),
    .y(_00713_)
  );
  al_ao21ftf _05246_ (
    .a(_00708_),
    .b(_00709_),
    .c(_00712_),
    .y(_00714_)
  );
  al_nand3 _05247_ (
    .a(_00448_),
    .b(_00714_),
    .c(_00713_),
    .y(_00715_)
  );
  al_aoi21 _05248_ (
    .a(TM0),
    .b(\DFF_175.Q ),
    .c(TM1),
    .y(_00716_)
  );
  al_ao21 _05249_ (
    .a(_00716_),
    .b(_00715_),
    .c(_00451_),
    .y(_00717_)
  );
  al_aoi21 _05250_ (
    .a(_00707_),
    .b(_00706_),
    .c(_00717_),
    .y(\DFF_48.D )
  );
  al_nand3 _05251_ (
    .a(_00448_),
    .b(_00251_),
    .c(_00248_),
    .y(_00718_)
  );
  al_aoi21ttf _05252_ (
    .a(TM0),
    .b(\DFF_17.Q ),
    .c(TM1),
    .y(_00719_)
  );
  al_and2ft _05253_ (
    .a(\DFF_273.Q ),
    .b(\DFF_305.Q ),
    .y(_00720_)
  );
  al_nand2ft _05254_ (
    .a(\DFF_305.Q ),
    .b(\DFF_273.Q ),
    .y(_00721_)
  );
  al_and2ft _05255_ (
    .a(\DFF_241.Q ),
    .b(\DFF_337.Q ),
    .y(_00722_)
  );
  al_nand2ft _05256_ (
    .a(\DFF_337.Q ),
    .b(\DFF_241.Q ),
    .y(_00723_)
  );
  al_nand2ft _05257_ (
    .a(_00722_),
    .b(_00723_),
    .y(_00724_)
  );
  al_or3ftt _05258_ (
    .a(_00721_),
    .b(_00720_),
    .c(_00724_),
    .y(_00725_)
  );
  al_ao21ftf _05259_ (
    .a(_00720_),
    .b(_00721_),
    .c(_00724_),
    .y(_00726_)
  );
  al_nand3 _05260_ (
    .a(_00448_),
    .b(_00726_),
    .c(_00725_),
    .y(_00727_)
  );
  al_aoi21 _05261_ (
    .a(TM0),
    .b(\DFF_174.Q ),
    .c(TM1),
    .y(_00728_)
  );
  al_ao21 _05262_ (
    .a(_00728_),
    .b(_00727_),
    .c(_00451_),
    .y(_00729_)
  );
  al_aoi21 _05263_ (
    .a(_00719_),
    .b(_00718_),
    .c(_00729_),
    .y(\DFF_49.D )
  );
  al_nand3 _05264_ (
    .a(_00448_),
    .b(_00265_),
    .c(_00262_),
    .y(_00730_)
  );
  al_aoi21ttf _05265_ (
    .a(TM0),
    .b(\DFF_18.Q ),
    .c(TM1),
    .y(_00731_)
  );
  al_and2ft _05266_ (
    .a(\DFF_274.Q ),
    .b(\DFF_306.Q ),
    .y(_00732_)
  );
  al_nand2ft _05267_ (
    .a(\DFF_306.Q ),
    .b(\DFF_274.Q ),
    .y(_00733_)
  );
  al_and2ft _05268_ (
    .a(\DFF_242.Q ),
    .b(\DFF_338.Q ),
    .y(_00734_)
  );
  al_nand2ft _05269_ (
    .a(\DFF_338.Q ),
    .b(\DFF_242.Q ),
    .y(_00735_)
  );
  al_nand2ft _05270_ (
    .a(_00734_),
    .b(_00735_),
    .y(_00736_)
  );
  al_or3ftt _05271_ (
    .a(_00733_),
    .b(_00732_),
    .c(_00736_),
    .y(_00737_)
  );
  al_ao21ftf _05272_ (
    .a(_00732_),
    .b(_00733_),
    .c(_00736_),
    .y(_00738_)
  );
  al_nand3 _05273_ (
    .a(_00448_),
    .b(_00738_),
    .c(_00737_),
    .y(_00739_)
  );
  al_aoi21 _05274_ (
    .a(TM0),
    .b(\DFF_173.Q ),
    .c(TM1),
    .y(_00740_)
  );
  al_ao21 _05275_ (
    .a(_00740_),
    .b(_00739_),
    .c(_00451_),
    .y(_00741_)
  );
  al_aoi21 _05276_ (
    .a(_00731_),
    .b(_00730_),
    .c(_00741_),
    .y(\DFF_50.D )
  );
  al_nand3 _05277_ (
    .a(_00448_),
    .b(_00279_),
    .c(_00276_),
    .y(_00742_)
  );
  al_aoi21ttf _05278_ (
    .a(TM0),
    .b(\DFF_19.Q ),
    .c(TM1),
    .y(_00743_)
  );
  al_and2ft _05279_ (
    .a(\DFF_275.Q ),
    .b(\DFF_307.Q ),
    .y(_00744_)
  );
  al_nand2ft _05280_ (
    .a(\DFF_307.Q ),
    .b(\DFF_275.Q ),
    .y(_00745_)
  );
  al_and2ft _05281_ (
    .a(\DFF_243.Q ),
    .b(\DFF_339.Q ),
    .y(_00746_)
  );
  al_nand2ft _05282_ (
    .a(\DFF_339.Q ),
    .b(\DFF_243.Q ),
    .y(_00747_)
  );
  al_nand2ft _05283_ (
    .a(_00746_),
    .b(_00747_),
    .y(_00748_)
  );
  al_or3ftt _05284_ (
    .a(_00745_),
    .b(_00744_),
    .c(_00748_),
    .y(_00749_)
  );
  al_ao21ftf _05285_ (
    .a(_00744_),
    .b(_00745_),
    .c(_00748_),
    .y(_00750_)
  );
  al_nand3 _05286_ (
    .a(_00448_),
    .b(_00750_),
    .c(_00749_),
    .y(_00751_)
  );
  al_aoi21 _05287_ (
    .a(TM0),
    .b(\DFF_172.Q ),
    .c(TM1),
    .y(_00752_)
  );
  al_ao21 _05288_ (
    .a(_00752_),
    .b(_00751_),
    .c(_00451_),
    .y(_00753_)
  );
  al_aoi21 _05289_ (
    .a(_00743_),
    .b(_00742_),
    .c(_00753_),
    .y(\DFF_51.D )
  );
  al_nand3 _05290_ (
    .a(_00448_),
    .b(_00293_),
    .c(_00290_),
    .y(_00754_)
  );
  al_aoi21ttf _05291_ (
    .a(TM0),
    .b(\DFF_20.Q ),
    .c(TM1),
    .y(_00755_)
  );
  al_and2ft _05292_ (
    .a(\DFF_276.Q ),
    .b(\DFF_308.Q ),
    .y(_00756_)
  );
  al_nand2ft _05293_ (
    .a(\DFF_308.Q ),
    .b(\DFF_276.Q ),
    .y(_00757_)
  );
  al_and2ft _05294_ (
    .a(\DFF_244.Q ),
    .b(\DFF_340.Q ),
    .y(_00758_)
  );
  al_nand2ft _05295_ (
    .a(\DFF_340.Q ),
    .b(\DFF_244.Q ),
    .y(_00759_)
  );
  al_nand2ft _05296_ (
    .a(_00758_),
    .b(_00759_),
    .y(_00760_)
  );
  al_or3ftt _05297_ (
    .a(_00757_),
    .b(_00756_),
    .c(_00760_),
    .y(_00761_)
  );
  al_ao21ftf _05298_ (
    .a(_00756_),
    .b(_00757_),
    .c(_00760_),
    .y(_00762_)
  );
  al_nand3 _05299_ (
    .a(_00448_),
    .b(_00762_),
    .c(_00761_),
    .y(_00763_)
  );
  al_aoi21 _05300_ (
    .a(TM0),
    .b(\DFF_171.Q ),
    .c(TM1),
    .y(_00764_)
  );
  al_ao21 _05301_ (
    .a(_00764_),
    .b(_00763_),
    .c(_00451_),
    .y(_00765_)
  );
  al_aoi21 _05302_ (
    .a(_00755_),
    .b(_00754_),
    .c(_00765_),
    .y(\DFF_52.D )
  );
  al_nand3 _05303_ (
    .a(_00448_),
    .b(_00307_),
    .c(_00304_),
    .y(_00766_)
  );
  al_aoi21ttf _05304_ (
    .a(TM0),
    .b(\DFF_21.Q ),
    .c(TM1),
    .y(_00767_)
  );
  al_and2ft _05305_ (
    .a(\DFF_277.Q ),
    .b(\DFF_309.Q ),
    .y(_00768_)
  );
  al_nand2ft _05306_ (
    .a(\DFF_309.Q ),
    .b(\DFF_277.Q ),
    .y(_00769_)
  );
  al_and2ft _05307_ (
    .a(\DFF_245.Q ),
    .b(\DFF_341.Q ),
    .y(_00770_)
  );
  al_nand2ft _05308_ (
    .a(\DFF_341.Q ),
    .b(\DFF_245.Q ),
    .y(_00771_)
  );
  al_nand2ft _05309_ (
    .a(_00770_),
    .b(_00771_),
    .y(_00772_)
  );
  al_or3ftt _05310_ (
    .a(_00769_),
    .b(_00768_),
    .c(_00772_),
    .y(_00773_)
  );
  al_ao21ftf _05311_ (
    .a(_00768_),
    .b(_00769_),
    .c(_00772_),
    .y(_00774_)
  );
  al_nand3 _05312_ (
    .a(_00448_),
    .b(_00774_),
    .c(_00773_),
    .y(_00775_)
  );
  al_aoi21 _05313_ (
    .a(TM0),
    .b(\DFF_170.Q ),
    .c(TM1),
    .y(_00776_)
  );
  al_ao21 _05314_ (
    .a(_00776_),
    .b(_00775_),
    .c(_00451_),
    .y(_00777_)
  );
  al_aoi21 _05315_ (
    .a(_00767_),
    .b(_00766_),
    .c(_00777_),
    .y(\DFF_53.D )
  );
  al_nand3 _05316_ (
    .a(_00448_),
    .b(_00321_),
    .c(_00318_),
    .y(_00778_)
  );
  al_aoi21ttf _05317_ (
    .a(TM0),
    .b(\DFF_22.Q ),
    .c(TM1),
    .y(_00779_)
  );
  al_and2ft _05318_ (
    .a(\DFF_278.Q ),
    .b(\DFF_310.Q ),
    .y(_00780_)
  );
  al_nand2ft _05319_ (
    .a(\DFF_310.Q ),
    .b(\DFF_278.Q ),
    .y(_00781_)
  );
  al_and2ft _05320_ (
    .a(\DFF_246.Q ),
    .b(\DFF_342.Q ),
    .y(_00782_)
  );
  al_nand2ft _05321_ (
    .a(\DFF_342.Q ),
    .b(\DFF_246.Q ),
    .y(_00783_)
  );
  al_nand2ft _05322_ (
    .a(_00782_),
    .b(_00783_),
    .y(_00784_)
  );
  al_or3ftt _05323_ (
    .a(_00781_),
    .b(_00780_),
    .c(_00784_),
    .y(_00785_)
  );
  al_ao21ftf _05324_ (
    .a(_00780_),
    .b(_00781_),
    .c(_00784_),
    .y(_00786_)
  );
  al_nand3 _05325_ (
    .a(_00448_),
    .b(_00786_),
    .c(_00785_),
    .y(_00787_)
  );
  al_aoi21 _05326_ (
    .a(TM0),
    .b(\DFF_169.Q ),
    .c(TM1),
    .y(_00788_)
  );
  al_ao21 _05327_ (
    .a(_00788_),
    .b(_00787_),
    .c(_00451_),
    .y(_00789_)
  );
  al_aoi21 _05328_ (
    .a(_00779_),
    .b(_00778_),
    .c(_00789_),
    .y(\DFF_54.D )
  );
  al_nand3 _05329_ (
    .a(_00448_),
    .b(_00335_),
    .c(_00332_),
    .y(_00790_)
  );
  al_aoi21ttf _05330_ (
    .a(TM0),
    .b(\DFF_23.Q ),
    .c(TM1),
    .y(_00791_)
  );
  al_and2ft _05331_ (
    .a(\DFF_279.Q ),
    .b(\DFF_311.Q ),
    .y(_00792_)
  );
  al_nand2ft _05332_ (
    .a(\DFF_311.Q ),
    .b(\DFF_279.Q ),
    .y(_00793_)
  );
  al_and2ft _05333_ (
    .a(\DFF_247.Q ),
    .b(\DFF_343.Q ),
    .y(_00794_)
  );
  al_nand2ft _05334_ (
    .a(\DFF_343.Q ),
    .b(\DFF_247.Q ),
    .y(_00795_)
  );
  al_nand2ft _05335_ (
    .a(_00794_),
    .b(_00795_),
    .y(_00796_)
  );
  al_or3ftt _05336_ (
    .a(_00793_),
    .b(_00792_),
    .c(_00796_),
    .y(_00797_)
  );
  al_ao21ftf _05337_ (
    .a(_00792_),
    .b(_00793_),
    .c(_00796_),
    .y(_00798_)
  );
  al_nand3 _05338_ (
    .a(_00448_),
    .b(_00798_),
    .c(_00797_),
    .y(_00799_)
  );
  al_aoi21 _05339_ (
    .a(TM0),
    .b(\DFF_168.Q ),
    .c(TM1),
    .y(_00800_)
  );
  al_ao21 _05340_ (
    .a(_00800_),
    .b(_00799_),
    .c(_00451_),
    .y(_00801_)
  );
  al_aoi21 _05341_ (
    .a(_00791_),
    .b(_00790_),
    .c(_00801_),
    .y(\DFF_55.D )
  );
  al_nand3 _05342_ (
    .a(_00448_),
    .b(_00349_),
    .c(_00346_),
    .y(_00802_)
  );
  al_aoi21ttf _05343_ (
    .a(TM0),
    .b(\DFF_24.Q ),
    .c(TM1),
    .y(_00803_)
  );
  al_and2ft _05344_ (
    .a(\DFF_280.Q ),
    .b(\DFF_312.Q ),
    .y(_00804_)
  );
  al_nand2ft _05345_ (
    .a(\DFF_312.Q ),
    .b(\DFF_280.Q ),
    .y(_00805_)
  );
  al_and2ft _05346_ (
    .a(\DFF_248.Q ),
    .b(\DFF_344.Q ),
    .y(_00806_)
  );
  al_nand2ft _05347_ (
    .a(\DFF_344.Q ),
    .b(\DFF_248.Q ),
    .y(_00807_)
  );
  al_nand2ft _05348_ (
    .a(_00806_),
    .b(_00807_),
    .y(_00808_)
  );
  al_or3ftt _05349_ (
    .a(_00805_),
    .b(_00804_),
    .c(_00808_),
    .y(_00809_)
  );
  al_ao21ftf _05350_ (
    .a(_00804_),
    .b(_00805_),
    .c(_00808_),
    .y(_00810_)
  );
  al_nand3 _05351_ (
    .a(_00448_),
    .b(_00810_),
    .c(_00809_),
    .y(_00811_)
  );
  al_aoi21 _05352_ (
    .a(TM0),
    .b(\DFF_167.Q ),
    .c(TM1),
    .y(_00812_)
  );
  al_ao21 _05353_ (
    .a(_00812_),
    .b(_00811_),
    .c(_00451_),
    .y(_00813_)
  );
  al_aoi21 _05354_ (
    .a(_00803_),
    .b(_00802_),
    .c(_00813_),
    .y(\DFF_56.D )
  );
  al_nand3 _05355_ (
    .a(_00448_),
    .b(_00363_),
    .c(_00360_),
    .y(_00814_)
  );
  al_aoi21ttf _05356_ (
    .a(TM0),
    .b(\DFF_25.Q ),
    .c(TM1),
    .y(_00815_)
  );
  al_and2ft _05357_ (
    .a(\DFF_281.Q ),
    .b(\DFF_313.Q ),
    .y(_00816_)
  );
  al_nand2ft _05358_ (
    .a(\DFF_313.Q ),
    .b(\DFF_281.Q ),
    .y(_00817_)
  );
  al_and2ft _05359_ (
    .a(\DFF_249.Q ),
    .b(\DFF_345.Q ),
    .y(_00818_)
  );
  al_nand2ft _05360_ (
    .a(\DFF_345.Q ),
    .b(\DFF_249.Q ),
    .y(_00819_)
  );
  al_nand2ft _05361_ (
    .a(_00818_),
    .b(_00819_),
    .y(_00820_)
  );
  al_or3ftt _05362_ (
    .a(_00817_),
    .b(_00816_),
    .c(_00820_),
    .y(_00821_)
  );
  al_ao21ftf _05363_ (
    .a(_00816_),
    .b(_00817_),
    .c(_00820_),
    .y(_00822_)
  );
  al_nand3 _05364_ (
    .a(_00448_),
    .b(_00822_),
    .c(_00821_),
    .y(_00823_)
  );
  al_aoi21 _05365_ (
    .a(TM0),
    .b(\DFF_166.Q ),
    .c(TM1),
    .y(_00824_)
  );
  al_ao21 _05366_ (
    .a(_00824_),
    .b(_00823_),
    .c(_00451_),
    .y(_00825_)
  );
  al_aoi21 _05367_ (
    .a(_00815_),
    .b(_00814_),
    .c(_00825_),
    .y(\DFF_57.D )
  );
  al_nand3 _05368_ (
    .a(_00448_),
    .b(_00377_),
    .c(_00374_),
    .y(_00826_)
  );
  al_aoi21ttf _05369_ (
    .a(TM0),
    .b(\DFF_26.Q ),
    .c(TM1),
    .y(_00827_)
  );
  al_and2ft _05370_ (
    .a(\DFF_282.Q ),
    .b(\DFF_314.Q ),
    .y(_00828_)
  );
  al_nand2ft _05371_ (
    .a(\DFF_314.Q ),
    .b(\DFF_282.Q ),
    .y(_00829_)
  );
  al_and2ft _05372_ (
    .a(\DFF_250.Q ),
    .b(\DFF_346.Q ),
    .y(_00830_)
  );
  al_nand2ft _05373_ (
    .a(\DFF_346.Q ),
    .b(\DFF_250.Q ),
    .y(_00831_)
  );
  al_nand2ft _05374_ (
    .a(_00830_),
    .b(_00831_),
    .y(_00832_)
  );
  al_or3ftt _05375_ (
    .a(_00829_),
    .b(_00828_),
    .c(_00832_),
    .y(_00833_)
  );
  al_ao21ftf _05376_ (
    .a(_00828_),
    .b(_00829_),
    .c(_00832_),
    .y(_00834_)
  );
  al_nand3 _05377_ (
    .a(_00448_),
    .b(_00834_),
    .c(_00833_),
    .y(_00835_)
  );
  al_aoi21 _05378_ (
    .a(TM0),
    .b(\DFF_165.Q ),
    .c(TM1),
    .y(_00836_)
  );
  al_ao21 _05379_ (
    .a(_00836_),
    .b(_00835_),
    .c(_00451_),
    .y(_00837_)
  );
  al_aoi21 _05380_ (
    .a(_00827_),
    .b(_00826_),
    .c(_00837_),
    .y(\DFF_58.D )
  );
  al_nand3 _05381_ (
    .a(_00448_),
    .b(_00391_),
    .c(_00388_),
    .y(_00838_)
  );
  al_aoi21ttf _05382_ (
    .a(TM0),
    .b(\DFF_27.Q ),
    .c(TM1),
    .y(_00839_)
  );
  al_and2ft _05383_ (
    .a(\DFF_283.Q ),
    .b(\DFF_315.Q ),
    .y(_00840_)
  );
  al_nand2ft _05384_ (
    .a(\DFF_315.Q ),
    .b(\DFF_283.Q ),
    .y(_00841_)
  );
  al_and2ft _05385_ (
    .a(\DFF_251.Q ),
    .b(\DFF_347.Q ),
    .y(_00842_)
  );
  al_nand2ft _05386_ (
    .a(\DFF_347.Q ),
    .b(\DFF_251.Q ),
    .y(_00843_)
  );
  al_nand2ft _05387_ (
    .a(_00842_),
    .b(_00843_),
    .y(_00844_)
  );
  al_or3ftt _05388_ (
    .a(_00841_),
    .b(_00840_),
    .c(_00844_),
    .y(_00845_)
  );
  al_ao21ftf _05389_ (
    .a(_00840_),
    .b(_00841_),
    .c(_00844_),
    .y(_00846_)
  );
  al_nand3 _05390_ (
    .a(_00448_),
    .b(_00846_),
    .c(_00845_),
    .y(_00847_)
  );
  al_aoi21 _05391_ (
    .a(TM0),
    .b(\DFF_164.Q ),
    .c(TM1),
    .y(_00848_)
  );
  al_ao21 _05392_ (
    .a(_00848_),
    .b(_00847_),
    .c(_00451_),
    .y(_00849_)
  );
  al_aoi21 _05393_ (
    .a(_00839_),
    .b(_00838_),
    .c(_00849_),
    .y(\DFF_59.D )
  );
  al_nand3 _05394_ (
    .a(_00448_),
    .b(_00405_),
    .c(_00402_),
    .y(_00850_)
  );
  al_aoi21ttf _05395_ (
    .a(TM0),
    .b(\DFF_28.Q ),
    .c(TM1),
    .y(_00851_)
  );
  al_and2ft _05396_ (
    .a(\DFF_284.Q ),
    .b(\DFF_316.Q ),
    .y(_00852_)
  );
  al_nand2ft _05397_ (
    .a(\DFF_316.Q ),
    .b(\DFF_284.Q ),
    .y(_00853_)
  );
  al_and2ft _05398_ (
    .a(\DFF_252.Q ),
    .b(\DFF_348.Q ),
    .y(_00854_)
  );
  al_nand2ft _05399_ (
    .a(\DFF_348.Q ),
    .b(\DFF_252.Q ),
    .y(_00855_)
  );
  al_nand2ft _05400_ (
    .a(_00854_),
    .b(_00855_),
    .y(_00856_)
  );
  al_or3ftt _05401_ (
    .a(_00853_),
    .b(_00852_),
    .c(_00856_),
    .y(_00857_)
  );
  al_ao21ftf _05402_ (
    .a(_00852_),
    .b(_00853_),
    .c(_00856_),
    .y(_00858_)
  );
  al_nand3 _05403_ (
    .a(_00448_),
    .b(_00858_),
    .c(_00857_),
    .y(_00859_)
  );
  al_aoi21 _05404_ (
    .a(TM0),
    .b(\DFF_163.Q ),
    .c(TM1),
    .y(_00860_)
  );
  al_ao21 _05405_ (
    .a(_00860_),
    .b(_00859_),
    .c(_00451_),
    .y(_00861_)
  );
  al_aoi21 _05406_ (
    .a(_00851_),
    .b(_00850_),
    .c(_00861_),
    .y(\DFF_60.D )
  );
  al_nand3 _05407_ (
    .a(_00448_),
    .b(_00419_),
    .c(_00416_),
    .y(_00862_)
  );
  al_aoi21ttf _05408_ (
    .a(TM0),
    .b(\DFF_29.Q ),
    .c(TM1),
    .y(_00863_)
  );
  al_and2ft _05409_ (
    .a(\DFF_285.Q ),
    .b(\DFF_317.Q ),
    .y(_00864_)
  );
  al_nand2ft _05410_ (
    .a(\DFF_317.Q ),
    .b(\DFF_285.Q ),
    .y(_00865_)
  );
  al_and2ft _05411_ (
    .a(\DFF_253.Q ),
    .b(\DFF_349.Q ),
    .y(_00866_)
  );
  al_nand2ft _05412_ (
    .a(\DFF_349.Q ),
    .b(\DFF_253.Q ),
    .y(_00867_)
  );
  al_nand2ft _05413_ (
    .a(_00866_),
    .b(_00867_),
    .y(_00868_)
  );
  al_or3ftt _05414_ (
    .a(_00865_),
    .b(_00864_),
    .c(_00868_),
    .y(_00869_)
  );
  al_ao21ftf _05415_ (
    .a(_00864_),
    .b(_00865_),
    .c(_00868_),
    .y(_00870_)
  );
  al_nand3 _05416_ (
    .a(_00448_),
    .b(_00870_),
    .c(_00869_),
    .y(_00871_)
  );
  al_aoi21 _05417_ (
    .a(TM0),
    .b(\DFF_162.Q ),
    .c(TM1),
    .y(_00872_)
  );
  al_ao21 _05418_ (
    .a(_00872_),
    .b(_00871_),
    .c(_00451_),
    .y(_00873_)
  );
  al_aoi21 _05419_ (
    .a(_00863_),
    .b(_00862_),
    .c(_00873_),
    .y(\DFF_61.D )
  );
  al_nand3 _05420_ (
    .a(_00448_),
    .b(_00433_),
    .c(_00430_),
    .y(_00874_)
  );
  al_aoi21ttf _05421_ (
    .a(TM0),
    .b(\DFF_30.Q ),
    .c(TM1),
    .y(_00875_)
  );
  al_and2ft _05422_ (
    .a(\DFF_286.Q ),
    .b(\DFF_318.Q ),
    .y(_00876_)
  );
  al_nand2ft _05423_ (
    .a(\DFF_318.Q ),
    .b(\DFF_286.Q ),
    .y(_00877_)
  );
  al_and2ft _05424_ (
    .a(\DFF_254.Q ),
    .b(\DFF_350.Q ),
    .y(_00878_)
  );
  al_nand2ft _05425_ (
    .a(\DFF_350.Q ),
    .b(\DFF_254.Q ),
    .y(_00879_)
  );
  al_nand2ft _05426_ (
    .a(_00878_),
    .b(_00879_),
    .y(_00880_)
  );
  al_or3ftt _05427_ (
    .a(_00877_),
    .b(_00876_),
    .c(_00880_),
    .y(_00881_)
  );
  al_ao21ftf _05428_ (
    .a(_00876_),
    .b(_00877_),
    .c(_00880_),
    .y(_00882_)
  );
  al_nand3 _05429_ (
    .a(_00448_),
    .b(_00882_),
    .c(_00881_),
    .y(_00883_)
  );
  al_aoi21 _05430_ (
    .a(TM0),
    .b(\DFF_161.Q ),
    .c(TM1),
    .y(_00884_)
  );
  al_ao21 _05431_ (
    .a(_00884_),
    .b(_00883_),
    .c(_00451_),
    .y(_00885_)
  );
  al_aoi21 _05432_ (
    .a(_00875_),
    .b(_00874_),
    .c(_00885_),
    .y(\DFF_62.D )
  );
  al_nand3 _05433_ (
    .a(_00448_),
    .b(_00447_),
    .c(_00444_),
    .y(_00886_)
  );
  al_aoi21ttf _05434_ (
    .a(TM0),
    .b(\DFF_31.Q ),
    .c(TM1),
    .y(_00887_)
  );
  al_and2ft _05435_ (
    .a(\DFF_287.Q ),
    .b(\DFF_319.Q ),
    .y(_00888_)
  );
  al_nand2ft _05436_ (
    .a(\DFF_319.Q ),
    .b(\DFF_287.Q ),
    .y(_00889_)
  );
  al_and2ft _05437_ (
    .a(\DFF_255.Q ),
    .b(\DFF_351.Q ),
    .y(_00890_)
  );
  al_nand2ft _05438_ (
    .a(\DFF_351.Q ),
    .b(\DFF_255.Q ),
    .y(_00891_)
  );
  al_nand2ft _05439_ (
    .a(_00890_),
    .b(_00891_),
    .y(_00892_)
  );
  al_or3ftt _05440_ (
    .a(_00889_),
    .b(_00888_),
    .c(_00892_),
    .y(_00893_)
  );
  al_ao21ftf _05441_ (
    .a(_00888_),
    .b(_00889_),
    .c(_00892_),
    .y(_00894_)
  );
  al_nand3 _05442_ (
    .a(_00448_),
    .b(_00894_),
    .c(_00893_),
    .y(_00895_)
  );
  al_aoi21 _05443_ (
    .a(TM0),
    .b(\DFF_160.Q ),
    .c(TM1),
    .y(_00896_)
  );
  al_ao21 _05444_ (
    .a(_00896_),
    .b(_00895_),
    .c(_00451_),
    .y(_00897_)
  );
  al_aoi21 _05445_ (
    .a(_00887_),
    .b(_00886_),
    .c(_00897_),
    .y(\DFF_63.D )
  );
  al_and2 _05446_ (
    .a(RESET),
    .b(\DFF_32.Q ),
    .y(\DFF_64.D )
  );
  al_and2 _05447_ (
    .a(RESET),
    .b(\DFF_33.Q ),
    .y(\DFF_65.D )
  );
  al_and2 _05448_ (
    .a(RESET),
    .b(\DFF_34.Q ),
    .y(\DFF_66.D )
  );
  al_and2 _05449_ (
    .a(RESET),
    .b(\DFF_35.Q ),
    .y(\DFF_67.D )
  );
  al_and2 _05450_ (
    .a(RESET),
    .b(\DFF_36.Q ),
    .y(\DFF_68.D )
  );
  al_and2 _05451_ (
    .a(RESET),
    .b(\DFF_37.Q ),
    .y(\DFF_69.D )
  );
  al_and2 _05452_ (
    .a(RESET),
    .b(\DFF_38.Q ),
    .y(\DFF_70.D )
  );
  al_and2 _05453_ (
    .a(RESET),
    .b(\DFF_39.Q ),
    .y(\DFF_71.D )
  );
  al_and2 _05454_ (
    .a(RESET),
    .b(\DFF_40.Q ),
    .y(\DFF_72.D )
  );
  al_and2 _05455_ (
    .a(RESET),
    .b(\DFF_41.Q ),
    .y(\DFF_73.D )
  );
  al_and2 _05456_ (
    .a(RESET),
    .b(\DFF_42.Q ),
    .y(\DFF_74.D )
  );
  al_and2 _05457_ (
    .a(RESET),
    .b(\DFF_43.Q ),
    .y(\DFF_75.D )
  );
  al_and2 _05458_ (
    .a(RESET),
    .b(\DFF_44.Q ),
    .y(\DFF_76.D )
  );
  al_and2 _05459_ (
    .a(RESET),
    .b(\DFF_45.Q ),
    .y(\DFF_77.D )
  );
  al_and2 _05460_ (
    .a(RESET),
    .b(\DFF_46.Q ),
    .y(\DFF_78.D )
  );
  al_and2 _05461_ (
    .a(RESET),
    .b(\DFF_47.Q ),
    .y(\DFF_79.D )
  );
  al_and2 _05462_ (
    .a(RESET),
    .b(\DFF_48.Q ),
    .y(\DFF_80.D )
  );
  al_and2 _05463_ (
    .a(RESET),
    .b(\DFF_49.Q ),
    .y(\DFF_81.D )
  );
  al_and2 _05464_ (
    .a(RESET),
    .b(\DFF_50.Q ),
    .y(\DFF_82.D )
  );
  al_and2 _05465_ (
    .a(RESET),
    .b(\DFF_51.Q ),
    .y(\DFF_83.D )
  );
  al_and2 _05466_ (
    .a(RESET),
    .b(\DFF_52.Q ),
    .y(\DFF_84.D )
  );
  al_and2 _05467_ (
    .a(RESET),
    .b(\DFF_53.Q ),
    .y(\DFF_85.D )
  );
  al_and2 _05468_ (
    .a(RESET),
    .b(\DFF_54.Q ),
    .y(\DFF_86.D )
  );
  al_and2 _05469_ (
    .a(RESET),
    .b(\DFF_55.Q ),
    .y(\DFF_87.D )
  );
  al_and2 _05470_ (
    .a(RESET),
    .b(\DFF_56.Q ),
    .y(\DFF_88.D )
  );
  al_and2 _05471_ (
    .a(RESET),
    .b(\DFF_57.Q ),
    .y(\DFF_89.D )
  );
  al_and2 _05472_ (
    .a(RESET),
    .b(\DFF_58.Q ),
    .y(\DFF_90.D )
  );
  al_and2 _05473_ (
    .a(RESET),
    .b(\DFF_59.Q ),
    .y(\DFF_91.D )
  );
  al_and2 _05474_ (
    .a(RESET),
    .b(\DFF_60.Q ),
    .y(\DFF_92.D )
  );
  al_and2 _05475_ (
    .a(RESET),
    .b(\DFF_61.Q ),
    .y(\DFF_93.D )
  );
  al_and2 _05476_ (
    .a(RESET),
    .b(\DFF_62.Q ),
    .y(\DFF_94.D )
  );
  al_and2 _05477_ (
    .a(RESET),
    .b(\DFF_63.Q ),
    .y(\DFF_95.D )
  );
  al_and2 _05478_ (
    .a(RESET),
    .b(\DFF_64.Q ),
    .y(\DFF_96.D )
  );
  al_and2 _05479_ (
    .a(RESET),
    .b(\DFF_65.Q ),
    .y(\DFF_97.D )
  );
  al_and2 _05480_ (
    .a(RESET),
    .b(\DFF_66.Q ),
    .y(\DFF_98.D )
  );
  al_and2 _05481_ (
    .a(RESET),
    .b(\DFF_67.Q ),
    .y(\DFF_99.D )
  );
  al_and2 _05482_ (
    .a(RESET),
    .b(\DFF_68.Q ),
    .y(\DFF_100.D )
  );
  al_and2 _05483_ (
    .a(RESET),
    .b(\DFF_69.Q ),
    .y(\DFF_101.D )
  );
  al_and2 _05484_ (
    .a(RESET),
    .b(\DFF_70.Q ),
    .y(\DFF_102.D )
  );
  al_and2 _05485_ (
    .a(RESET),
    .b(\DFF_71.Q ),
    .y(\DFF_103.D )
  );
  al_and2 _05486_ (
    .a(RESET),
    .b(\DFF_72.Q ),
    .y(\DFF_104.D )
  );
  al_and2 _05487_ (
    .a(RESET),
    .b(\DFF_73.Q ),
    .y(\DFF_105.D )
  );
  al_and2 _05488_ (
    .a(RESET),
    .b(\DFF_74.Q ),
    .y(\DFF_106.D )
  );
  al_and2 _05489_ (
    .a(RESET),
    .b(\DFF_75.Q ),
    .y(\DFF_107.D )
  );
  al_and2 _05490_ (
    .a(RESET),
    .b(\DFF_76.Q ),
    .y(\DFF_108.D )
  );
  al_and2 _05491_ (
    .a(RESET),
    .b(\DFF_77.Q ),
    .y(\DFF_109.D )
  );
  al_and2 _05492_ (
    .a(RESET),
    .b(\DFF_78.Q ),
    .y(\DFF_110.D )
  );
  al_and2 _05493_ (
    .a(RESET),
    .b(\DFF_79.Q ),
    .y(\DFF_111.D )
  );
  al_and2 _05494_ (
    .a(RESET),
    .b(\DFF_80.Q ),
    .y(\DFF_112.D )
  );
  al_and2 _05495_ (
    .a(RESET),
    .b(\DFF_81.Q ),
    .y(\DFF_113.D )
  );
  al_and2 _05496_ (
    .a(RESET),
    .b(\DFF_82.Q ),
    .y(\DFF_114.D )
  );
  al_and2 _05497_ (
    .a(RESET),
    .b(\DFF_83.Q ),
    .y(\DFF_115.D )
  );
  al_and2 _05498_ (
    .a(RESET),
    .b(\DFF_84.Q ),
    .y(\DFF_116.D )
  );
  al_and2 _05499_ (
    .a(RESET),
    .b(\DFF_85.Q ),
    .y(\DFF_117.D )
  );
  al_and2 _05500_ (
    .a(RESET),
    .b(\DFF_86.Q ),
    .y(\DFF_118.D )
  );
  al_and2 _05501_ (
    .a(RESET),
    .b(\DFF_87.Q ),
    .y(\DFF_119.D )
  );
  al_and2 _05502_ (
    .a(RESET),
    .b(\DFF_88.Q ),
    .y(\DFF_120.D )
  );
  al_and2 _05503_ (
    .a(RESET),
    .b(\DFF_89.Q ),
    .y(\DFF_121.D )
  );
  al_and2 _05504_ (
    .a(RESET),
    .b(\DFF_90.Q ),
    .y(\DFF_122.D )
  );
  al_and2 _05505_ (
    .a(RESET),
    .b(\DFF_91.Q ),
    .y(\DFF_123.D )
  );
  al_and2 _05506_ (
    .a(RESET),
    .b(\DFF_92.Q ),
    .y(\DFF_124.D )
  );
  al_and2 _05507_ (
    .a(RESET),
    .b(\DFF_93.Q ),
    .y(\DFF_125.D )
  );
  al_and2 _05508_ (
    .a(RESET),
    .b(\DFF_94.Q ),
    .y(\DFF_126.D )
  );
  al_and2 _05509_ (
    .a(RESET),
    .b(\DFF_95.Q ),
    .y(\DFF_127.D )
  );
  al_and2 _05510_ (
    .a(RESET),
    .b(\DFF_96.Q ),
    .y(\DFF_128.D )
  );
  al_and2 _05511_ (
    .a(RESET),
    .b(\DFF_97.Q ),
    .y(\DFF_129.D )
  );
  al_and2 _05512_ (
    .a(RESET),
    .b(\DFF_98.Q ),
    .y(\DFF_130.D )
  );
  al_and2 _05513_ (
    .a(RESET),
    .b(\DFF_99.Q ),
    .y(\DFF_131.D )
  );
  al_and2 _05514_ (
    .a(RESET),
    .b(\DFF_100.Q ),
    .y(\DFF_132.D )
  );
  al_and2 _05515_ (
    .a(RESET),
    .b(\DFF_101.Q ),
    .y(\DFF_133.D )
  );
  al_and2 _05516_ (
    .a(RESET),
    .b(\DFF_102.Q ),
    .y(\DFF_134.D )
  );
  al_and2 _05517_ (
    .a(RESET),
    .b(\DFF_103.Q ),
    .y(\DFF_135.D )
  );
  al_and2 _05518_ (
    .a(RESET),
    .b(\DFF_104.Q ),
    .y(\DFF_136.D )
  );
  al_and2 _05519_ (
    .a(RESET),
    .b(\DFF_105.Q ),
    .y(\DFF_137.D )
  );
  al_and2 _05520_ (
    .a(RESET),
    .b(\DFF_106.Q ),
    .y(\DFF_138.D )
  );
  al_and2 _05521_ (
    .a(RESET),
    .b(\DFF_107.Q ),
    .y(\DFF_139.D )
  );
  al_and2 _05522_ (
    .a(RESET),
    .b(\DFF_108.Q ),
    .y(\DFF_140.D )
  );
  al_and2 _05523_ (
    .a(RESET),
    .b(\DFF_109.Q ),
    .y(\DFF_141.D )
  );
  al_and2 _05524_ (
    .a(RESET),
    .b(\DFF_110.Q ),
    .y(\DFF_142.D )
  );
  al_and2 _05525_ (
    .a(RESET),
    .b(\DFF_111.Q ),
    .y(\DFF_143.D )
  );
  al_and2 _05526_ (
    .a(RESET),
    .b(\DFF_112.Q ),
    .y(\DFF_144.D )
  );
  al_and2 _05527_ (
    .a(RESET),
    .b(\DFF_113.Q ),
    .y(\DFF_145.D )
  );
  al_and2 _05528_ (
    .a(RESET),
    .b(\DFF_114.Q ),
    .y(\DFF_146.D )
  );
  al_and2 _05529_ (
    .a(RESET),
    .b(\DFF_115.Q ),
    .y(\DFF_147.D )
  );
  al_and2 _05530_ (
    .a(RESET),
    .b(\DFF_116.Q ),
    .y(\DFF_148.D )
  );
  al_and2 _05531_ (
    .a(RESET),
    .b(\DFF_117.Q ),
    .y(\DFF_149.D )
  );
  al_and2 _05532_ (
    .a(RESET),
    .b(\DFF_118.Q ),
    .y(\DFF_150.D )
  );
  al_and2 _05533_ (
    .a(RESET),
    .b(\DFF_119.Q ),
    .y(\DFF_151.D )
  );
  al_and2 _05534_ (
    .a(RESET),
    .b(\DFF_120.Q ),
    .y(\DFF_152.D )
  );
  al_and2 _05535_ (
    .a(RESET),
    .b(\DFF_121.Q ),
    .y(\DFF_153.D )
  );
  al_and2 _05536_ (
    .a(RESET),
    .b(\DFF_122.Q ),
    .y(\DFF_154.D )
  );
  al_and2 _05537_ (
    .a(RESET),
    .b(\DFF_123.Q ),
    .y(\DFF_155.D )
  );
  al_and2 _05538_ (
    .a(RESET),
    .b(\DFF_124.Q ),
    .y(\DFF_156.D )
  );
  al_and2 _05539_ (
    .a(RESET),
    .b(\DFF_125.Q ),
    .y(\DFF_157.D )
  );
  al_and2 _05540_ (
    .a(RESET),
    .b(\DFF_126.Q ),
    .y(\DFF_158.D )
  );
  al_and2 _05541_ (
    .a(RESET),
    .b(\DFF_127.Q ),
    .y(\DFF_159.D )
  );
  al_oa21ftt _05542_ (
    .a(\DFF_159.Q ),
    .b(\DFF_191.Q ),
    .c(RESET),
    .y(_00898_)
  );
  al_aoi21ftf _05543_ (
    .a(\DFF_159.Q ),
    .b(\DFF_191.Q ),
    .c(_00898_),
    .y(\DFF_160.D )
  );
  al_oa21ftt _05544_ (
    .a(\DFF_158.Q ),
    .b(\DFF_160.Q ),
    .c(RESET),
    .y(_00899_)
  );
  al_aoi21ftf _05545_ (
    .a(\DFF_158.Q ),
    .b(\DFF_160.Q ),
    .c(_00899_),
    .y(\DFF_161.D )
  );
  al_oa21ftt _05546_ (
    .a(\DFF_157.Q ),
    .b(\DFF_161.Q ),
    .c(RESET),
    .y(_00900_)
  );
  al_aoi21ftf _05547_ (
    .a(\DFF_157.Q ),
    .b(\DFF_161.Q ),
    .c(_00900_),
    .y(\DFF_162.D )
  );
  al_oa21ftt _05548_ (
    .a(\DFF_156.Q ),
    .b(\DFF_162.Q ),
    .c(RESET),
    .y(_00901_)
  );
  al_aoi21ftf _05549_ (
    .a(\DFF_156.Q ),
    .b(\DFF_162.Q ),
    .c(_00901_),
    .y(\DFF_163.D )
  );
  al_nand2ft _05550_ (
    .a(\DFF_155.Q ),
    .b(\DFF_191.Q ),
    .y(_00902_)
  );
  al_nand2ft _05551_ (
    .a(\DFF_191.Q ),
    .b(\DFF_155.Q ),
    .y(_00903_)
  );
  al_ao21ttf _05552_ (
    .a(_00902_),
    .b(_00903_),
    .c(\DFF_163.Q ),
    .y(_00904_)
  );
  al_nand3ftt _05553_ (
    .a(\DFF_163.Q ),
    .b(_00902_),
    .c(_00903_),
    .y(_00905_)
  );
  al_aoi21 _05554_ (
    .a(_00905_),
    .b(_00904_),
    .c(_00451_),
    .y(\DFF_164.D )
  );
  al_oa21ftt _05555_ (
    .a(\DFF_154.Q ),
    .b(\DFF_164.Q ),
    .c(RESET),
    .y(_00906_)
  );
  al_aoi21ftf _05556_ (
    .a(\DFF_154.Q ),
    .b(\DFF_164.Q ),
    .c(_00906_),
    .y(\DFF_165.D )
  );
  al_oa21ftt _05557_ (
    .a(\DFF_153.Q ),
    .b(\DFF_165.Q ),
    .c(RESET),
    .y(_00907_)
  );
  al_aoi21ftf _05558_ (
    .a(\DFF_153.Q ),
    .b(\DFF_165.Q ),
    .c(_00907_),
    .y(\DFF_166.D )
  );
  al_oa21ftt _05559_ (
    .a(\DFF_152.Q ),
    .b(\DFF_166.Q ),
    .c(RESET),
    .y(_00908_)
  );
  al_aoi21ftf _05560_ (
    .a(\DFF_152.Q ),
    .b(\DFF_166.Q ),
    .c(_00908_),
    .y(\DFF_167.D )
  );
  al_oa21ftt _05561_ (
    .a(\DFF_151.Q ),
    .b(\DFF_167.Q ),
    .c(RESET),
    .y(_00909_)
  );
  al_aoi21ftf _05562_ (
    .a(\DFF_151.Q ),
    .b(\DFF_167.Q ),
    .c(_00909_),
    .y(\DFF_168.D )
  );
  al_oa21ftt _05563_ (
    .a(\DFF_150.Q ),
    .b(\DFF_168.Q ),
    .c(RESET),
    .y(_00910_)
  );
  al_aoi21ftf _05564_ (
    .a(\DFF_150.Q ),
    .b(\DFF_168.Q ),
    .c(_00910_),
    .y(\DFF_169.D )
  );
  al_oa21ftt _05565_ (
    .a(\DFF_149.Q ),
    .b(\DFF_169.Q ),
    .c(RESET),
    .y(_00911_)
  );
  al_aoi21ftf _05566_ (
    .a(\DFF_149.Q ),
    .b(\DFF_169.Q ),
    .c(_00911_),
    .y(\DFF_170.D )
  );
  al_nand2ft _05567_ (
    .a(\DFF_148.Q ),
    .b(\DFF_191.Q ),
    .y(_00912_)
  );
  al_nand2ft _05568_ (
    .a(\DFF_191.Q ),
    .b(\DFF_148.Q ),
    .y(_00913_)
  );
  al_ao21ttf _05569_ (
    .a(_00912_),
    .b(_00913_),
    .c(\DFF_170.Q ),
    .y(_00914_)
  );
  al_nand3ftt _05570_ (
    .a(\DFF_170.Q ),
    .b(_00912_),
    .c(_00913_),
    .y(_00915_)
  );
  al_aoi21 _05571_ (
    .a(_00915_),
    .b(_00914_),
    .c(_00451_),
    .y(\DFF_171.D )
  );
  al_oa21ftt _05572_ (
    .a(\DFF_147.Q ),
    .b(\DFF_171.Q ),
    .c(RESET),
    .y(_00916_)
  );
  al_aoi21ftf _05573_ (
    .a(\DFF_147.Q ),
    .b(\DFF_171.Q ),
    .c(_00916_),
    .y(\DFF_172.D )
  );
  al_oa21ftt _05574_ (
    .a(\DFF_146.Q ),
    .b(\DFF_172.Q ),
    .c(RESET),
    .y(_00917_)
  );
  al_aoi21ftf _05575_ (
    .a(\DFF_146.Q ),
    .b(\DFF_172.Q ),
    .c(_00917_),
    .y(\DFF_173.D )
  );
  al_oa21ftt _05576_ (
    .a(\DFF_145.Q ),
    .b(\DFF_173.Q ),
    .c(RESET),
    .y(_00918_)
  );
  al_aoi21ftf _05577_ (
    .a(\DFF_145.Q ),
    .b(\DFF_173.Q ),
    .c(_00918_),
    .y(\DFF_174.D )
  );
  al_oa21ftt _05578_ (
    .a(\DFF_144.Q ),
    .b(\DFF_174.Q ),
    .c(RESET),
    .y(_00919_)
  );
  al_aoi21ftf _05579_ (
    .a(\DFF_144.Q ),
    .b(\DFF_174.Q ),
    .c(_00919_),
    .y(\DFF_175.D )
  );
  al_nand2ft _05580_ (
    .a(\DFF_143.Q ),
    .b(\DFF_191.Q ),
    .y(_00920_)
  );
  al_nand2ft _05581_ (
    .a(\DFF_191.Q ),
    .b(\DFF_143.Q ),
    .y(_00921_)
  );
  al_ao21ttf _05582_ (
    .a(_00920_),
    .b(_00921_),
    .c(\DFF_175.Q ),
    .y(_00922_)
  );
  al_nand3ftt _05583_ (
    .a(\DFF_175.Q ),
    .b(_00920_),
    .c(_00921_),
    .y(_00923_)
  );
  al_aoi21 _05584_ (
    .a(_00923_),
    .b(_00922_),
    .c(_00451_),
    .y(\DFF_176.D )
  );
  al_oa21ftt _05585_ (
    .a(\DFF_142.Q ),
    .b(\DFF_176.Q ),
    .c(RESET),
    .y(_00924_)
  );
  al_aoi21ftf _05586_ (
    .a(\DFF_142.Q ),
    .b(\DFF_176.Q ),
    .c(_00924_),
    .y(\DFF_177.D )
  );
  al_oa21ftt _05587_ (
    .a(\DFF_141.Q ),
    .b(\DFF_177.Q ),
    .c(RESET),
    .y(_00925_)
  );
  al_aoi21ftf _05588_ (
    .a(\DFF_141.Q ),
    .b(\DFF_177.Q ),
    .c(_00925_),
    .y(\DFF_178.D )
  );
  al_oa21ftt _05589_ (
    .a(\DFF_140.Q ),
    .b(\DFF_178.Q ),
    .c(RESET),
    .y(_00926_)
  );
  al_aoi21ftf _05590_ (
    .a(\DFF_140.Q ),
    .b(\DFF_178.Q ),
    .c(_00926_),
    .y(\DFF_179.D )
  );
  al_oa21ftt _05591_ (
    .a(\DFF_139.Q ),
    .b(\DFF_179.Q ),
    .c(RESET),
    .y(_00927_)
  );
  al_aoi21ftf _05592_ (
    .a(\DFF_139.Q ),
    .b(\DFF_179.Q ),
    .c(_00927_),
    .y(\DFF_180.D )
  );
  al_oa21ftt _05593_ (
    .a(\DFF_138.Q ),
    .b(\DFF_180.Q ),
    .c(RESET),
    .y(_00928_)
  );
  al_aoi21ftf _05594_ (
    .a(\DFF_138.Q ),
    .b(\DFF_180.Q ),
    .c(_00928_),
    .y(\DFF_181.D )
  );
  al_oa21ftt _05595_ (
    .a(\DFF_137.Q ),
    .b(\DFF_181.Q ),
    .c(RESET),
    .y(_00929_)
  );
  al_aoi21ftf _05596_ (
    .a(\DFF_137.Q ),
    .b(\DFF_181.Q ),
    .c(_00929_),
    .y(\DFF_182.D )
  );
  al_oa21ftt _05597_ (
    .a(\DFF_136.Q ),
    .b(\DFF_182.Q ),
    .c(RESET),
    .y(_00930_)
  );
  al_aoi21ftf _05598_ (
    .a(\DFF_136.Q ),
    .b(\DFF_182.Q ),
    .c(_00930_),
    .y(\DFF_183.D )
  );
  al_oa21ftt _05599_ (
    .a(\DFF_135.Q ),
    .b(\DFF_183.Q ),
    .c(RESET),
    .y(_00931_)
  );
  al_aoi21ftf _05600_ (
    .a(\DFF_135.Q ),
    .b(\DFF_183.Q ),
    .c(_00931_),
    .y(\DFF_184.D )
  );
  al_oa21ftt _05601_ (
    .a(\DFF_134.Q ),
    .b(\DFF_184.Q ),
    .c(RESET),
    .y(_00932_)
  );
  al_aoi21ftf _05602_ (
    .a(\DFF_134.Q ),
    .b(\DFF_184.Q ),
    .c(_00932_),
    .y(\DFF_185.D )
  );
  al_oa21ftt _05603_ (
    .a(\DFF_133.Q ),
    .b(\DFF_185.Q ),
    .c(RESET),
    .y(_00933_)
  );
  al_aoi21ftf _05604_ (
    .a(\DFF_133.Q ),
    .b(\DFF_185.Q ),
    .c(_00933_),
    .y(\DFF_186.D )
  );
  al_oa21ftt _05605_ (
    .a(\DFF_132.Q ),
    .b(\DFF_186.Q ),
    .c(RESET),
    .y(_00934_)
  );
  al_aoi21ftf _05606_ (
    .a(\DFF_132.Q ),
    .b(\DFF_186.Q ),
    .c(_00934_),
    .y(\DFF_187.D )
  );
  al_oa21ftt _05607_ (
    .a(\DFF_131.Q ),
    .b(\DFF_187.Q ),
    .c(RESET),
    .y(_00935_)
  );
  al_aoi21ftf _05608_ (
    .a(\DFF_131.Q ),
    .b(\DFF_187.Q ),
    .c(_00935_),
    .y(\DFF_188.D )
  );
  al_oa21ftt _05609_ (
    .a(\DFF_130.Q ),
    .b(\DFF_188.Q ),
    .c(RESET),
    .y(_00936_)
  );
  al_aoi21ftf _05610_ (
    .a(\DFF_130.Q ),
    .b(\DFF_188.Q ),
    .c(_00936_),
    .y(\DFF_189.D )
  );
  al_oa21ftt _05611_ (
    .a(\DFF_129.Q ),
    .b(\DFF_189.Q ),
    .c(RESET),
    .y(_00937_)
  );
  al_aoi21ftf _05612_ (
    .a(\DFF_129.Q ),
    .b(\DFF_189.Q ),
    .c(_00937_),
    .y(\DFF_190.D )
  );
  al_oa21ftt _05613_ (
    .a(\DFF_128.Q ),
    .b(\DFF_190.Q ),
    .c(RESET),
    .y(_00938_)
  );
  al_aoi21ftf _05614_ (
    .a(\DFF_128.Q ),
    .b(\DFF_190.Q ),
    .c(_00938_),
    .y(\DFF_191.D )
  );
  al_and2 _05615_ (
    .a(RESET),
    .b(\DFF_193.Q ),
    .y(\DFF_192.D )
  );
  al_and2 _05616_ (
    .a(RESET),
    .b(\DFF_194.Q ),
    .y(\DFF_193.D )
  );
  al_and2 _05617_ (
    .a(RESET),
    .b(\DFF_195.Q ),
    .y(\DFF_194.D )
  );
  al_and2 _05618_ (
    .a(RESET),
    .b(\DFF_196.Q ),
    .y(\DFF_195.D )
  );
  al_and2 _05619_ (
    .a(RESET),
    .b(\DFF_197.Q ),
    .y(\DFF_196.D )
  );
  al_and2 _05620_ (
    .a(RESET),
    .b(\DFF_198.Q ),
    .y(\DFF_197.D )
  );
  al_and2 _05621_ (
    .a(RESET),
    .b(\DFF_199.Q ),
    .y(\DFF_198.D )
  );
  al_and2 _05622_ (
    .a(RESET),
    .b(\DFF_200.Q ),
    .y(\DFF_199.D )
  );
  al_and2 _05623_ (
    .a(RESET),
    .b(\DFF_201.Q ),
    .y(\DFF_200.D )
  );
  al_and2 _05624_ (
    .a(RESET),
    .b(\DFF_202.Q ),
    .y(\DFF_201.D )
  );
  al_and2 _05625_ (
    .a(RESET),
    .b(\DFF_203.Q ),
    .y(\DFF_202.D )
  );
  al_and2 _05626_ (
    .a(RESET),
    .b(\DFF_204.Q ),
    .y(\DFF_203.D )
  );
  al_and2 _05627_ (
    .a(RESET),
    .b(\DFF_205.Q ),
    .y(\DFF_204.D )
  );
  al_and2 _05628_ (
    .a(RESET),
    .b(\DFF_206.Q ),
    .y(\DFF_205.D )
  );
  al_and2 _05629_ (
    .a(RESET),
    .b(\DFF_207.Q ),
    .y(\DFF_206.D )
  );
  al_and2 _05630_ (
    .a(RESET),
    .b(\DFF_208.Q ),
    .y(\DFF_207.D )
  );
  al_and2 _05631_ (
    .a(RESET),
    .b(\DFF_209.Q ),
    .y(\DFF_208.D )
  );
  al_and2 _05632_ (
    .a(RESET),
    .b(\DFF_210.Q ),
    .y(\DFF_209.D )
  );
  al_and2 _05633_ (
    .a(RESET),
    .b(\DFF_211.Q ),
    .y(\DFF_210.D )
  );
  al_and2 _05634_ (
    .a(RESET),
    .b(\DFF_212.Q ),
    .y(\DFF_211.D )
  );
  al_and2 _05635_ (
    .a(RESET),
    .b(\DFF_213.Q ),
    .y(\DFF_212.D )
  );
  al_and2 _05636_ (
    .a(RESET),
    .b(\DFF_214.Q ),
    .y(\DFF_213.D )
  );
  al_and2 _05637_ (
    .a(RESET),
    .b(\DFF_215.Q ),
    .y(\DFF_214.D )
  );
  al_and2 _05638_ (
    .a(RESET),
    .b(\DFF_216.Q ),
    .y(\DFF_215.D )
  );
  al_and2 _05639_ (
    .a(RESET),
    .b(\DFF_217.Q ),
    .y(\DFF_216.D )
  );
  al_and2 _05640_ (
    .a(RESET),
    .b(\DFF_218.Q ),
    .y(\DFF_217.D )
  );
  al_and2 _05641_ (
    .a(RESET),
    .b(\DFF_219.Q ),
    .y(\DFF_218.D )
  );
  al_and2 _05642_ (
    .a(RESET),
    .b(\DFF_220.Q ),
    .y(\DFF_219.D )
  );
  al_and2 _05643_ (
    .a(RESET),
    .b(\DFF_221.Q ),
    .y(\DFF_220.D )
  );
  al_and2 _05644_ (
    .a(RESET),
    .b(\DFF_222.Q ),
    .y(\DFF_221.D )
  );
  al_and2 _05645_ (
    .a(RESET),
    .b(\DFF_223.Q ),
    .y(\DFF_222.D )
  );
  al_and2ft _05646_ (
    .a(\DFF_192.Q ),
    .b(RESET),
    .y(\DFF_223.D )
  );
  al_or2 _05647_ (
    .a(TM1),
    .b(\DFF_480.Q ),
    .y(_00939_)
  );
  al_nand2 _05648_ (
    .a(TM1),
    .b(\DFF_480.Q ),
    .y(_00940_)
  );
  al_nand3 _05649_ (
    .a(\DFF_512.Q ),
    .b(_00939_),
    .c(_00940_),
    .y(_00941_)
  );
  al_nand2ft _05650_ (
    .a(TM1),
    .b(\DFF_480.Q ),
    .y(_00942_)
  );
  al_and2ft _05651_ (
    .a(\DFF_480.Q ),
    .b(TM1),
    .y(_00943_)
  );
  al_and3fft _05652_ (
    .a(\DFF_512.Q ),
    .b(_00943_),
    .c(_00942_),
    .y(_00944_)
  );
  al_and2ft _05653_ (
    .a(\DFF_448.Q ),
    .b(\DFF_416.Q ),
    .y(_00945_)
  );
  al_nand2ft _05654_ (
    .a(\DFF_416.Q ),
    .b(\DFF_448.Q ),
    .y(_00946_)
  );
  al_nand2ft _05655_ (
    .a(_00945_),
    .b(_00946_),
    .y(_00947_)
  );
  al_oai21ftf _05656_ (
    .a(_00941_),
    .b(_00944_),
    .c(_00947_),
    .y(_00948_)
  );
  al_nand3ftt _05657_ (
    .a(_00944_),
    .b(_00941_),
    .c(_00947_),
    .y(_00949_)
  );
  al_nand3 _05658_ (
    .a(_00448_),
    .b(_00948_),
    .c(_00949_),
    .y(_00950_)
  );
  al_ao21 _05659_ (
    .a(TM0),
    .b(\DFF_383.Q ),
    .c(TM1),
    .y(_00951_)
  );
  al_aoi21ttf _05660_ (
    .a(\DFF_192.Q ),
    .b(TM0),
    .c(TM1),
    .y(_00952_)
  );
  al_aoi21 _05661_ (
    .a(_00952_),
    .b(_00463_),
    .c(_00451_),
    .y(_00953_)
  );
  al_aoi21ftf _05662_ (
    .a(_00951_),
    .b(_00950_),
    .c(_00953_),
    .y(\DFF_224.D )
  );
  al_or2 _05663_ (
    .a(TM1),
    .b(\DFF_481.Q ),
    .y(_00954_)
  );
  al_nand2 _05664_ (
    .a(TM1),
    .b(\DFF_481.Q ),
    .y(_00955_)
  );
  al_nand3 _05665_ (
    .a(\DFF_513.Q ),
    .b(_00954_),
    .c(_00955_),
    .y(_00956_)
  );
  al_nand2ft _05666_ (
    .a(TM1),
    .b(\DFF_481.Q ),
    .y(_00957_)
  );
  al_and2ft _05667_ (
    .a(\DFF_481.Q ),
    .b(TM1),
    .y(_00958_)
  );
  al_and3fft _05668_ (
    .a(\DFF_513.Q ),
    .b(_00958_),
    .c(_00957_),
    .y(_00959_)
  );
  al_and2ft _05669_ (
    .a(\DFF_449.Q ),
    .b(\DFF_417.Q ),
    .y(_00960_)
  );
  al_nand2ft _05670_ (
    .a(\DFF_417.Q ),
    .b(\DFF_449.Q ),
    .y(_00961_)
  );
  al_nand2ft _05671_ (
    .a(_00960_),
    .b(_00961_),
    .y(_00962_)
  );
  al_oai21ftf _05672_ (
    .a(_00956_),
    .b(_00959_),
    .c(_00962_),
    .y(_00963_)
  );
  al_nand3ftt _05673_ (
    .a(_00959_),
    .b(_00956_),
    .c(_00962_),
    .y(_00964_)
  );
  al_nand3 _05674_ (
    .a(_00448_),
    .b(_00963_),
    .c(_00964_),
    .y(_00965_)
  );
  al_ao21 _05675_ (
    .a(TM0),
    .b(\DFF_382.Q ),
    .c(TM1),
    .y(_00966_)
  );
  al_aoi21ttf _05676_ (
    .a(TM0),
    .b(\DFF_193.Q ),
    .c(TM1),
    .y(_00967_)
  );
  al_aoi21 _05677_ (
    .a(_00967_),
    .b(_00479_),
    .c(_00451_),
    .y(_00968_)
  );
  al_aoi21ftf _05678_ (
    .a(_00966_),
    .b(_00965_),
    .c(_00968_),
    .y(\DFF_225.D )
  );
  al_or2 _05679_ (
    .a(TM1),
    .b(\DFF_482.Q ),
    .y(_00969_)
  );
  al_nand2 _05680_ (
    .a(TM1),
    .b(\DFF_482.Q ),
    .y(_00970_)
  );
  al_nand3 _05681_ (
    .a(\DFF_514.Q ),
    .b(_00969_),
    .c(_00970_),
    .y(_00971_)
  );
  al_nand2ft _05682_ (
    .a(TM1),
    .b(\DFF_482.Q ),
    .y(_00972_)
  );
  al_and2ft _05683_ (
    .a(\DFF_482.Q ),
    .b(TM1),
    .y(_00973_)
  );
  al_and3fft _05684_ (
    .a(\DFF_514.Q ),
    .b(_00973_),
    .c(_00972_),
    .y(_00974_)
  );
  al_and2ft _05685_ (
    .a(\DFF_450.Q ),
    .b(\DFF_418.Q ),
    .y(_00975_)
  );
  al_nand2ft _05686_ (
    .a(\DFF_418.Q ),
    .b(\DFF_450.Q ),
    .y(_00976_)
  );
  al_nand2ft _05687_ (
    .a(_00975_),
    .b(_00976_),
    .y(_00977_)
  );
  al_oai21ftf _05688_ (
    .a(_00971_),
    .b(_00974_),
    .c(_00977_),
    .y(_00978_)
  );
  al_nand3ftt _05689_ (
    .a(_00974_),
    .b(_00971_),
    .c(_00977_),
    .y(_00979_)
  );
  al_nand3 _05690_ (
    .a(_00448_),
    .b(_00978_),
    .c(_00979_),
    .y(_00980_)
  );
  al_ao21 _05691_ (
    .a(TM0),
    .b(\DFF_381.Q ),
    .c(TM1),
    .y(_00981_)
  );
  al_aoi21ttf _05692_ (
    .a(TM0),
    .b(\DFF_194.Q ),
    .c(TM1),
    .y(_00982_)
  );
  al_aoi21 _05693_ (
    .a(_00982_),
    .b(_00495_),
    .c(_00451_),
    .y(_00983_)
  );
  al_aoi21ftf _05694_ (
    .a(_00981_),
    .b(_00980_),
    .c(_00983_),
    .y(\DFF_226.D )
  );
  al_or2 _05695_ (
    .a(TM1),
    .b(\DFF_483.Q ),
    .y(_00984_)
  );
  al_nand2 _05696_ (
    .a(TM1),
    .b(\DFF_483.Q ),
    .y(_00985_)
  );
  al_nand3 _05697_ (
    .a(\DFF_515.Q ),
    .b(_00984_),
    .c(_00985_),
    .y(_00986_)
  );
  al_nand2ft _05698_ (
    .a(TM1),
    .b(\DFF_483.Q ),
    .y(_00987_)
  );
  al_and2ft _05699_ (
    .a(\DFF_483.Q ),
    .b(TM1),
    .y(_00988_)
  );
  al_and3fft _05700_ (
    .a(\DFF_515.Q ),
    .b(_00988_),
    .c(_00987_),
    .y(_00989_)
  );
  al_and2ft _05701_ (
    .a(\DFF_451.Q ),
    .b(\DFF_419.Q ),
    .y(_00990_)
  );
  al_nand2ft _05702_ (
    .a(\DFF_419.Q ),
    .b(\DFF_451.Q ),
    .y(_00991_)
  );
  al_nand2ft _05703_ (
    .a(_00990_),
    .b(_00991_),
    .y(_00992_)
  );
  al_oai21ftf _05704_ (
    .a(_00986_),
    .b(_00989_),
    .c(_00992_),
    .y(_00993_)
  );
  al_nand3ftt _05705_ (
    .a(_00989_),
    .b(_00986_),
    .c(_00992_),
    .y(_00994_)
  );
  al_nand3 _05706_ (
    .a(_00448_),
    .b(_00993_),
    .c(_00994_),
    .y(_00995_)
  );
  al_ao21 _05707_ (
    .a(TM0),
    .b(\DFF_380.Q ),
    .c(TM1),
    .y(_00996_)
  );
  al_aoi21ttf _05708_ (
    .a(TM0),
    .b(\DFF_195.Q ),
    .c(TM1),
    .y(_00997_)
  );
  al_aoi21 _05709_ (
    .a(_00997_),
    .b(_00511_),
    .c(_00451_),
    .y(_00998_)
  );
  al_aoi21ftf _05710_ (
    .a(_00996_),
    .b(_00995_),
    .c(_00998_),
    .y(\DFF_227.D )
  );
  al_or2 _05711_ (
    .a(TM1),
    .b(\DFF_484.Q ),
    .y(_00999_)
  );
  al_nand2 _05712_ (
    .a(TM1),
    .b(\DFF_484.Q ),
    .y(_01000_)
  );
  al_nand3 _05713_ (
    .a(\DFF_516.Q ),
    .b(_00999_),
    .c(_01000_),
    .y(_01001_)
  );
  al_nand2ft _05714_ (
    .a(TM1),
    .b(\DFF_484.Q ),
    .y(_01002_)
  );
  al_and2ft _05715_ (
    .a(\DFF_484.Q ),
    .b(TM1),
    .y(_01003_)
  );
  al_and3fft _05716_ (
    .a(\DFF_516.Q ),
    .b(_01003_),
    .c(_01002_),
    .y(_01004_)
  );
  al_and2ft _05717_ (
    .a(\DFF_452.Q ),
    .b(\DFF_420.Q ),
    .y(_01005_)
  );
  al_nand2ft _05718_ (
    .a(\DFF_420.Q ),
    .b(\DFF_452.Q ),
    .y(_01006_)
  );
  al_nand2ft _05719_ (
    .a(_01005_),
    .b(_01006_),
    .y(_01007_)
  );
  al_oai21ftf _05720_ (
    .a(_01001_),
    .b(_01004_),
    .c(_01007_),
    .y(_01008_)
  );
  al_nand3ftt _05721_ (
    .a(_01004_),
    .b(_01001_),
    .c(_01007_),
    .y(_01009_)
  );
  al_nand3 _05722_ (
    .a(_00448_),
    .b(_01008_),
    .c(_01009_),
    .y(_01010_)
  );
  al_ao21 _05723_ (
    .a(TM0),
    .b(\DFF_379.Q ),
    .c(TM1),
    .y(_01011_)
  );
  al_aoi21ttf _05724_ (
    .a(TM0),
    .b(\DFF_196.Q ),
    .c(TM1),
    .y(_01012_)
  );
  al_aoi21 _05725_ (
    .a(_01012_),
    .b(_00527_),
    .c(_00451_),
    .y(_01013_)
  );
  al_aoi21ftf _05726_ (
    .a(_01011_),
    .b(_01010_),
    .c(_01013_),
    .y(\DFF_228.D )
  );
  al_or2 _05727_ (
    .a(TM1),
    .b(\DFF_485.Q ),
    .y(_01014_)
  );
  al_nand2 _05728_ (
    .a(TM1),
    .b(\DFF_485.Q ),
    .y(_01015_)
  );
  al_nand3 _05729_ (
    .a(\DFF_517.Q ),
    .b(_01014_),
    .c(_01015_),
    .y(_01016_)
  );
  al_nand2ft _05730_ (
    .a(TM1),
    .b(\DFF_485.Q ),
    .y(_01017_)
  );
  al_and2ft _05731_ (
    .a(\DFF_485.Q ),
    .b(TM1),
    .y(_01018_)
  );
  al_and3fft _05732_ (
    .a(\DFF_517.Q ),
    .b(_01018_),
    .c(_01017_),
    .y(_01019_)
  );
  al_and2ft _05733_ (
    .a(\DFF_453.Q ),
    .b(\DFF_421.Q ),
    .y(_01020_)
  );
  al_nand2ft _05734_ (
    .a(\DFF_421.Q ),
    .b(\DFF_453.Q ),
    .y(_01021_)
  );
  al_nand2ft _05735_ (
    .a(_01020_),
    .b(_01021_),
    .y(_01022_)
  );
  al_oai21ftf _05736_ (
    .a(_01016_),
    .b(_01019_),
    .c(_01022_),
    .y(_01023_)
  );
  al_nand3ftt _05737_ (
    .a(_01019_),
    .b(_01016_),
    .c(_01022_),
    .y(_01024_)
  );
  al_nand3 _05738_ (
    .a(_00448_),
    .b(_01023_),
    .c(_01024_),
    .y(_01025_)
  );
  al_ao21 _05739_ (
    .a(TM0),
    .b(\DFF_378.Q ),
    .c(TM1),
    .y(_01026_)
  );
  al_aoi21ttf _05740_ (
    .a(TM0),
    .b(\DFF_197.Q ),
    .c(TM1),
    .y(_01027_)
  );
  al_aoi21 _05741_ (
    .a(_01027_),
    .b(_00543_),
    .c(_00451_),
    .y(_01028_)
  );
  al_aoi21ftf _05742_ (
    .a(_01026_),
    .b(_01025_),
    .c(_01028_),
    .y(\DFF_229.D )
  );
  al_or2 _05743_ (
    .a(TM1),
    .b(\DFF_486.Q ),
    .y(_01029_)
  );
  al_nand2 _05744_ (
    .a(TM1),
    .b(\DFF_486.Q ),
    .y(_01030_)
  );
  al_nand3 _05745_ (
    .a(\DFF_518.Q ),
    .b(_01029_),
    .c(_01030_),
    .y(_01031_)
  );
  al_nand2ft _05746_ (
    .a(TM1),
    .b(\DFF_486.Q ),
    .y(_01032_)
  );
  al_and2ft _05747_ (
    .a(\DFF_486.Q ),
    .b(TM1),
    .y(_01033_)
  );
  al_and3fft _05748_ (
    .a(\DFF_518.Q ),
    .b(_01033_),
    .c(_01032_),
    .y(_01034_)
  );
  al_and2ft _05749_ (
    .a(\DFF_454.Q ),
    .b(\DFF_422.Q ),
    .y(_01035_)
  );
  al_nand2ft _05750_ (
    .a(\DFF_422.Q ),
    .b(\DFF_454.Q ),
    .y(_01036_)
  );
  al_nand2ft _05751_ (
    .a(_01035_),
    .b(_01036_),
    .y(_01037_)
  );
  al_oai21ftf _05752_ (
    .a(_01031_),
    .b(_01034_),
    .c(_01037_),
    .y(_01038_)
  );
  al_nand3ftt _05753_ (
    .a(_01034_),
    .b(_01031_),
    .c(_01037_),
    .y(_01039_)
  );
  al_nand3 _05754_ (
    .a(_00448_),
    .b(_01038_),
    .c(_01039_),
    .y(_01040_)
  );
  al_ao21 _05755_ (
    .a(TM0),
    .b(\DFF_377.Q ),
    .c(TM1),
    .y(_01041_)
  );
  al_aoi21ttf _05756_ (
    .a(TM0),
    .b(\DFF_198.Q ),
    .c(TM1),
    .y(_01042_)
  );
  al_aoi21 _05757_ (
    .a(_01042_),
    .b(_00559_),
    .c(_00451_),
    .y(_01043_)
  );
  al_aoi21ftf _05758_ (
    .a(_01041_),
    .b(_01040_),
    .c(_01043_),
    .y(\DFF_230.D )
  );
  al_or2 _05759_ (
    .a(TM1),
    .b(\DFF_487.Q ),
    .y(_01044_)
  );
  al_nand2 _05760_ (
    .a(TM1),
    .b(\DFF_487.Q ),
    .y(_01045_)
  );
  al_nand3 _05761_ (
    .a(\DFF_519.Q ),
    .b(_01044_),
    .c(_01045_),
    .y(_01046_)
  );
  al_nand2ft _05762_ (
    .a(TM1),
    .b(\DFF_487.Q ),
    .y(_01047_)
  );
  al_and2ft _05763_ (
    .a(\DFF_487.Q ),
    .b(TM1),
    .y(_01048_)
  );
  al_and3fft _05764_ (
    .a(\DFF_519.Q ),
    .b(_01048_),
    .c(_01047_),
    .y(_01049_)
  );
  al_and2ft _05765_ (
    .a(\DFF_455.Q ),
    .b(\DFF_423.Q ),
    .y(_01050_)
  );
  al_nand2ft _05766_ (
    .a(\DFF_423.Q ),
    .b(\DFF_455.Q ),
    .y(_01051_)
  );
  al_nand2ft _05767_ (
    .a(_01050_),
    .b(_01051_),
    .y(_01052_)
  );
  al_oai21ftf _05768_ (
    .a(_01046_),
    .b(_01049_),
    .c(_01052_),
    .y(_01053_)
  );
  al_nand3ftt _05769_ (
    .a(_01049_),
    .b(_01046_),
    .c(_01052_),
    .y(_01054_)
  );
  al_nand3 _05770_ (
    .a(_00448_),
    .b(_01053_),
    .c(_01054_),
    .y(_01055_)
  );
  al_ao21 _05771_ (
    .a(TM0),
    .b(\DFF_376.Q ),
    .c(TM1),
    .y(_01056_)
  );
  al_aoi21ttf _05772_ (
    .a(TM0),
    .b(\DFF_199.Q ),
    .c(TM1),
    .y(_01057_)
  );
  al_aoi21 _05773_ (
    .a(_01057_),
    .b(_00575_),
    .c(_00451_),
    .y(_01058_)
  );
  al_aoi21ftf _05774_ (
    .a(_01056_),
    .b(_01055_),
    .c(_01058_),
    .y(\DFF_231.D )
  );
  al_or2 _05775_ (
    .a(TM1),
    .b(\DFF_488.Q ),
    .y(_01059_)
  );
  al_nand2 _05776_ (
    .a(TM1),
    .b(\DFF_488.Q ),
    .y(_01060_)
  );
  al_nand3 _05777_ (
    .a(\DFF_520.Q ),
    .b(_01059_),
    .c(_01060_),
    .y(_01061_)
  );
  al_nand2ft _05778_ (
    .a(TM1),
    .b(\DFF_488.Q ),
    .y(_01062_)
  );
  al_and2ft _05779_ (
    .a(\DFF_488.Q ),
    .b(TM1),
    .y(_01063_)
  );
  al_and3fft _05780_ (
    .a(\DFF_520.Q ),
    .b(_01063_),
    .c(_01062_),
    .y(_01064_)
  );
  al_and2ft _05781_ (
    .a(\DFF_456.Q ),
    .b(\DFF_424.Q ),
    .y(_01065_)
  );
  al_nand2ft _05782_ (
    .a(\DFF_424.Q ),
    .b(\DFF_456.Q ),
    .y(_01066_)
  );
  al_nand2ft _05783_ (
    .a(_01065_),
    .b(_01066_),
    .y(_01067_)
  );
  al_oai21ftf _05784_ (
    .a(_01061_),
    .b(_01064_),
    .c(_01067_),
    .y(_01068_)
  );
  al_nand3ftt _05785_ (
    .a(_01064_),
    .b(_01061_),
    .c(_01067_),
    .y(_01069_)
  );
  al_nand3 _05786_ (
    .a(_00448_),
    .b(_01068_),
    .c(_01069_),
    .y(_01070_)
  );
  al_ao21 _05787_ (
    .a(TM0),
    .b(\DFF_375.Q ),
    .c(TM1),
    .y(_01071_)
  );
  al_aoi21ttf _05788_ (
    .a(TM0),
    .b(\DFF_200.Q ),
    .c(TM1),
    .y(_01072_)
  );
  al_aoi21 _05789_ (
    .a(_01072_),
    .b(_00591_),
    .c(_00451_),
    .y(_01073_)
  );
  al_aoi21ftf _05790_ (
    .a(_01071_),
    .b(_01070_),
    .c(_01073_),
    .y(\DFF_232.D )
  );
  al_or2 _05791_ (
    .a(TM1),
    .b(\DFF_489.Q ),
    .y(_01074_)
  );
  al_nand2 _05792_ (
    .a(TM1),
    .b(\DFF_489.Q ),
    .y(_01075_)
  );
  al_nand3 _05793_ (
    .a(\DFF_521.Q ),
    .b(_01074_),
    .c(_01075_),
    .y(_01076_)
  );
  al_nand2ft _05794_ (
    .a(TM1),
    .b(\DFF_489.Q ),
    .y(_01077_)
  );
  al_and2ft _05795_ (
    .a(\DFF_489.Q ),
    .b(TM1),
    .y(_01078_)
  );
  al_and3fft _05796_ (
    .a(\DFF_521.Q ),
    .b(_01078_),
    .c(_01077_),
    .y(_01079_)
  );
  al_and2ft _05797_ (
    .a(\DFF_457.Q ),
    .b(\DFF_425.Q ),
    .y(_01080_)
  );
  al_nand2ft _05798_ (
    .a(\DFF_425.Q ),
    .b(\DFF_457.Q ),
    .y(_01081_)
  );
  al_nand2ft _05799_ (
    .a(_01080_),
    .b(_01081_),
    .y(_01082_)
  );
  al_oai21ftf _05800_ (
    .a(_01076_),
    .b(_01079_),
    .c(_01082_),
    .y(_01083_)
  );
  al_nand3ftt _05801_ (
    .a(_01079_),
    .b(_01076_),
    .c(_01082_),
    .y(_01084_)
  );
  al_nand3 _05802_ (
    .a(_00448_),
    .b(_01083_),
    .c(_01084_),
    .y(_01085_)
  );
  al_ao21 _05803_ (
    .a(TM0),
    .b(\DFF_374.Q ),
    .c(TM1),
    .y(_01086_)
  );
  al_aoi21ttf _05804_ (
    .a(TM0),
    .b(\DFF_201.Q ),
    .c(TM1),
    .y(_01087_)
  );
  al_aoi21 _05805_ (
    .a(_01087_),
    .b(_00607_),
    .c(_00451_),
    .y(_01088_)
  );
  al_aoi21ftf _05806_ (
    .a(_01086_),
    .b(_01085_),
    .c(_01088_),
    .y(\DFF_233.D )
  );
  al_or2 _05807_ (
    .a(TM1),
    .b(\DFF_490.Q ),
    .y(_01089_)
  );
  al_nand2 _05808_ (
    .a(TM1),
    .b(\DFF_490.Q ),
    .y(_01090_)
  );
  al_nand3 _05809_ (
    .a(\DFF_522.Q ),
    .b(_01089_),
    .c(_01090_),
    .y(_01091_)
  );
  al_nand2ft _05810_ (
    .a(TM1),
    .b(\DFF_490.Q ),
    .y(_01092_)
  );
  al_and2ft _05811_ (
    .a(\DFF_490.Q ),
    .b(TM1),
    .y(_01093_)
  );
  al_and3fft _05812_ (
    .a(\DFF_522.Q ),
    .b(_01093_),
    .c(_01092_),
    .y(_01094_)
  );
  al_and2ft _05813_ (
    .a(\DFF_458.Q ),
    .b(\DFF_426.Q ),
    .y(_01095_)
  );
  al_nand2ft _05814_ (
    .a(\DFF_426.Q ),
    .b(\DFF_458.Q ),
    .y(_01096_)
  );
  al_nand2ft _05815_ (
    .a(_01095_),
    .b(_01096_),
    .y(_01097_)
  );
  al_oai21ftf _05816_ (
    .a(_01091_),
    .b(_01094_),
    .c(_01097_),
    .y(_01098_)
  );
  al_nand3ftt _05817_ (
    .a(_01094_),
    .b(_01091_),
    .c(_01097_),
    .y(_01099_)
  );
  al_nand3 _05818_ (
    .a(_00448_),
    .b(_01098_),
    .c(_01099_),
    .y(_01100_)
  );
  al_ao21 _05819_ (
    .a(TM0),
    .b(\DFF_373.Q ),
    .c(TM1),
    .y(_01101_)
  );
  al_aoi21ttf _05820_ (
    .a(TM0),
    .b(\DFF_202.Q ),
    .c(TM1),
    .y(_01102_)
  );
  al_aoi21 _05821_ (
    .a(_01102_),
    .b(_00623_),
    .c(_00451_),
    .y(_01103_)
  );
  al_aoi21ftf _05822_ (
    .a(_01101_),
    .b(_01100_),
    .c(_01103_),
    .y(\DFF_234.D )
  );
  al_or2 _05823_ (
    .a(TM1),
    .b(\DFF_491.Q ),
    .y(_01104_)
  );
  al_nand2 _05824_ (
    .a(TM1),
    .b(\DFF_491.Q ),
    .y(_01105_)
  );
  al_nand3 _05825_ (
    .a(\DFF_523.Q ),
    .b(_01104_),
    .c(_01105_),
    .y(_01106_)
  );
  al_nand2ft _05826_ (
    .a(TM1),
    .b(\DFF_491.Q ),
    .y(_01107_)
  );
  al_and2ft _05827_ (
    .a(\DFF_491.Q ),
    .b(TM1),
    .y(_01108_)
  );
  al_and3fft _05828_ (
    .a(\DFF_523.Q ),
    .b(_01108_),
    .c(_01107_),
    .y(_01109_)
  );
  al_and2ft _05829_ (
    .a(\DFF_459.Q ),
    .b(\DFF_427.Q ),
    .y(_01110_)
  );
  al_nand2ft _05830_ (
    .a(\DFF_427.Q ),
    .b(\DFF_459.Q ),
    .y(_01111_)
  );
  al_nand2ft _05831_ (
    .a(_01110_),
    .b(_01111_),
    .y(_01112_)
  );
  al_oai21ftf _05832_ (
    .a(_01106_),
    .b(_01109_),
    .c(_01112_),
    .y(_01113_)
  );
  al_nand3ftt _05833_ (
    .a(_01109_),
    .b(_01106_),
    .c(_01112_),
    .y(_01114_)
  );
  al_nand3 _05834_ (
    .a(_00448_),
    .b(_01113_),
    .c(_01114_),
    .y(_01115_)
  );
  al_ao21 _05835_ (
    .a(TM0),
    .b(\DFF_372.Q ),
    .c(TM1),
    .y(_01116_)
  );
  al_aoi21ttf _05836_ (
    .a(TM0),
    .b(\DFF_203.Q ),
    .c(TM1),
    .y(_01117_)
  );
  al_aoi21 _05837_ (
    .a(_01117_),
    .b(_00639_),
    .c(_00451_),
    .y(_01118_)
  );
  al_aoi21ftf _05838_ (
    .a(_01116_),
    .b(_01115_),
    .c(_01118_),
    .y(\DFF_235.D )
  );
  al_or2 _05839_ (
    .a(TM1),
    .b(\DFF_492.Q ),
    .y(_01119_)
  );
  al_nand2 _05840_ (
    .a(TM1),
    .b(\DFF_492.Q ),
    .y(_01120_)
  );
  al_nand3 _05841_ (
    .a(\DFF_524.Q ),
    .b(_01119_),
    .c(_01120_),
    .y(_01121_)
  );
  al_nand2ft _05842_ (
    .a(TM1),
    .b(\DFF_492.Q ),
    .y(_01122_)
  );
  al_and2ft _05843_ (
    .a(\DFF_492.Q ),
    .b(TM1),
    .y(_01123_)
  );
  al_and3fft _05844_ (
    .a(\DFF_524.Q ),
    .b(_01123_),
    .c(_01122_),
    .y(_01124_)
  );
  al_and2ft _05845_ (
    .a(\DFF_460.Q ),
    .b(\DFF_428.Q ),
    .y(_01125_)
  );
  al_nand2ft _05846_ (
    .a(\DFF_428.Q ),
    .b(\DFF_460.Q ),
    .y(_01126_)
  );
  al_nand2ft _05847_ (
    .a(_01125_),
    .b(_01126_),
    .y(_01127_)
  );
  al_oai21ftf _05848_ (
    .a(_01121_),
    .b(_01124_),
    .c(_01127_),
    .y(_01128_)
  );
  al_nand3ftt _05849_ (
    .a(_01124_),
    .b(_01121_),
    .c(_01127_),
    .y(_01129_)
  );
  al_nand3 _05850_ (
    .a(_00448_),
    .b(_01128_),
    .c(_01129_),
    .y(_01130_)
  );
  al_ao21 _05851_ (
    .a(TM0),
    .b(\DFF_371.Q ),
    .c(TM1),
    .y(_01131_)
  );
  al_aoi21ttf _05852_ (
    .a(TM0),
    .b(\DFF_204.Q ),
    .c(TM1),
    .y(_01132_)
  );
  al_aoi21 _05853_ (
    .a(_01132_),
    .b(_00655_),
    .c(_00451_),
    .y(_01133_)
  );
  al_aoi21ftf _05854_ (
    .a(_01131_),
    .b(_01130_),
    .c(_01133_),
    .y(\DFF_236.D )
  );
  al_or2 _05855_ (
    .a(TM1),
    .b(\DFF_493.Q ),
    .y(_01134_)
  );
  al_nand2 _05856_ (
    .a(TM1),
    .b(\DFF_493.Q ),
    .y(_01135_)
  );
  al_nand3 _05857_ (
    .a(\DFF_525.Q ),
    .b(_01134_),
    .c(_01135_),
    .y(_01136_)
  );
  al_nand2ft _05858_ (
    .a(TM1),
    .b(\DFF_493.Q ),
    .y(_01137_)
  );
  al_and2ft _05859_ (
    .a(\DFF_493.Q ),
    .b(TM1),
    .y(_01138_)
  );
  al_and3fft _05860_ (
    .a(\DFF_525.Q ),
    .b(_01138_),
    .c(_01137_),
    .y(_01139_)
  );
  al_and2ft _05861_ (
    .a(\DFF_461.Q ),
    .b(\DFF_429.Q ),
    .y(_01140_)
  );
  al_nand2ft _05862_ (
    .a(\DFF_429.Q ),
    .b(\DFF_461.Q ),
    .y(_01141_)
  );
  al_nand2ft _05863_ (
    .a(_01140_),
    .b(_01141_),
    .y(_01142_)
  );
  al_oai21ftf _05864_ (
    .a(_01136_),
    .b(_01139_),
    .c(_01142_),
    .y(_01143_)
  );
  al_nand3ftt _05865_ (
    .a(_01139_),
    .b(_01136_),
    .c(_01142_),
    .y(_01144_)
  );
  al_nand3 _05866_ (
    .a(_00448_),
    .b(_01143_),
    .c(_01144_),
    .y(_01145_)
  );
  al_ao21 _05867_ (
    .a(TM0),
    .b(\DFF_370.Q ),
    .c(TM1),
    .y(_01146_)
  );
  al_aoi21ttf _05868_ (
    .a(TM0),
    .b(\DFF_205.Q ),
    .c(TM1),
    .y(_01147_)
  );
  al_aoi21 _05869_ (
    .a(_01147_),
    .b(_00671_),
    .c(_00451_),
    .y(_01148_)
  );
  al_aoi21ftf _05870_ (
    .a(_01146_),
    .b(_01145_),
    .c(_01148_),
    .y(\DFF_237.D )
  );
  al_or2 _05871_ (
    .a(TM1),
    .b(\DFF_494.Q ),
    .y(_01149_)
  );
  al_nand2 _05872_ (
    .a(TM1),
    .b(\DFF_494.Q ),
    .y(_01150_)
  );
  al_nand3 _05873_ (
    .a(\DFF_526.Q ),
    .b(_01149_),
    .c(_01150_),
    .y(_01151_)
  );
  al_nand2ft _05874_ (
    .a(TM1),
    .b(\DFF_494.Q ),
    .y(_01152_)
  );
  al_and2ft _05875_ (
    .a(\DFF_494.Q ),
    .b(TM1),
    .y(_01153_)
  );
  al_and3fft _05876_ (
    .a(\DFF_526.Q ),
    .b(_01153_),
    .c(_01152_),
    .y(_01154_)
  );
  al_and2ft _05877_ (
    .a(\DFF_462.Q ),
    .b(\DFF_430.Q ),
    .y(_01155_)
  );
  al_nand2ft _05878_ (
    .a(\DFF_430.Q ),
    .b(\DFF_462.Q ),
    .y(_01156_)
  );
  al_nand2ft _05879_ (
    .a(_01155_),
    .b(_01156_),
    .y(_01157_)
  );
  al_oai21ftf _05880_ (
    .a(_01151_),
    .b(_01154_),
    .c(_01157_),
    .y(_01158_)
  );
  al_nand3ftt _05881_ (
    .a(_01154_),
    .b(_01151_),
    .c(_01157_),
    .y(_01159_)
  );
  al_nand3 _05882_ (
    .a(_00448_),
    .b(_01158_),
    .c(_01159_),
    .y(_01160_)
  );
  al_ao21 _05883_ (
    .a(TM0),
    .b(\DFF_369.Q ),
    .c(TM1),
    .y(_01161_)
  );
  al_aoi21ttf _05884_ (
    .a(TM0),
    .b(\DFF_206.Q ),
    .c(TM1),
    .y(_01162_)
  );
  al_aoi21 _05885_ (
    .a(_01162_),
    .b(_00687_),
    .c(_00451_),
    .y(_01163_)
  );
  al_aoi21ftf _05886_ (
    .a(_01161_),
    .b(_01160_),
    .c(_01163_),
    .y(\DFF_238.D )
  );
  al_or2 _05887_ (
    .a(TM1),
    .b(\DFF_495.Q ),
    .y(_01164_)
  );
  al_nand2 _05888_ (
    .a(TM1),
    .b(\DFF_495.Q ),
    .y(_01165_)
  );
  al_nand3 _05889_ (
    .a(\DFF_527.Q ),
    .b(_01164_),
    .c(_01165_),
    .y(_01166_)
  );
  al_nand2ft _05890_ (
    .a(TM1),
    .b(\DFF_495.Q ),
    .y(_01167_)
  );
  al_and2ft _05891_ (
    .a(\DFF_495.Q ),
    .b(TM1),
    .y(_01168_)
  );
  al_and3fft _05892_ (
    .a(\DFF_527.Q ),
    .b(_01168_),
    .c(_01167_),
    .y(_01169_)
  );
  al_and2ft _05893_ (
    .a(\DFF_463.Q ),
    .b(\DFF_431.Q ),
    .y(_01170_)
  );
  al_nand2ft _05894_ (
    .a(\DFF_431.Q ),
    .b(\DFF_463.Q ),
    .y(_01171_)
  );
  al_nand2ft _05895_ (
    .a(_01170_),
    .b(_01171_),
    .y(_01172_)
  );
  al_oai21ftf _05896_ (
    .a(_01166_),
    .b(_01169_),
    .c(_01172_),
    .y(_01173_)
  );
  al_nand3ftt _05897_ (
    .a(_01169_),
    .b(_01166_),
    .c(_01172_),
    .y(_01174_)
  );
  al_nand3 _05898_ (
    .a(_00448_),
    .b(_01173_),
    .c(_01174_),
    .y(_01175_)
  );
  al_ao21 _05899_ (
    .a(TM0),
    .b(\DFF_368.Q ),
    .c(TM1),
    .y(_01176_)
  );
  al_aoi21ttf _05900_ (
    .a(TM0),
    .b(\DFF_207.Q ),
    .c(TM1),
    .y(_01177_)
  );
  al_aoi21 _05901_ (
    .a(_01177_),
    .b(_00703_),
    .c(_00451_),
    .y(_01178_)
  );
  al_aoi21ftf _05902_ (
    .a(_01176_),
    .b(_01175_),
    .c(_01178_),
    .y(\DFF_239.D )
  );
  al_nor2 _05903_ (
    .a(\DFF_464.Q ),
    .b(\DFF_496.Q ),
    .y(_01179_)
  );
  al_and2 _05904_ (
    .a(\DFF_464.Q ),
    .b(\DFF_496.Q ),
    .y(_01180_)
  );
  al_and2ft _05905_ (
    .a(\DFF_432.Q ),
    .b(\DFF_528.Q ),
    .y(_01181_)
  );
  al_nand2ft _05906_ (
    .a(\DFF_528.Q ),
    .b(\DFF_432.Q ),
    .y(_01182_)
  );
  al_nand2ft _05907_ (
    .a(_01181_),
    .b(_01182_),
    .y(_01183_)
  );
  al_oa21ttf _05908_ (
    .a(_01179_),
    .b(_01180_),
    .c(_01183_),
    .y(_01184_)
  );
  al_nand3fft _05909_ (
    .a(_01179_),
    .b(_01180_),
    .c(_01183_),
    .y(_01185_)
  );
  al_and3fft _05910_ (
    .a(TM0),
    .b(_01184_),
    .c(_01185_),
    .y(_01186_)
  );
  al_aoi21 _05911_ (
    .a(TM0),
    .b(\DFF_367.Q ),
    .c(TM1),
    .y(_01187_)
  );
  al_aoi21ttf _05912_ (
    .a(TM0),
    .b(\DFF_208.Q ),
    .c(TM1),
    .y(_01188_)
  );
  al_aoi21 _05913_ (
    .a(_01188_),
    .b(_00715_),
    .c(_00451_),
    .y(_01189_)
  );
  al_aoi21ftf _05914_ (
    .a(_01186_),
    .b(_01187_),
    .c(_01189_),
    .y(\DFF_240.D )
  );
  al_nor2 _05915_ (
    .a(\DFF_465.Q ),
    .b(\DFF_497.Q ),
    .y(_01190_)
  );
  al_and2 _05916_ (
    .a(\DFF_465.Q ),
    .b(\DFF_497.Q ),
    .y(_01191_)
  );
  al_and2ft _05917_ (
    .a(\DFF_433.Q ),
    .b(\DFF_529.Q ),
    .y(_01192_)
  );
  al_nand2ft _05918_ (
    .a(\DFF_529.Q ),
    .b(\DFF_433.Q ),
    .y(_01193_)
  );
  al_nand2ft _05919_ (
    .a(_01192_),
    .b(_01193_),
    .y(_01194_)
  );
  al_oa21ttf _05920_ (
    .a(_01190_),
    .b(_01191_),
    .c(_01194_),
    .y(_01195_)
  );
  al_nand3fft _05921_ (
    .a(_01190_),
    .b(_01191_),
    .c(_01194_),
    .y(_01196_)
  );
  al_and3fft _05922_ (
    .a(TM0),
    .b(_01195_),
    .c(_01196_),
    .y(_01197_)
  );
  al_aoi21 _05923_ (
    .a(TM0),
    .b(\DFF_366.Q ),
    .c(TM1),
    .y(_01198_)
  );
  al_aoi21ttf _05924_ (
    .a(TM0),
    .b(\DFF_209.Q ),
    .c(TM1),
    .y(_01199_)
  );
  al_aoi21 _05925_ (
    .a(_01199_),
    .b(_00727_),
    .c(_00451_),
    .y(_01200_)
  );
  al_aoi21ftf _05926_ (
    .a(_01197_),
    .b(_01198_),
    .c(_01200_),
    .y(\DFF_241.D )
  );
  al_nor2 _05927_ (
    .a(\DFF_466.Q ),
    .b(\DFF_498.Q ),
    .y(_01201_)
  );
  al_and2 _05928_ (
    .a(\DFF_466.Q ),
    .b(\DFF_498.Q ),
    .y(_01202_)
  );
  al_and2ft _05929_ (
    .a(\DFF_434.Q ),
    .b(\DFF_530.Q ),
    .y(_01203_)
  );
  al_nand2ft _05930_ (
    .a(\DFF_530.Q ),
    .b(\DFF_434.Q ),
    .y(_01204_)
  );
  al_nand2ft _05931_ (
    .a(_01203_),
    .b(_01204_),
    .y(_01205_)
  );
  al_oa21ttf _05932_ (
    .a(_01201_),
    .b(_01202_),
    .c(_01205_),
    .y(_01206_)
  );
  al_nand3fft _05933_ (
    .a(_01201_),
    .b(_01202_),
    .c(_01205_),
    .y(_01207_)
  );
  al_and3fft _05934_ (
    .a(TM0),
    .b(_01206_),
    .c(_01207_),
    .y(_01208_)
  );
  al_aoi21 _05935_ (
    .a(TM0),
    .b(\DFF_365.Q ),
    .c(TM1),
    .y(_01209_)
  );
  al_aoi21ttf _05936_ (
    .a(TM0),
    .b(\DFF_210.Q ),
    .c(TM1),
    .y(_01210_)
  );
  al_aoi21 _05937_ (
    .a(_01210_),
    .b(_00739_),
    .c(_00451_),
    .y(_01211_)
  );
  al_aoi21ftf _05938_ (
    .a(_01208_),
    .b(_01209_),
    .c(_01211_),
    .y(\DFF_242.D )
  );
  al_nor2 _05939_ (
    .a(\DFF_467.Q ),
    .b(\DFF_499.Q ),
    .y(_01212_)
  );
  al_and2 _05940_ (
    .a(\DFF_467.Q ),
    .b(\DFF_499.Q ),
    .y(_01213_)
  );
  al_and2ft _05941_ (
    .a(\DFF_435.Q ),
    .b(\DFF_531.Q ),
    .y(_01214_)
  );
  al_nand2ft _05942_ (
    .a(\DFF_531.Q ),
    .b(\DFF_435.Q ),
    .y(_01215_)
  );
  al_nand2ft _05943_ (
    .a(_01214_),
    .b(_01215_),
    .y(_01216_)
  );
  al_oa21ttf _05944_ (
    .a(_01212_),
    .b(_01213_),
    .c(_01216_),
    .y(_01217_)
  );
  al_nand3fft _05945_ (
    .a(_01212_),
    .b(_01213_),
    .c(_01216_),
    .y(_01218_)
  );
  al_and3fft _05946_ (
    .a(TM0),
    .b(_01217_),
    .c(_01218_),
    .y(_01219_)
  );
  al_aoi21 _05947_ (
    .a(TM0),
    .b(\DFF_364.Q ),
    .c(TM1),
    .y(_01220_)
  );
  al_aoi21ttf _05948_ (
    .a(TM0),
    .b(\DFF_211.Q ),
    .c(TM1),
    .y(_01221_)
  );
  al_aoi21 _05949_ (
    .a(_01221_),
    .b(_00751_),
    .c(_00451_),
    .y(_01222_)
  );
  al_aoi21ftf _05950_ (
    .a(_01219_),
    .b(_01220_),
    .c(_01222_),
    .y(\DFF_243.D )
  );
  al_nor2 _05951_ (
    .a(\DFF_468.Q ),
    .b(\DFF_500.Q ),
    .y(_01223_)
  );
  al_and2 _05952_ (
    .a(\DFF_468.Q ),
    .b(\DFF_500.Q ),
    .y(_01224_)
  );
  al_and2ft _05953_ (
    .a(\DFF_436.Q ),
    .b(\DFF_532.Q ),
    .y(_01225_)
  );
  al_nand2ft _05954_ (
    .a(\DFF_532.Q ),
    .b(\DFF_436.Q ),
    .y(_01226_)
  );
  al_nand2ft _05955_ (
    .a(_01225_),
    .b(_01226_),
    .y(_01227_)
  );
  al_oa21ttf _05956_ (
    .a(_01223_),
    .b(_01224_),
    .c(_01227_),
    .y(_01228_)
  );
  al_nand3fft _05957_ (
    .a(_01223_),
    .b(_01224_),
    .c(_01227_),
    .y(_01229_)
  );
  al_and3fft _05958_ (
    .a(TM0),
    .b(_01228_),
    .c(_01229_),
    .y(_01230_)
  );
  al_aoi21 _05959_ (
    .a(TM0),
    .b(\DFF_363.Q ),
    .c(TM1),
    .y(_01231_)
  );
  al_aoi21ttf _05960_ (
    .a(TM0),
    .b(\DFF_212.Q ),
    .c(TM1),
    .y(_01232_)
  );
  al_aoi21 _05961_ (
    .a(_01232_),
    .b(_00763_),
    .c(_00451_),
    .y(_01233_)
  );
  al_aoi21ftf _05962_ (
    .a(_01230_),
    .b(_01231_),
    .c(_01233_),
    .y(\DFF_244.D )
  );
  al_nor2 _05963_ (
    .a(\DFF_469.Q ),
    .b(\DFF_501.Q ),
    .y(_01234_)
  );
  al_and2 _05964_ (
    .a(\DFF_469.Q ),
    .b(\DFF_501.Q ),
    .y(_01235_)
  );
  al_and2ft _05965_ (
    .a(\DFF_437.Q ),
    .b(\DFF_533.Q ),
    .y(_01236_)
  );
  al_nand2ft _05966_ (
    .a(\DFF_533.Q ),
    .b(\DFF_437.Q ),
    .y(_01237_)
  );
  al_nand2ft _05967_ (
    .a(_01236_),
    .b(_01237_),
    .y(_01238_)
  );
  al_oa21ttf _05968_ (
    .a(_01234_),
    .b(_01235_),
    .c(_01238_),
    .y(_01239_)
  );
  al_nand3fft _05969_ (
    .a(_01234_),
    .b(_01235_),
    .c(_01238_),
    .y(_01240_)
  );
  al_and3fft _05970_ (
    .a(TM0),
    .b(_01239_),
    .c(_01240_),
    .y(_01241_)
  );
  al_aoi21 _05971_ (
    .a(TM0),
    .b(\DFF_362.Q ),
    .c(TM1),
    .y(_01242_)
  );
  al_aoi21ttf _05972_ (
    .a(TM0),
    .b(\DFF_213.Q ),
    .c(TM1),
    .y(_01243_)
  );
  al_aoi21 _05973_ (
    .a(_01243_),
    .b(_00775_),
    .c(_00451_),
    .y(_01244_)
  );
  al_aoi21ftf _05974_ (
    .a(_01241_),
    .b(_01242_),
    .c(_01244_),
    .y(\DFF_245.D )
  );
  al_nor2 _05975_ (
    .a(\DFF_470.Q ),
    .b(\DFF_502.Q ),
    .y(_01245_)
  );
  al_and2 _05976_ (
    .a(\DFF_470.Q ),
    .b(\DFF_502.Q ),
    .y(_01246_)
  );
  al_and2ft _05977_ (
    .a(\DFF_438.Q ),
    .b(\DFF_534.Q ),
    .y(_01247_)
  );
  al_nand2ft _05978_ (
    .a(\DFF_534.Q ),
    .b(\DFF_438.Q ),
    .y(_01248_)
  );
  al_nand2ft _05979_ (
    .a(_01247_),
    .b(_01248_),
    .y(_01249_)
  );
  al_oa21ttf _05980_ (
    .a(_01245_),
    .b(_01246_),
    .c(_01249_),
    .y(_01250_)
  );
  al_nand3fft _05981_ (
    .a(_01245_),
    .b(_01246_),
    .c(_01249_),
    .y(_01251_)
  );
  al_and3fft _05982_ (
    .a(TM0),
    .b(_01250_),
    .c(_01251_),
    .y(_01252_)
  );
  al_aoi21 _05983_ (
    .a(TM0),
    .b(\DFF_361.Q ),
    .c(TM1),
    .y(_01253_)
  );
  al_aoi21ttf _05984_ (
    .a(TM0),
    .b(\DFF_214.Q ),
    .c(TM1),
    .y(_01254_)
  );
  al_aoi21 _05985_ (
    .a(_01254_),
    .b(_00787_),
    .c(_00451_),
    .y(_01255_)
  );
  al_aoi21ftf _05986_ (
    .a(_01252_),
    .b(_01253_),
    .c(_01255_),
    .y(\DFF_246.D )
  );
  al_nor2 _05987_ (
    .a(\DFF_471.Q ),
    .b(\DFF_503.Q ),
    .y(_01256_)
  );
  al_and2 _05988_ (
    .a(\DFF_471.Q ),
    .b(\DFF_503.Q ),
    .y(_01257_)
  );
  al_and2ft _05989_ (
    .a(\DFF_439.Q ),
    .b(\DFF_535.Q ),
    .y(_01258_)
  );
  al_nand2ft _05990_ (
    .a(\DFF_535.Q ),
    .b(\DFF_439.Q ),
    .y(_01259_)
  );
  al_nand2ft _05991_ (
    .a(_01258_),
    .b(_01259_),
    .y(_01260_)
  );
  al_oa21ttf _05992_ (
    .a(_01256_),
    .b(_01257_),
    .c(_01260_),
    .y(_01261_)
  );
  al_nand3fft _05993_ (
    .a(_01256_),
    .b(_01257_),
    .c(_01260_),
    .y(_01262_)
  );
  al_and3fft _05994_ (
    .a(TM0),
    .b(_01261_),
    .c(_01262_),
    .y(_01263_)
  );
  al_aoi21 _05995_ (
    .a(TM0),
    .b(\DFF_360.Q ),
    .c(TM1),
    .y(_01264_)
  );
  al_aoi21ttf _05996_ (
    .a(TM0),
    .b(\DFF_215.Q ),
    .c(TM1),
    .y(_01265_)
  );
  al_aoi21 _05997_ (
    .a(_01265_),
    .b(_00799_),
    .c(_00451_),
    .y(_01266_)
  );
  al_aoi21ftf _05998_ (
    .a(_01263_),
    .b(_01264_),
    .c(_01266_),
    .y(\DFF_247.D )
  );
  al_nor2 _05999_ (
    .a(\DFF_472.Q ),
    .b(\DFF_504.Q ),
    .y(_01267_)
  );
  al_and2 _06000_ (
    .a(\DFF_472.Q ),
    .b(\DFF_504.Q ),
    .y(_01268_)
  );
  al_and2ft _06001_ (
    .a(\DFF_440.Q ),
    .b(\DFF_536.Q ),
    .y(_01269_)
  );
  al_nand2ft _06002_ (
    .a(\DFF_536.Q ),
    .b(\DFF_440.Q ),
    .y(_01270_)
  );
  al_nand2ft _06003_ (
    .a(_01269_),
    .b(_01270_),
    .y(_01271_)
  );
  al_oa21ttf _06004_ (
    .a(_01267_),
    .b(_01268_),
    .c(_01271_),
    .y(_01272_)
  );
  al_nand3fft _06005_ (
    .a(_01267_),
    .b(_01268_),
    .c(_01271_),
    .y(_01273_)
  );
  al_and3fft _06006_ (
    .a(TM0),
    .b(_01272_),
    .c(_01273_),
    .y(_01274_)
  );
  al_aoi21 _06007_ (
    .a(TM0),
    .b(\DFF_359.Q ),
    .c(TM1),
    .y(_01275_)
  );
  al_aoi21ttf _06008_ (
    .a(TM0),
    .b(\DFF_216.Q ),
    .c(TM1),
    .y(_01276_)
  );
  al_aoi21 _06009_ (
    .a(_01276_),
    .b(_00811_),
    .c(_00451_),
    .y(_01277_)
  );
  al_aoi21ftf _06010_ (
    .a(_01274_),
    .b(_01275_),
    .c(_01277_),
    .y(\DFF_248.D )
  );
  al_nor2 _06011_ (
    .a(\DFF_473.Q ),
    .b(\DFF_505.Q ),
    .y(_01278_)
  );
  al_and2 _06012_ (
    .a(\DFF_473.Q ),
    .b(\DFF_505.Q ),
    .y(_01279_)
  );
  al_and2ft _06013_ (
    .a(\DFF_441.Q ),
    .b(\DFF_537.Q ),
    .y(_01280_)
  );
  al_nand2ft _06014_ (
    .a(\DFF_537.Q ),
    .b(\DFF_441.Q ),
    .y(_01281_)
  );
  al_nand2ft _06015_ (
    .a(_01280_),
    .b(_01281_),
    .y(_01282_)
  );
  al_oa21ttf _06016_ (
    .a(_01278_),
    .b(_01279_),
    .c(_01282_),
    .y(_01283_)
  );
  al_nand3fft _06017_ (
    .a(_01278_),
    .b(_01279_),
    .c(_01282_),
    .y(_01284_)
  );
  al_and3fft _06018_ (
    .a(TM0),
    .b(_01283_),
    .c(_01284_),
    .y(_01285_)
  );
  al_aoi21 _06019_ (
    .a(TM0),
    .b(\DFF_358.Q ),
    .c(TM1),
    .y(_01286_)
  );
  al_aoi21ttf _06020_ (
    .a(TM0),
    .b(\DFF_217.Q ),
    .c(TM1),
    .y(_01287_)
  );
  al_aoi21 _06021_ (
    .a(_01287_),
    .b(_00823_),
    .c(_00451_),
    .y(_01288_)
  );
  al_aoi21ftf _06022_ (
    .a(_01285_),
    .b(_01286_),
    .c(_01288_),
    .y(\DFF_249.D )
  );
  al_nor2 _06023_ (
    .a(\DFF_474.Q ),
    .b(\DFF_506.Q ),
    .y(_01289_)
  );
  al_and2 _06024_ (
    .a(\DFF_474.Q ),
    .b(\DFF_506.Q ),
    .y(_01290_)
  );
  al_and2ft _06025_ (
    .a(\DFF_442.Q ),
    .b(\DFF_538.Q ),
    .y(_01291_)
  );
  al_nand2ft _06026_ (
    .a(\DFF_538.Q ),
    .b(\DFF_442.Q ),
    .y(_01292_)
  );
  al_nand2ft _06027_ (
    .a(_01291_),
    .b(_01292_),
    .y(_01293_)
  );
  al_oa21ttf _06028_ (
    .a(_01289_),
    .b(_01290_),
    .c(_01293_),
    .y(_01294_)
  );
  al_nand3fft _06029_ (
    .a(_01289_),
    .b(_01290_),
    .c(_01293_),
    .y(_01295_)
  );
  al_and3fft _06030_ (
    .a(TM0),
    .b(_01294_),
    .c(_01295_),
    .y(_01296_)
  );
  al_aoi21 _06031_ (
    .a(TM0),
    .b(\DFF_357.Q ),
    .c(TM1),
    .y(_01297_)
  );
  al_aoi21ttf _06032_ (
    .a(TM0),
    .b(\DFF_218.Q ),
    .c(TM1),
    .y(_01298_)
  );
  al_aoi21 _06033_ (
    .a(_01298_),
    .b(_00835_),
    .c(_00451_),
    .y(_01299_)
  );
  al_aoi21ftf _06034_ (
    .a(_01296_),
    .b(_01297_),
    .c(_01299_),
    .y(\DFF_250.D )
  );
  al_nor2 _06035_ (
    .a(\DFF_475.Q ),
    .b(\DFF_507.Q ),
    .y(_01300_)
  );
  al_and2 _06036_ (
    .a(\DFF_475.Q ),
    .b(\DFF_507.Q ),
    .y(_01301_)
  );
  al_and2ft _06037_ (
    .a(\DFF_443.Q ),
    .b(\DFF_539.Q ),
    .y(_01302_)
  );
  al_nand2ft _06038_ (
    .a(\DFF_539.Q ),
    .b(\DFF_443.Q ),
    .y(_01303_)
  );
  al_nand2ft _06039_ (
    .a(_01302_),
    .b(_01303_),
    .y(_01304_)
  );
  al_oa21ttf _06040_ (
    .a(_01300_),
    .b(_01301_),
    .c(_01304_),
    .y(_01305_)
  );
  al_nand3fft _06041_ (
    .a(_01300_),
    .b(_01301_),
    .c(_01304_),
    .y(_01306_)
  );
  al_and3fft _06042_ (
    .a(TM0),
    .b(_01305_),
    .c(_01306_),
    .y(_01307_)
  );
  al_aoi21 _06043_ (
    .a(TM0),
    .b(\DFF_356.Q ),
    .c(TM1),
    .y(_01308_)
  );
  al_aoi21ttf _06044_ (
    .a(TM0),
    .b(\DFF_219.Q ),
    .c(TM1),
    .y(_01309_)
  );
  al_aoi21 _06045_ (
    .a(_01309_),
    .b(_00847_),
    .c(_00451_),
    .y(_01310_)
  );
  al_aoi21ftf _06046_ (
    .a(_01307_),
    .b(_01308_),
    .c(_01310_),
    .y(\DFF_251.D )
  );
  al_nor2 _06047_ (
    .a(\DFF_476.Q ),
    .b(\DFF_508.Q ),
    .y(_01311_)
  );
  al_and2 _06048_ (
    .a(\DFF_476.Q ),
    .b(\DFF_508.Q ),
    .y(_01312_)
  );
  al_and2ft _06049_ (
    .a(\DFF_444.Q ),
    .b(\DFF_540.Q ),
    .y(_01313_)
  );
  al_nand2ft _06050_ (
    .a(\DFF_540.Q ),
    .b(\DFF_444.Q ),
    .y(_01314_)
  );
  al_nand2ft _06051_ (
    .a(_01313_),
    .b(_01314_),
    .y(_01315_)
  );
  al_oa21ttf _06052_ (
    .a(_01311_),
    .b(_01312_),
    .c(_01315_),
    .y(_01316_)
  );
  al_nand3fft _06053_ (
    .a(_01311_),
    .b(_01312_),
    .c(_01315_),
    .y(_01317_)
  );
  al_and3fft _06054_ (
    .a(TM0),
    .b(_01316_),
    .c(_01317_),
    .y(_01318_)
  );
  al_aoi21 _06055_ (
    .a(TM0),
    .b(\DFF_355.Q ),
    .c(TM1),
    .y(_01319_)
  );
  al_aoi21ttf _06056_ (
    .a(TM0),
    .b(\DFF_220.Q ),
    .c(TM1),
    .y(_01320_)
  );
  al_aoi21 _06057_ (
    .a(_01320_),
    .b(_00859_),
    .c(_00451_),
    .y(_01321_)
  );
  al_aoi21ftf _06058_ (
    .a(_01318_),
    .b(_01319_),
    .c(_01321_),
    .y(\DFF_252.D )
  );
  al_nor2 _06059_ (
    .a(\DFF_477.Q ),
    .b(\DFF_509.Q ),
    .y(_01322_)
  );
  al_and2 _06060_ (
    .a(\DFF_477.Q ),
    .b(\DFF_509.Q ),
    .y(_01323_)
  );
  al_and2ft _06061_ (
    .a(\DFF_445.Q ),
    .b(\DFF_541.Q ),
    .y(_01324_)
  );
  al_nand2ft _06062_ (
    .a(\DFF_541.Q ),
    .b(\DFF_445.Q ),
    .y(_01325_)
  );
  al_nand2ft _06063_ (
    .a(_01324_),
    .b(_01325_),
    .y(_01326_)
  );
  al_oa21ttf _06064_ (
    .a(_01322_),
    .b(_01323_),
    .c(_01326_),
    .y(_01327_)
  );
  al_nand3fft _06065_ (
    .a(_01322_),
    .b(_01323_),
    .c(_01326_),
    .y(_01328_)
  );
  al_and3fft _06066_ (
    .a(TM0),
    .b(_01327_),
    .c(_01328_),
    .y(_01329_)
  );
  al_aoi21 _06067_ (
    .a(TM0),
    .b(\DFF_354.Q ),
    .c(TM1),
    .y(_01330_)
  );
  al_aoi21ttf _06068_ (
    .a(TM0),
    .b(\DFF_221.Q ),
    .c(TM1),
    .y(_01331_)
  );
  al_aoi21 _06069_ (
    .a(_01331_),
    .b(_00871_),
    .c(_00451_),
    .y(_01332_)
  );
  al_aoi21ftf _06070_ (
    .a(_01329_),
    .b(_01330_),
    .c(_01332_),
    .y(\DFF_253.D )
  );
  al_nor2 _06071_ (
    .a(\DFF_478.Q ),
    .b(\DFF_510.Q ),
    .y(_01333_)
  );
  al_and2 _06072_ (
    .a(\DFF_478.Q ),
    .b(\DFF_510.Q ),
    .y(_01334_)
  );
  al_and2ft _06073_ (
    .a(\DFF_446.Q ),
    .b(\DFF_542.Q ),
    .y(_01335_)
  );
  al_nand2ft _06074_ (
    .a(\DFF_542.Q ),
    .b(\DFF_446.Q ),
    .y(_01336_)
  );
  al_nand2ft _06075_ (
    .a(_01335_),
    .b(_01336_),
    .y(_01337_)
  );
  al_oa21ttf _06076_ (
    .a(_01333_),
    .b(_01334_),
    .c(_01337_),
    .y(_01338_)
  );
  al_nand3fft _06077_ (
    .a(_01333_),
    .b(_01334_),
    .c(_01337_),
    .y(_01339_)
  );
  al_and3fft _06078_ (
    .a(TM0),
    .b(_01338_),
    .c(_01339_),
    .y(_01340_)
  );
  al_aoi21 _06079_ (
    .a(TM0),
    .b(\DFF_353.Q ),
    .c(TM1),
    .y(_01341_)
  );
  al_aoi21ttf _06080_ (
    .a(TM0),
    .b(\DFF_222.Q ),
    .c(TM1),
    .y(_01342_)
  );
  al_aoi21 _06081_ (
    .a(_01342_),
    .b(_00883_),
    .c(_00451_),
    .y(_01343_)
  );
  al_aoi21ftf _06082_ (
    .a(_01340_),
    .b(_01341_),
    .c(_01343_),
    .y(\DFF_254.D )
  );
  al_nor2 _06083_ (
    .a(\DFF_479.Q ),
    .b(\DFF_511.Q ),
    .y(_01344_)
  );
  al_and2 _06084_ (
    .a(\DFF_479.Q ),
    .b(\DFF_511.Q ),
    .y(_01345_)
  );
  al_and2ft _06085_ (
    .a(\DFF_447.Q ),
    .b(\DFF_543.Q ),
    .y(_01346_)
  );
  al_nand2ft _06086_ (
    .a(\DFF_543.Q ),
    .b(\DFF_447.Q ),
    .y(_01347_)
  );
  al_nand2ft _06087_ (
    .a(_01346_),
    .b(_01347_),
    .y(_01348_)
  );
  al_oa21ttf _06088_ (
    .a(_01344_),
    .b(_01345_),
    .c(_01348_),
    .y(_01349_)
  );
  al_nand3fft _06089_ (
    .a(_01344_),
    .b(_01345_),
    .c(_01348_),
    .y(_01350_)
  );
  al_and3fft _06090_ (
    .a(TM0),
    .b(_01349_),
    .c(_01350_),
    .y(_01351_)
  );
  al_aoi21 _06091_ (
    .a(TM0),
    .b(\DFF_352.Q ),
    .c(TM1),
    .y(_01352_)
  );
  al_aoi21ttf _06092_ (
    .a(TM0),
    .b(\DFF_223.Q ),
    .c(TM1),
    .y(_01353_)
  );
  al_aoi21 _06093_ (
    .a(_01353_),
    .b(_00895_),
    .c(_00451_),
    .y(_01354_)
  );
  al_aoi21ftf _06094_ (
    .a(_01351_),
    .b(_01352_),
    .c(_01354_),
    .y(\DFF_255.D )
  );
  al_and2 _06095_ (
    .a(RESET),
    .b(\DFF_224.Q ),
    .y(\DFF_256.D )
  );
  al_and2 _06096_ (
    .a(RESET),
    .b(\DFF_225.Q ),
    .y(\DFF_257.D )
  );
  al_and2 _06097_ (
    .a(RESET),
    .b(\DFF_226.Q ),
    .y(\DFF_258.D )
  );
  al_and2 _06098_ (
    .a(RESET),
    .b(\DFF_227.Q ),
    .y(\DFF_259.D )
  );
  al_and2 _06099_ (
    .a(RESET),
    .b(\DFF_228.Q ),
    .y(\DFF_260.D )
  );
  al_and2 _06100_ (
    .a(RESET),
    .b(\DFF_229.Q ),
    .y(\DFF_261.D )
  );
  al_and2 _06101_ (
    .a(RESET),
    .b(\DFF_230.Q ),
    .y(\DFF_262.D )
  );
  al_and2 _06102_ (
    .a(RESET),
    .b(\DFF_231.Q ),
    .y(\DFF_263.D )
  );
  al_and2 _06103_ (
    .a(RESET),
    .b(\DFF_232.Q ),
    .y(\DFF_264.D )
  );
  al_and2 _06104_ (
    .a(RESET),
    .b(\DFF_233.Q ),
    .y(\DFF_265.D )
  );
  al_and2 _06105_ (
    .a(RESET),
    .b(\DFF_234.Q ),
    .y(\DFF_266.D )
  );
  al_and2 _06106_ (
    .a(RESET),
    .b(\DFF_235.Q ),
    .y(\DFF_267.D )
  );
  al_and2 _06107_ (
    .a(RESET),
    .b(\DFF_236.Q ),
    .y(\DFF_268.D )
  );
  al_and2 _06108_ (
    .a(RESET),
    .b(\DFF_237.Q ),
    .y(\DFF_269.D )
  );
  al_and2 _06109_ (
    .a(RESET),
    .b(\DFF_238.Q ),
    .y(\DFF_270.D )
  );
  al_and2 _06110_ (
    .a(RESET),
    .b(\DFF_239.Q ),
    .y(\DFF_271.D )
  );
  al_and2 _06111_ (
    .a(RESET),
    .b(\DFF_240.Q ),
    .y(\DFF_272.D )
  );
  al_and2 _06112_ (
    .a(RESET),
    .b(\DFF_241.Q ),
    .y(\DFF_273.D )
  );
  al_and2 _06113_ (
    .a(RESET),
    .b(\DFF_242.Q ),
    .y(\DFF_274.D )
  );
  al_and2 _06114_ (
    .a(RESET),
    .b(\DFF_243.Q ),
    .y(\DFF_275.D )
  );
  al_and2 _06115_ (
    .a(RESET),
    .b(\DFF_244.Q ),
    .y(\DFF_276.D )
  );
  al_and2 _06116_ (
    .a(RESET),
    .b(\DFF_245.Q ),
    .y(\DFF_277.D )
  );
  al_and2 _06117_ (
    .a(RESET),
    .b(\DFF_246.Q ),
    .y(\DFF_278.D )
  );
  al_and2 _06118_ (
    .a(RESET),
    .b(\DFF_247.Q ),
    .y(\DFF_279.D )
  );
  al_and2 _06119_ (
    .a(RESET),
    .b(\DFF_248.Q ),
    .y(\DFF_280.D )
  );
  al_and2 _06120_ (
    .a(RESET),
    .b(\DFF_249.Q ),
    .y(\DFF_281.D )
  );
  al_and2 _06121_ (
    .a(RESET),
    .b(\DFF_250.Q ),
    .y(\DFF_282.D )
  );
  al_and2 _06122_ (
    .a(RESET),
    .b(\DFF_251.Q ),
    .y(\DFF_283.D )
  );
  al_and2 _06123_ (
    .a(RESET),
    .b(\DFF_252.Q ),
    .y(\DFF_284.D )
  );
  al_and2 _06124_ (
    .a(RESET),
    .b(\DFF_253.Q ),
    .y(\DFF_285.D )
  );
  al_and2 _06125_ (
    .a(RESET),
    .b(\DFF_254.Q ),
    .y(\DFF_286.D )
  );
  al_and2 _06126_ (
    .a(RESET),
    .b(\DFF_255.Q ),
    .y(\DFF_287.D )
  );
  al_and2 _06127_ (
    .a(RESET),
    .b(\DFF_256.Q ),
    .y(\DFF_288.D )
  );
  al_and2 _06128_ (
    .a(RESET),
    .b(\DFF_257.Q ),
    .y(\DFF_289.D )
  );
  al_and2 _06129_ (
    .a(RESET),
    .b(\DFF_258.Q ),
    .y(\DFF_290.D )
  );
  al_and2 _06130_ (
    .a(RESET),
    .b(\DFF_259.Q ),
    .y(\DFF_291.D )
  );
  al_and2 _06131_ (
    .a(RESET),
    .b(\DFF_260.Q ),
    .y(\DFF_292.D )
  );
  al_and2 _06132_ (
    .a(RESET),
    .b(\DFF_261.Q ),
    .y(\DFF_293.D )
  );
  al_and2 _06133_ (
    .a(RESET),
    .b(\DFF_262.Q ),
    .y(\DFF_294.D )
  );
  al_and2 _06134_ (
    .a(RESET),
    .b(\DFF_263.Q ),
    .y(\DFF_295.D )
  );
  al_and2 _06135_ (
    .a(RESET),
    .b(\DFF_264.Q ),
    .y(\DFF_296.D )
  );
  al_and2 _06136_ (
    .a(RESET),
    .b(\DFF_265.Q ),
    .y(\DFF_297.D )
  );
  al_and2 _06137_ (
    .a(RESET),
    .b(\DFF_266.Q ),
    .y(\DFF_298.D )
  );
  al_and2 _06138_ (
    .a(RESET),
    .b(\DFF_267.Q ),
    .y(\DFF_299.D )
  );
  al_and2 _06139_ (
    .a(RESET),
    .b(\DFF_268.Q ),
    .y(\DFF_300.D )
  );
  al_and2 _06140_ (
    .a(RESET),
    .b(\DFF_269.Q ),
    .y(\DFF_301.D )
  );
  al_and2 _06141_ (
    .a(RESET),
    .b(\DFF_270.Q ),
    .y(\DFF_302.D )
  );
  al_and2 _06142_ (
    .a(RESET),
    .b(\DFF_271.Q ),
    .y(\DFF_303.D )
  );
  al_and2 _06143_ (
    .a(RESET),
    .b(\DFF_272.Q ),
    .y(\DFF_304.D )
  );
  al_and2 _06144_ (
    .a(RESET),
    .b(\DFF_273.Q ),
    .y(\DFF_305.D )
  );
  al_and2 _06145_ (
    .a(RESET),
    .b(\DFF_274.Q ),
    .y(\DFF_306.D )
  );
  al_and2 _06146_ (
    .a(RESET),
    .b(\DFF_275.Q ),
    .y(\DFF_307.D )
  );
  al_and2 _06147_ (
    .a(RESET),
    .b(\DFF_276.Q ),
    .y(\DFF_308.D )
  );
  al_and2 _06148_ (
    .a(RESET),
    .b(\DFF_277.Q ),
    .y(\DFF_309.D )
  );
  al_and2 _06149_ (
    .a(RESET),
    .b(\DFF_278.Q ),
    .y(\DFF_310.D )
  );
  al_and2 _06150_ (
    .a(RESET),
    .b(\DFF_279.Q ),
    .y(\DFF_311.D )
  );
  al_and2 _06151_ (
    .a(RESET),
    .b(\DFF_280.Q ),
    .y(\DFF_312.D )
  );
  al_and2 _06152_ (
    .a(RESET),
    .b(\DFF_281.Q ),
    .y(\DFF_313.D )
  );
  al_and2 _06153_ (
    .a(RESET),
    .b(\DFF_282.Q ),
    .y(\DFF_314.D )
  );
  al_and2 _06154_ (
    .a(RESET),
    .b(\DFF_283.Q ),
    .y(\DFF_315.D )
  );
  al_and2 _06155_ (
    .a(RESET),
    .b(\DFF_284.Q ),
    .y(\DFF_316.D )
  );
  al_and2 _06156_ (
    .a(RESET),
    .b(\DFF_285.Q ),
    .y(\DFF_317.D )
  );
  al_and2 _06157_ (
    .a(RESET),
    .b(\DFF_286.Q ),
    .y(\DFF_318.D )
  );
  al_and2 _06158_ (
    .a(RESET),
    .b(\DFF_287.Q ),
    .y(\DFF_319.D )
  );
  al_and2 _06159_ (
    .a(RESET),
    .b(\DFF_288.Q ),
    .y(\DFF_320.D )
  );
  al_and2 _06160_ (
    .a(RESET),
    .b(\DFF_289.Q ),
    .y(\DFF_321.D )
  );
  al_and2 _06161_ (
    .a(RESET),
    .b(\DFF_290.Q ),
    .y(\DFF_322.D )
  );
  al_and2 _06162_ (
    .a(RESET),
    .b(\DFF_291.Q ),
    .y(\DFF_323.D )
  );
  al_and2 _06163_ (
    .a(RESET),
    .b(\DFF_292.Q ),
    .y(\DFF_324.D )
  );
  al_and2 _06164_ (
    .a(RESET),
    .b(\DFF_293.Q ),
    .y(\DFF_325.D )
  );
  al_and2 _06165_ (
    .a(RESET),
    .b(\DFF_294.Q ),
    .y(\DFF_326.D )
  );
  al_and2 _06166_ (
    .a(RESET),
    .b(\DFF_295.Q ),
    .y(\DFF_327.D )
  );
  al_and2 _06167_ (
    .a(RESET),
    .b(\DFF_296.Q ),
    .y(\DFF_328.D )
  );
  al_and2 _06168_ (
    .a(RESET),
    .b(\DFF_297.Q ),
    .y(\DFF_329.D )
  );
  al_and2 _06169_ (
    .a(RESET),
    .b(\DFF_298.Q ),
    .y(\DFF_330.D )
  );
  al_and2 _06170_ (
    .a(RESET),
    .b(\DFF_299.Q ),
    .y(\DFF_331.D )
  );
  al_and2 _06171_ (
    .a(RESET),
    .b(\DFF_300.Q ),
    .y(\DFF_332.D )
  );
  al_and2 _06172_ (
    .a(RESET),
    .b(\DFF_301.Q ),
    .y(\DFF_333.D )
  );
  al_and2 _06173_ (
    .a(RESET),
    .b(\DFF_302.Q ),
    .y(\DFF_334.D )
  );
  al_and2 _06174_ (
    .a(RESET),
    .b(\DFF_303.Q ),
    .y(\DFF_335.D )
  );
  al_and2 _06175_ (
    .a(RESET),
    .b(\DFF_304.Q ),
    .y(\DFF_336.D )
  );
  al_and2 _06176_ (
    .a(RESET),
    .b(\DFF_305.Q ),
    .y(\DFF_337.D )
  );
  al_and2 _06177_ (
    .a(RESET),
    .b(\DFF_306.Q ),
    .y(\DFF_338.D )
  );
  al_and2 _06178_ (
    .a(RESET),
    .b(\DFF_307.Q ),
    .y(\DFF_339.D )
  );
  al_and2 _06179_ (
    .a(RESET),
    .b(\DFF_308.Q ),
    .y(\DFF_340.D )
  );
  al_and2 _06180_ (
    .a(RESET),
    .b(\DFF_309.Q ),
    .y(\DFF_341.D )
  );
  al_and2 _06181_ (
    .a(RESET),
    .b(\DFF_310.Q ),
    .y(\DFF_342.D )
  );
  al_and2 _06182_ (
    .a(RESET),
    .b(\DFF_311.Q ),
    .y(\DFF_343.D )
  );
  al_and2 _06183_ (
    .a(RESET),
    .b(\DFF_312.Q ),
    .y(\DFF_344.D )
  );
  al_and2 _06184_ (
    .a(RESET),
    .b(\DFF_313.Q ),
    .y(\DFF_345.D )
  );
  al_and2 _06185_ (
    .a(RESET),
    .b(\DFF_314.Q ),
    .y(\DFF_346.D )
  );
  al_and2 _06186_ (
    .a(RESET),
    .b(\DFF_315.Q ),
    .y(\DFF_347.D )
  );
  al_and2 _06187_ (
    .a(RESET),
    .b(\DFF_316.Q ),
    .y(\DFF_348.D )
  );
  al_and2 _06188_ (
    .a(RESET),
    .b(\DFF_317.Q ),
    .y(\DFF_349.D )
  );
  al_and2 _06189_ (
    .a(RESET),
    .b(\DFF_318.Q ),
    .y(\DFF_350.D )
  );
  al_and2 _06190_ (
    .a(RESET),
    .b(\DFF_319.Q ),
    .y(\DFF_351.D )
  );
  al_oa21ftt _06191_ (
    .a(\DFF_351.Q ),
    .b(\DFF_383.Q ),
    .c(RESET),
    .y(_01355_)
  );
  al_aoi21ftf _06192_ (
    .a(\DFF_351.Q ),
    .b(\DFF_383.Q ),
    .c(_01355_),
    .y(\DFF_352.D )
  );
  al_oa21ftt _06193_ (
    .a(\DFF_350.Q ),
    .b(\DFF_352.Q ),
    .c(RESET),
    .y(_01356_)
  );
  al_aoi21ftf _06194_ (
    .a(\DFF_350.Q ),
    .b(\DFF_352.Q ),
    .c(_01356_),
    .y(\DFF_353.D )
  );
  al_oa21ftt _06195_ (
    .a(\DFF_349.Q ),
    .b(\DFF_353.Q ),
    .c(RESET),
    .y(_01357_)
  );
  al_aoi21ftf _06196_ (
    .a(\DFF_349.Q ),
    .b(\DFF_353.Q ),
    .c(_01357_),
    .y(\DFF_354.D )
  );
  al_oa21ftt _06197_ (
    .a(\DFF_348.Q ),
    .b(\DFF_354.Q ),
    .c(RESET),
    .y(_01358_)
  );
  al_aoi21ftf _06198_ (
    .a(\DFF_348.Q ),
    .b(\DFF_354.Q ),
    .c(_01358_),
    .y(\DFF_355.D )
  );
  al_nand2ft _06199_ (
    .a(\DFF_347.Q ),
    .b(\DFF_355.Q ),
    .y(_01359_)
  );
  al_nand2ft _06200_ (
    .a(\DFF_355.Q ),
    .b(\DFF_347.Q ),
    .y(_01360_)
  );
  al_ao21ttf _06201_ (
    .a(_01359_),
    .b(_01360_),
    .c(\DFF_383.Q ),
    .y(_01361_)
  );
  al_nand3ftt _06202_ (
    .a(\DFF_383.Q ),
    .b(_01359_),
    .c(_01360_),
    .y(_01362_)
  );
  al_aoi21 _06203_ (
    .a(_01362_),
    .b(_01361_),
    .c(_00451_),
    .y(\DFF_356.D )
  );
  al_oa21ftt _06204_ (
    .a(\DFF_346.Q ),
    .b(\DFF_356.Q ),
    .c(RESET),
    .y(_01363_)
  );
  al_aoi21ftf _06205_ (
    .a(\DFF_346.Q ),
    .b(\DFF_356.Q ),
    .c(_01363_),
    .y(\DFF_357.D )
  );
  al_oa21ftt _06206_ (
    .a(\DFF_345.Q ),
    .b(\DFF_357.Q ),
    .c(RESET),
    .y(_01364_)
  );
  al_aoi21ftf _06207_ (
    .a(\DFF_345.Q ),
    .b(\DFF_357.Q ),
    .c(_01364_),
    .y(\DFF_358.D )
  );
  al_oa21ftt _06208_ (
    .a(\DFF_344.Q ),
    .b(\DFF_358.Q ),
    .c(RESET),
    .y(_01365_)
  );
  al_aoi21ftf _06209_ (
    .a(\DFF_344.Q ),
    .b(\DFF_358.Q ),
    .c(_01365_),
    .y(\DFF_359.D )
  );
  al_oa21ftt _06210_ (
    .a(\DFF_343.Q ),
    .b(\DFF_359.Q ),
    .c(RESET),
    .y(_01366_)
  );
  al_aoi21ftf _06211_ (
    .a(\DFF_343.Q ),
    .b(\DFF_359.Q ),
    .c(_01366_),
    .y(\DFF_360.D )
  );
  al_oa21ftt _06212_ (
    .a(\DFF_342.Q ),
    .b(\DFF_360.Q ),
    .c(RESET),
    .y(_01367_)
  );
  al_aoi21ftf _06213_ (
    .a(\DFF_342.Q ),
    .b(\DFF_360.Q ),
    .c(_01367_),
    .y(\DFF_361.D )
  );
  al_oa21ftt _06214_ (
    .a(\DFF_341.Q ),
    .b(\DFF_361.Q ),
    .c(RESET),
    .y(_01368_)
  );
  al_aoi21ftf _06215_ (
    .a(\DFF_341.Q ),
    .b(\DFF_361.Q ),
    .c(_01368_),
    .y(\DFF_362.D )
  );
  al_nand2ft _06216_ (
    .a(\DFF_340.Q ),
    .b(\DFF_362.Q ),
    .y(_01369_)
  );
  al_nand2ft _06217_ (
    .a(\DFF_362.Q ),
    .b(\DFF_340.Q ),
    .y(_01370_)
  );
  al_ao21ttf _06218_ (
    .a(_01369_),
    .b(_01370_),
    .c(\DFF_383.Q ),
    .y(_01371_)
  );
  al_nand3ftt _06219_ (
    .a(\DFF_383.Q ),
    .b(_01369_),
    .c(_01370_),
    .y(_01372_)
  );
  al_aoi21 _06220_ (
    .a(_01372_),
    .b(_01371_),
    .c(_00451_),
    .y(\DFF_363.D )
  );
  al_oa21ftt _06221_ (
    .a(\DFF_339.Q ),
    .b(\DFF_363.Q ),
    .c(RESET),
    .y(_01373_)
  );
  al_aoi21ftf _06222_ (
    .a(\DFF_339.Q ),
    .b(\DFF_363.Q ),
    .c(_01373_),
    .y(\DFF_364.D )
  );
  al_oa21ftt _06223_ (
    .a(\DFF_338.Q ),
    .b(\DFF_364.Q ),
    .c(RESET),
    .y(_01374_)
  );
  al_aoi21ftf _06224_ (
    .a(\DFF_338.Q ),
    .b(\DFF_364.Q ),
    .c(_01374_),
    .y(\DFF_365.D )
  );
  al_oa21ftt _06225_ (
    .a(\DFF_337.Q ),
    .b(\DFF_365.Q ),
    .c(RESET),
    .y(_01375_)
  );
  al_aoi21ftf _06226_ (
    .a(\DFF_337.Q ),
    .b(\DFF_365.Q ),
    .c(_01375_),
    .y(\DFF_366.D )
  );
  al_oa21ftt _06227_ (
    .a(\DFF_336.Q ),
    .b(\DFF_366.Q ),
    .c(RESET),
    .y(_01376_)
  );
  al_aoi21ftf _06228_ (
    .a(\DFF_336.Q ),
    .b(\DFF_366.Q ),
    .c(_01376_),
    .y(\DFF_367.D )
  );
  al_nand2ft _06229_ (
    .a(\DFF_335.Q ),
    .b(\DFF_367.Q ),
    .y(_01377_)
  );
  al_nand2ft _06230_ (
    .a(\DFF_367.Q ),
    .b(\DFF_335.Q ),
    .y(_01378_)
  );
  al_ao21ttf _06231_ (
    .a(_01377_),
    .b(_01378_),
    .c(\DFF_383.Q ),
    .y(_01379_)
  );
  al_nand3ftt _06232_ (
    .a(\DFF_383.Q ),
    .b(_01377_),
    .c(_01378_),
    .y(_01380_)
  );
  al_aoi21 _06233_ (
    .a(_01380_),
    .b(_01379_),
    .c(_00451_),
    .y(\DFF_368.D )
  );
  al_oa21ftt _06234_ (
    .a(\DFF_334.Q ),
    .b(\DFF_368.Q ),
    .c(RESET),
    .y(_01381_)
  );
  al_aoi21ftf _06235_ (
    .a(\DFF_334.Q ),
    .b(\DFF_368.Q ),
    .c(_01381_),
    .y(\DFF_369.D )
  );
  al_oa21ftt _06236_ (
    .a(\DFF_333.Q ),
    .b(\DFF_369.Q ),
    .c(RESET),
    .y(_01382_)
  );
  al_aoi21ftf _06237_ (
    .a(\DFF_333.Q ),
    .b(\DFF_369.Q ),
    .c(_01382_),
    .y(\DFF_370.D )
  );
  al_oa21ftt _06238_ (
    .a(\DFF_332.Q ),
    .b(\DFF_370.Q ),
    .c(RESET),
    .y(_01383_)
  );
  al_aoi21ftf _06239_ (
    .a(\DFF_332.Q ),
    .b(\DFF_370.Q ),
    .c(_01383_),
    .y(\DFF_371.D )
  );
  al_oa21ftt _06240_ (
    .a(\DFF_331.Q ),
    .b(\DFF_371.Q ),
    .c(RESET),
    .y(_01384_)
  );
  al_aoi21ftf _06241_ (
    .a(\DFF_331.Q ),
    .b(\DFF_371.Q ),
    .c(_01384_),
    .y(\DFF_372.D )
  );
  al_oa21ftt _06242_ (
    .a(\DFF_330.Q ),
    .b(\DFF_372.Q ),
    .c(RESET),
    .y(_01385_)
  );
  al_aoi21ftf _06243_ (
    .a(\DFF_330.Q ),
    .b(\DFF_372.Q ),
    .c(_01385_),
    .y(\DFF_373.D )
  );
  al_oa21ftt _06244_ (
    .a(\DFF_329.Q ),
    .b(\DFF_373.Q ),
    .c(RESET),
    .y(_01386_)
  );
  al_aoi21ftf _06245_ (
    .a(\DFF_329.Q ),
    .b(\DFF_373.Q ),
    .c(_01386_),
    .y(\DFF_374.D )
  );
  al_oa21ftt _06246_ (
    .a(\DFF_328.Q ),
    .b(\DFF_374.Q ),
    .c(RESET),
    .y(_01387_)
  );
  al_aoi21ftf _06247_ (
    .a(\DFF_328.Q ),
    .b(\DFF_374.Q ),
    .c(_01387_),
    .y(\DFF_375.D )
  );
  al_oa21ftt _06248_ (
    .a(\DFF_327.Q ),
    .b(\DFF_375.Q ),
    .c(RESET),
    .y(_01388_)
  );
  al_aoi21ftf _06249_ (
    .a(\DFF_327.Q ),
    .b(\DFF_375.Q ),
    .c(_01388_),
    .y(\DFF_376.D )
  );
  al_oa21ftt _06250_ (
    .a(\DFF_326.Q ),
    .b(\DFF_376.Q ),
    .c(RESET),
    .y(_01389_)
  );
  al_aoi21ftf _06251_ (
    .a(\DFF_326.Q ),
    .b(\DFF_376.Q ),
    .c(_01389_),
    .y(\DFF_377.D )
  );
  al_oa21ftt _06252_ (
    .a(\DFF_325.Q ),
    .b(\DFF_377.Q ),
    .c(RESET),
    .y(_01390_)
  );
  al_aoi21ftf _06253_ (
    .a(\DFF_325.Q ),
    .b(\DFF_377.Q ),
    .c(_01390_),
    .y(\DFF_378.D )
  );
  al_oa21ftt _06254_ (
    .a(\DFF_324.Q ),
    .b(\DFF_378.Q ),
    .c(RESET),
    .y(_01391_)
  );
  al_aoi21ftf _06255_ (
    .a(\DFF_324.Q ),
    .b(\DFF_378.Q ),
    .c(_01391_),
    .y(\DFF_379.D )
  );
  al_oa21ftt _06256_ (
    .a(\DFF_323.Q ),
    .b(\DFF_379.Q ),
    .c(RESET),
    .y(_01392_)
  );
  al_aoi21ftf _06257_ (
    .a(\DFF_323.Q ),
    .b(\DFF_379.Q ),
    .c(_01392_),
    .y(\DFF_380.D )
  );
  al_oa21ftt _06258_ (
    .a(\DFF_322.Q ),
    .b(\DFF_380.Q ),
    .c(RESET),
    .y(_01393_)
  );
  al_aoi21ftf _06259_ (
    .a(\DFF_322.Q ),
    .b(\DFF_380.Q ),
    .c(_01393_),
    .y(\DFF_381.D )
  );
  al_oa21ftt _06260_ (
    .a(\DFF_321.Q ),
    .b(\DFF_381.Q ),
    .c(RESET),
    .y(_01394_)
  );
  al_aoi21ftf _06261_ (
    .a(\DFF_321.Q ),
    .b(\DFF_381.Q ),
    .c(_01394_),
    .y(\DFF_382.D )
  );
  al_oa21ftt _06262_ (
    .a(\DFF_320.Q ),
    .b(\DFF_382.Q ),
    .c(RESET),
    .y(_01395_)
  );
  al_aoi21ftf _06263_ (
    .a(\DFF_320.Q ),
    .b(\DFF_382.Q ),
    .c(_01395_),
    .y(\DFF_383.D )
  );
  al_and2 _06264_ (
    .a(RESET),
    .b(\DFF_385.Q ),
    .y(\DFF_384.D )
  );
  al_and2 _06265_ (
    .a(RESET),
    .b(\DFF_386.Q ),
    .y(\DFF_385.D )
  );
  al_and2 _06266_ (
    .a(RESET),
    .b(\DFF_387.Q ),
    .y(\DFF_386.D )
  );
  al_and2 _06267_ (
    .a(RESET),
    .b(\DFF_388.Q ),
    .y(\DFF_387.D )
  );
  al_and2 _06268_ (
    .a(RESET),
    .b(\DFF_389.Q ),
    .y(\DFF_388.D )
  );
  al_and2 _06269_ (
    .a(RESET),
    .b(\DFF_390.Q ),
    .y(\DFF_389.D )
  );
  al_and2 _06270_ (
    .a(RESET),
    .b(\DFF_391.Q ),
    .y(\DFF_390.D )
  );
  al_and2 _06271_ (
    .a(RESET),
    .b(\DFF_392.Q ),
    .y(\DFF_391.D )
  );
  al_and2 _06272_ (
    .a(RESET),
    .b(\DFF_393.Q ),
    .y(\DFF_392.D )
  );
  al_and2 _06273_ (
    .a(RESET),
    .b(\DFF_394.Q ),
    .y(\DFF_393.D )
  );
  al_and2 _06274_ (
    .a(RESET),
    .b(\DFF_395.Q ),
    .y(\DFF_394.D )
  );
  al_and2 _06275_ (
    .a(RESET),
    .b(\DFF_396.Q ),
    .y(\DFF_395.D )
  );
  al_and2 _06276_ (
    .a(RESET),
    .b(\DFF_397.Q ),
    .y(\DFF_396.D )
  );
  al_and2 _06277_ (
    .a(RESET),
    .b(\DFF_398.Q ),
    .y(\DFF_397.D )
  );
  al_and2 _06278_ (
    .a(RESET),
    .b(\DFF_399.Q ),
    .y(\DFF_398.D )
  );
  al_and2 _06279_ (
    .a(RESET),
    .b(\DFF_400.Q ),
    .y(\DFF_399.D )
  );
  al_and2 _06280_ (
    .a(RESET),
    .b(\DFF_401.Q ),
    .y(\DFF_400.D )
  );
  al_and2 _06281_ (
    .a(RESET),
    .b(\DFF_402.Q ),
    .y(\DFF_401.D )
  );
  al_and2 _06282_ (
    .a(RESET),
    .b(\DFF_403.Q ),
    .y(\DFF_402.D )
  );
  al_and2 _06283_ (
    .a(RESET),
    .b(\DFF_404.Q ),
    .y(\DFF_403.D )
  );
  al_and2 _06284_ (
    .a(RESET),
    .b(\DFF_405.Q ),
    .y(\DFF_404.D )
  );
  al_and2 _06285_ (
    .a(RESET),
    .b(\DFF_406.Q ),
    .y(\DFF_405.D )
  );
  al_and2 _06286_ (
    .a(RESET),
    .b(\DFF_407.Q ),
    .y(\DFF_406.D )
  );
  al_and2 _06287_ (
    .a(RESET),
    .b(\DFF_408.Q ),
    .y(\DFF_407.D )
  );
  al_and2 _06288_ (
    .a(RESET),
    .b(\DFF_409.Q ),
    .y(\DFF_408.D )
  );
  al_and2 _06289_ (
    .a(RESET),
    .b(\DFF_410.Q ),
    .y(\DFF_409.D )
  );
  al_and2 _06290_ (
    .a(RESET),
    .b(\DFF_411.Q ),
    .y(\DFF_410.D )
  );
  al_and2 _06291_ (
    .a(RESET),
    .b(\DFF_412.Q ),
    .y(\DFF_411.D )
  );
  al_and2 _06292_ (
    .a(RESET),
    .b(\DFF_413.Q ),
    .y(\DFF_412.D )
  );
  al_and2 _06293_ (
    .a(RESET),
    .b(\DFF_414.Q ),
    .y(\DFF_413.D )
  );
  al_and2 _06294_ (
    .a(RESET),
    .b(\DFF_415.Q ),
    .y(\DFF_414.D )
  );
  al_and2ft _06295_ (
    .a(\DFF_384.Q ),
    .b(RESET),
    .y(\DFF_415.D )
  );
  al_or2 _06296_ (
    .a(TM1),
    .b(\DFF_672.Q ),
    .y(_01396_)
  );
  al_nand2 _06297_ (
    .a(TM1),
    .b(\DFF_672.Q ),
    .y(_01397_)
  );
  al_nand3 _06298_ (
    .a(\DFF_704.Q ),
    .b(_01396_),
    .c(_01397_),
    .y(_01398_)
  );
  al_nand2ft _06299_ (
    .a(TM1),
    .b(\DFF_672.Q ),
    .y(_01399_)
  );
  al_and2ft _06300_ (
    .a(\DFF_672.Q ),
    .b(TM1),
    .y(_01400_)
  );
  al_and3fft _06301_ (
    .a(\DFF_704.Q ),
    .b(_01400_),
    .c(_01399_),
    .y(_01401_)
  );
  al_and2ft _06302_ (
    .a(\DFF_640.Q ),
    .b(\DFF_608.Q ),
    .y(_01402_)
  );
  al_nand2ft _06303_ (
    .a(\DFF_608.Q ),
    .b(\DFF_640.Q ),
    .y(_01403_)
  );
  al_nand2ft _06304_ (
    .a(_01402_),
    .b(_01403_),
    .y(_01404_)
  );
  al_oai21ftf _06305_ (
    .a(_01398_),
    .b(_01401_),
    .c(_01404_),
    .y(_01405_)
  );
  al_nand3ftt _06306_ (
    .a(_01401_),
    .b(_01398_),
    .c(_01404_),
    .y(_01406_)
  );
  al_nand3 _06307_ (
    .a(_00448_),
    .b(_01405_),
    .c(_01406_),
    .y(_01407_)
  );
  al_aoi21 _06308_ (
    .a(TM0),
    .b(\DFF_575.Q ),
    .c(TM1),
    .y(_01408_)
  );
  al_nand2 _06309_ (
    .a(_01408_),
    .b(_01407_),
    .y(_01409_)
  );
  al_aoi21ttf _06310_ (
    .a(\DFF_384.Q ),
    .b(TM0),
    .c(TM1),
    .y(_01410_)
  );
  al_and2 _06311_ (
    .a(_01410_),
    .b(_00950_),
    .y(_01411_)
  );
  al_nor3fft _06312_ (
    .a(RESET),
    .b(_01409_),
    .c(_01411_),
    .y(\DFF_416.D )
  );
  al_or2 _06313_ (
    .a(TM1),
    .b(\DFF_673.Q ),
    .y(_01412_)
  );
  al_nand2 _06314_ (
    .a(TM1),
    .b(\DFF_673.Q ),
    .y(_01413_)
  );
  al_nand3 _06315_ (
    .a(\DFF_705.Q ),
    .b(_01412_),
    .c(_01413_),
    .y(_01414_)
  );
  al_nand2ft _06316_ (
    .a(TM1),
    .b(\DFF_673.Q ),
    .y(_01415_)
  );
  al_and2ft _06317_ (
    .a(\DFF_673.Q ),
    .b(TM1),
    .y(_01416_)
  );
  al_and3fft _06318_ (
    .a(\DFF_705.Q ),
    .b(_01416_),
    .c(_01415_),
    .y(_01417_)
  );
  al_and2ft _06319_ (
    .a(\DFF_641.Q ),
    .b(\DFF_609.Q ),
    .y(_01418_)
  );
  al_nand2ft _06320_ (
    .a(\DFF_609.Q ),
    .b(\DFF_641.Q ),
    .y(_01419_)
  );
  al_nand2ft _06321_ (
    .a(_01418_),
    .b(_01419_),
    .y(_01420_)
  );
  al_oai21ftf _06322_ (
    .a(_01414_),
    .b(_01417_),
    .c(_01420_),
    .y(_01421_)
  );
  al_nand3ftt _06323_ (
    .a(_01417_),
    .b(_01414_),
    .c(_01420_),
    .y(_01422_)
  );
  al_nand3 _06324_ (
    .a(_00448_),
    .b(_01421_),
    .c(_01422_),
    .y(_01423_)
  );
  al_aoi21 _06325_ (
    .a(TM0),
    .b(\DFF_574.Q ),
    .c(TM1),
    .y(_01424_)
  );
  al_nand2 _06326_ (
    .a(_01424_),
    .b(_01423_),
    .y(_01425_)
  );
  al_aoi21ttf _06327_ (
    .a(TM0),
    .b(\DFF_385.Q ),
    .c(TM1),
    .y(_01426_)
  );
  al_and2 _06328_ (
    .a(_01426_),
    .b(_00965_),
    .y(_01427_)
  );
  al_nor3fft _06329_ (
    .a(RESET),
    .b(_01425_),
    .c(_01427_),
    .y(\DFF_417.D )
  );
  al_or2 _06330_ (
    .a(TM1),
    .b(\DFF_674.Q ),
    .y(_01428_)
  );
  al_nand2 _06331_ (
    .a(TM1),
    .b(\DFF_674.Q ),
    .y(_01429_)
  );
  al_nand3 _06332_ (
    .a(\DFF_706.Q ),
    .b(_01428_),
    .c(_01429_),
    .y(_01430_)
  );
  al_nand2ft _06333_ (
    .a(TM1),
    .b(\DFF_674.Q ),
    .y(_01431_)
  );
  al_and2ft _06334_ (
    .a(\DFF_674.Q ),
    .b(TM1),
    .y(_01432_)
  );
  al_and3fft _06335_ (
    .a(\DFF_706.Q ),
    .b(_01432_),
    .c(_01431_),
    .y(_01433_)
  );
  al_and2ft _06336_ (
    .a(\DFF_642.Q ),
    .b(\DFF_610.Q ),
    .y(_01434_)
  );
  al_nand2ft _06337_ (
    .a(\DFF_610.Q ),
    .b(\DFF_642.Q ),
    .y(_01435_)
  );
  al_nand2ft _06338_ (
    .a(_01434_),
    .b(_01435_),
    .y(_01436_)
  );
  al_oai21ftf _06339_ (
    .a(_01430_),
    .b(_01433_),
    .c(_01436_),
    .y(_01437_)
  );
  al_nand3ftt _06340_ (
    .a(_01433_),
    .b(_01430_),
    .c(_01436_),
    .y(_01438_)
  );
  al_nand3 _06341_ (
    .a(_00448_),
    .b(_01437_),
    .c(_01438_),
    .y(_01439_)
  );
  al_aoi21 _06342_ (
    .a(TM0),
    .b(\DFF_573.Q ),
    .c(TM1),
    .y(_01440_)
  );
  al_nand2 _06343_ (
    .a(_01440_),
    .b(_01439_),
    .y(_01441_)
  );
  al_aoi21ttf _06344_ (
    .a(TM0),
    .b(\DFF_386.Q ),
    .c(TM1),
    .y(_01442_)
  );
  al_and2 _06345_ (
    .a(_01442_),
    .b(_00980_),
    .y(_01443_)
  );
  al_nor3fft _06346_ (
    .a(RESET),
    .b(_01441_),
    .c(_01443_),
    .y(\DFF_418.D )
  );
  al_or2 _06347_ (
    .a(TM1),
    .b(\DFF_675.Q ),
    .y(_01444_)
  );
  al_nand2 _06348_ (
    .a(TM1),
    .b(\DFF_675.Q ),
    .y(_01445_)
  );
  al_nand3 _06349_ (
    .a(\DFF_707.Q ),
    .b(_01444_),
    .c(_01445_),
    .y(_01446_)
  );
  al_nand2ft _06350_ (
    .a(TM1),
    .b(\DFF_675.Q ),
    .y(_01447_)
  );
  al_and2ft _06351_ (
    .a(\DFF_675.Q ),
    .b(TM1),
    .y(_01448_)
  );
  al_and3fft _06352_ (
    .a(\DFF_707.Q ),
    .b(_01448_),
    .c(_01447_),
    .y(_01449_)
  );
  al_and2ft _06353_ (
    .a(\DFF_643.Q ),
    .b(\DFF_611.Q ),
    .y(_01450_)
  );
  al_nand2ft _06354_ (
    .a(\DFF_611.Q ),
    .b(\DFF_643.Q ),
    .y(_01451_)
  );
  al_nand2ft _06355_ (
    .a(_01450_),
    .b(_01451_),
    .y(_01452_)
  );
  al_oai21ftf _06356_ (
    .a(_01446_),
    .b(_01449_),
    .c(_01452_),
    .y(_01453_)
  );
  al_nand3ftt _06357_ (
    .a(_01449_),
    .b(_01446_),
    .c(_01452_),
    .y(_01454_)
  );
  al_nand3 _06358_ (
    .a(_00448_),
    .b(_01453_),
    .c(_01454_),
    .y(_01455_)
  );
  al_aoi21 _06359_ (
    .a(TM0),
    .b(\DFF_572.Q ),
    .c(TM1),
    .y(_01456_)
  );
  al_nand2 _06360_ (
    .a(_01456_),
    .b(_01455_),
    .y(_01457_)
  );
  al_aoi21ttf _06361_ (
    .a(TM0),
    .b(\DFF_387.Q ),
    .c(TM1),
    .y(_01458_)
  );
  al_and2 _06362_ (
    .a(_01458_),
    .b(_00995_),
    .y(_01459_)
  );
  al_nor3fft _06363_ (
    .a(RESET),
    .b(_01457_),
    .c(_01459_),
    .y(\DFF_419.D )
  );
  al_or2 _06364_ (
    .a(TM1),
    .b(\DFF_676.Q ),
    .y(_01460_)
  );
  al_nand2 _06365_ (
    .a(TM1),
    .b(\DFF_676.Q ),
    .y(_01461_)
  );
  al_nand3 _06366_ (
    .a(\DFF_708.Q ),
    .b(_01460_),
    .c(_01461_),
    .y(_01462_)
  );
  al_nand2ft _06367_ (
    .a(TM1),
    .b(\DFF_676.Q ),
    .y(_01463_)
  );
  al_and2ft _06368_ (
    .a(\DFF_676.Q ),
    .b(TM1),
    .y(_01464_)
  );
  al_and3fft _06369_ (
    .a(\DFF_708.Q ),
    .b(_01464_),
    .c(_01463_),
    .y(_01465_)
  );
  al_and2ft _06370_ (
    .a(\DFF_644.Q ),
    .b(\DFF_612.Q ),
    .y(_01466_)
  );
  al_nand2ft _06371_ (
    .a(\DFF_612.Q ),
    .b(\DFF_644.Q ),
    .y(_01467_)
  );
  al_nand2ft _06372_ (
    .a(_01466_),
    .b(_01467_),
    .y(_01468_)
  );
  al_oai21ftf _06373_ (
    .a(_01462_),
    .b(_01465_),
    .c(_01468_),
    .y(_01469_)
  );
  al_nand3ftt _06374_ (
    .a(_01465_),
    .b(_01462_),
    .c(_01468_),
    .y(_01470_)
  );
  al_nand3 _06375_ (
    .a(_00448_),
    .b(_01469_),
    .c(_01470_),
    .y(_01471_)
  );
  al_aoi21 _06376_ (
    .a(TM0),
    .b(\DFF_571.Q ),
    .c(TM1),
    .y(_01472_)
  );
  al_nand2 _06377_ (
    .a(_01472_),
    .b(_01471_),
    .y(_01473_)
  );
  al_aoi21ttf _06378_ (
    .a(TM0),
    .b(\DFF_388.Q ),
    .c(TM1),
    .y(_01474_)
  );
  al_and2 _06379_ (
    .a(_01474_),
    .b(_01010_),
    .y(_01475_)
  );
  al_nor3fft _06380_ (
    .a(RESET),
    .b(_01473_),
    .c(_01475_),
    .y(\DFF_420.D )
  );
  al_or2 _06381_ (
    .a(TM1),
    .b(\DFF_677.Q ),
    .y(_01476_)
  );
  al_nand2 _06382_ (
    .a(TM1),
    .b(\DFF_677.Q ),
    .y(_01477_)
  );
  al_nand3 _06383_ (
    .a(\DFF_709.Q ),
    .b(_01476_),
    .c(_01477_),
    .y(_01478_)
  );
  al_nand2ft _06384_ (
    .a(TM1),
    .b(\DFF_677.Q ),
    .y(_01479_)
  );
  al_and2ft _06385_ (
    .a(\DFF_677.Q ),
    .b(TM1),
    .y(_01480_)
  );
  al_and3fft _06386_ (
    .a(\DFF_709.Q ),
    .b(_01480_),
    .c(_01479_),
    .y(_01481_)
  );
  al_and2ft _06387_ (
    .a(\DFF_645.Q ),
    .b(\DFF_613.Q ),
    .y(_01482_)
  );
  al_nand2ft _06388_ (
    .a(\DFF_613.Q ),
    .b(\DFF_645.Q ),
    .y(_01483_)
  );
  al_nand2ft _06389_ (
    .a(_01482_),
    .b(_01483_),
    .y(_01484_)
  );
  al_oai21ftf _06390_ (
    .a(_01478_),
    .b(_01481_),
    .c(_01484_),
    .y(_01485_)
  );
  al_nand3ftt _06391_ (
    .a(_01481_),
    .b(_01478_),
    .c(_01484_),
    .y(_01486_)
  );
  al_nand3 _06392_ (
    .a(_00448_),
    .b(_01485_),
    .c(_01486_),
    .y(_01487_)
  );
  al_aoi21 _06393_ (
    .a(TM0),
    .b(\DFF_570.Q ),
    .c(TM1),
    .y(_01488_)
  );
  al_nand2 _06394_ (
    .a(_01488_),
    .b(_01487_),
    .y(_01489_)
  );
  al_aoi21ttf _06395_ (
    .a(TM0),
    .b(\DFF_389.Q ),
    .c(TM1),
    .y(_01490_)
  );
  al_and2 _06396_ (
    .a(_01490_),
    .b(_01025_),
    .y(_01491_)
  );
  al_nor3fft _06397_ (
    .a(RESET),
    .b(_01489_),
    .c(_01491_),
    .y(\DFF_421.D )
  );
  al_or2 _06398_ (
    .a(TM1),
    .b(\DFF_678.Q ),
    .y(_01492_)
  );
  al_nand2 _06399_ (
    .a(TM1),
    .b(\DFF_678.Q ),
    .y(_01493_)
  );
  al_nand3 _06400_ (
    .a(\DFF_710.Q ),
    .b(_01492_),
    .c(_01493_),
    .y(_01494_)
  );
  al_nand2ft _06401_ (
    .a(TM1),
    .b(\DFF_678.Q ),
    .y(_01495_)
  );
  al_and2ft _06402_ (
    .a(\DFF_678.Q ),
    .b(TM1),
    .y(_01496_)
  );
  al_and3fft _06403_ (
    .a(\DFF_710.Q ),
    .b(_01496_),
    .c(_01495_),
    .y(_01497_)
  );
  al_and2ft _06404_ (
    .a(\DFF_646.Q ),
    .b(\DFF_614.Q ),
    .y(_01498_)
  );
  al_nand2ft _06405_ (
    .a(\DFF_614.Q ),
    .b(\DFF_646.Q ),
    .y(_01499_)
  );
  al_nand2ft _06406_ (
    .a(_01498_),
    .b(_01499_),
    .y(_01500_)
  );
  al_oai21ftf _06407_ (
    .a(_01494_),
    .b(_01497_),
    .c(_01500_),
    .y(_01501_)
  );
  al_nand3ftt _06408_ (
    .a(_01497_),
    .b(_01494_),
    .c(_01500_),
    .y(_01502_)
  );
  al_nand3 _06409_ (
    .a(_00448_),
    .b(_01501_),
    .c(_01502_),
    .y(_01503_)
  );
  al_aoi21 _06410_ (
    .a(TM0),
    .b(\DFF_569.Q ),
    .c(TM1),
    .y(_01504_)
  );
  al_nand2 _06411_ (
    .a(_01504_),
    .b(_01503_),
    .y(_01505_)
  );
  al_aoi21ttf _06412_ (
    .a(TM0),
    .b(\DFF_390.Q ),
    .c(TM1),
    .y(_01506_)
  );
  al_and2 _06413_ (
    .a(_01506_),
    .b(_01040_),
    .y(_01507_)
  );
  al_nor3fft _06414_ (
    .a(RESET),
    .b(_01505_),
    .c(_01507_),
    .y(\DFF_422.D )
  );
  al_or2 _06415_ (
    .a(TM1),
    .b(\DFF_679.Q ),
    .y(_01508_)
  );
  al_nand2 _06416_ (
    .a(TM1),
    .b(\DFF_679.Q ),
    .y(_01509_)
  );
  al_nand3 _06417_ (
    .a(\DFF_711.Q ),
    .b(_01508_),
    .c(_01509_),
    .y(_01510_)
  );
  al_nand2ft _06418_ (
    .a(TM1),
    .b(\DFF_679.Q ),
    .y(_01511_)
  );
  al_and2ft _06419_ (
    .a(\DFF_679.Q ),
    .b(TM1),
    .y(_01512_)
  );
  al_and3fft _06420_ (
    .a(\DFF_711.Q ),
    .b(_01512_),
    .c(_01511_),
    .y(_01513_)
  );
  al_and2ft _06421_ (
    .a(\DFF_647.Q ),
    .b(\DFF_615.Q ),
    .y(_01514_)
  );
  al_nand2ft _06422_ (
    .a(\DFF_615.Q ),
    .b(\DFF_647.Q ),
    .y(_01515_)
  );
  al_nand2ft _06423_ (
    .a(_01514_),
    .b(_01515_),
    .y(_01516_)
  );
  al_oai21ftf _06424_ (
    .a(_01510_),
    .b(_01513_),
    .c(_01516_),
    .y(_01517_)
  );
  al_nand3ftt _06425_ (
    .a(_01513_),
    .b(_01510_),
    .c(_01516_),
    .y(_01518_)
  );
  al_nand3 _06426_ (
    .a(_00448_),
    .b(_01517_),
    .c(_01518_),
    .y(_01519_)
  );
  al_aoi21 _06427_ (
    .a(TM0),
    .b(\DFF_568.Q ),
    .c(TM1),
    .y(_01520_)
  );
  al_nand2 _06428_ (
    .a(_01520_),
    .b(_01519_),
    .y(_01521_)
  );
  al_aoi21ttf _06429_ (
    .a(TM0),
    .b(\DFF_391.Q ),
    .c(TM1),
    .y(_01522_)
  );
  al_and2 _06430_ (
    .a(_01522_),
    .b(_01055_),
    .y(_01523_)
  );
  al_nor3fft _06431_ (
    .a(RESET),
    .b(_01521_),
    .c(_01523_),
    .y(\DFF_423.D )
  );
  al_or2 _06432_ (
    .a(TM1),
    .b(\DFF_680.Q ),
    .y(_01524_)
  );
  al_nand2 _06433_ (
    .a(TM1),
    .b(\DFF_680.Q ),
    .y(_01525_)
  );
  al_nand3 _06434_ (
    .a(\DFF_712.Q ),
    .b(_01524_),
    .c(_01525_),
    .y(_01526_)
  );
  al_nand2ft _06435_ (
    .a(TM1),
    .b(\DFF_680.Q ),
    .y(_01527_)
  );
  al_and2ft _06436_ (
    .a(\DFF_680.Q ),
    .b(TM1),
    .y(_01528_)
  );
  al_and3fft _06437_ (
    .a(\DFF_712.Q ),
    .b(_01528_),
    .c(_01527_),
    .y(_01529_)
  );
  al_and2ft _06438_ (
    .a(\DFF_648.Q ),
    .b(\DFF_616.Q ),
    .y(_01530_)
  );
  al_nand2ft _06439_ (
    .a(\DFF_616.Q ),
    .b(\DFF_648.Q ),
    .y(_01531_)
  );
  al_nand2ft _06440_ (
    .a(_01530_),
    .b(_01531_),
    .y(_01532_)
  );
  al_oai21ftf _06441_ (
    .a(_01526_),
    .b(_01529_),
    .c(_01532_),
    .y(_01533_)
  );
  al_nand3ftt _06442_ (
    .a(_01529_),
    .b(_01526_),
    .c(_01532_),
    .y(_01534_)
  );
  al_nand3 _06443_ (
    .a(_00448_),
    .b(_01533_),
    .c(_01534_),
    .y(_01535_)
  );
  al_aoi21 _06444_ (
    .a(TM0),
    .b(\DFF_567.Q ),
    .c(TM1),
    .y(_01536_)
  );
  al_nand2 _06445_ (
    .a(_01536_),
    .b(_01535_),
    .y(_01537_)
  );
  al_aoi21ttf _06446_ (
    .a(TM0),
    .b(\DFF_392.Q ),
    .c(TM1),
    .y(_01538_)
  );
  al_and2 _06447_ (
    .a(_01538_),
    .b(_01070_),
    .y(_01539_)
  );
  al_nor3fft _06448_ (
    .a(RESET),
    .b(_01537_),
    .c(_01539_),
    .y(\DFF_424.D )
  );
  al_or2 _06449_ (
    .a(TM1),
    .b(\DFF_681.Q ),
    .y(_01540_)
  );
  al_nand2 _06450_ (
    .a(TM1),
    .b(\DFF_681.Q ),
    .y(_01541_)
  );
  al_nand3 _06451_ (
    .a(\DFF_713.Q ),
    .b(_01540_),
    .c(_01541_),
    .y(_01542_)
  );
  al_nand2ft _06452_ (
    .a(TM1),
    .b(\DFF_681.Q ),
    .y(_01543_)
  );
  al_and2ft _06453_ (
    .a(\DFF_681.Q ),
    .b(TM1),
    .y(_01544_)
  );
  al_and3fft _06454_ (
    .a(\DFF_713.Q ),
    .b(_01544_),
    .c(_01543_),
    .y(_01545_)
  );
  al_and2ft _06455_ (
    .a(\DFF_649.Q ),
    .b(\DFF_617.Q ),
    .y(_01546_)
  );
  al_nand2ft _06456_ (
    .a(\DFF_617.Q ),
    .b(\DFF_649.Q ),
    .y(_01547_)
  );
  al_nand2ft _06457_ (
    .a(_01546_),
    .b(_01547_),
    .y(_01548_)
  );
  al_oai21ftf _06458_ (
    .a(_01542_),
    .b(_01545_),
    .c(_01548_),
    .y(_01549_)
  );
  al_nand3ftt _06459_ (
    .a(_01545_),
    .b(_01542_),
    .c(_01548_),
    .y(_01550_)
  );
  al_nand3 _06460_ (
    .a(_00448_),
    .b(_01549_),
    .c(_01550_),
    .y(_01551_)
  );
  al_aoi21 _06461_ (
    .a(TM0),
    .b(\DFF_566.Q ),
    .c(TM1),
    .y(_01552_)
  );
  al_nand2 _06462_ (
    .a(_01552_),
    .b(_01551_),
    .y(_01553_)
  );
  al_aoi21ttf _06463_ (
    .a(TM0),
    .b(\DFF_393.Q ),
    .c(TM1),
    .y(_01554_)
  );
  al_and2 _06464_ (
    .a(_01554_),
    .b(_01085_),
    .y(_01555_)
  );
  al_nor3fft _06465_ (
    .a(RESET),
    .b(_01553_),
    .c(_01555_),
    .y(\DFF_425.D )
  );
  al_or2 _06466_ (
    .a(TM1),
    .b(\DFF_682.Q ),
    .y(_01556_)
  );
  al_nand2 _06467_ (
    .a(TM1),
    .b(\DFF_682.Q ),
    .y(_01557_)
  );
  al_nand3 _06468_ (
    .a(\DFF_714.Q ),
    .b(_01556_),
    .c(_01557_),
    .y(_01558_)
  );
  al_nand2ft _06469_ (
    .a(TM1),
    .b(\DFF_682.Q ),
    .y(_01559_)
  );
  al_and2ft _06470_ (
    .a(\DFF_682.Q ),
    .b(TM1),
    .y(_01560_)
  );
  al_and3fft _06471_ (
    .a(\DFF_714.Q ),
    .b(_01560_),
    .c(_01559_),
    .y(_01561_)
  );
  al_and2ft _06472_ (
    .a(\DFF_650.Q ),
    .b(\DFF_618.Q ),
    .y(_01562_)
  );
  al_nand2ft _06473_ (
    .a(\DFF_618.Q ),
    .b(\DFF_650.Q ),
    .y(_01563_)
  );
  al_nand2ft _06474_ (
    .a(_01562_),
    .b(_01563_),
    .y(_01564_)
  );
  al_oai21ftf _06475_ (
    .a(_01558_),
    .b(_01561_),
    .c(_01564_),
    .y(_01565_)
  );
  al_nand3ftt _06476_ (
    .a(_01561_),
    .b(_01558_),
    .c(_01564_),
    .y(_01566_)
  );
  al_nand3 _06477_ (
    .a(_00448_),
    .b(_01565_),
    .c(_01566_),
    .y(_01567_)
  );
  al_aoi21 _06478_ (
    .a(TM0),
    .b(\DFF_565.Q ),
    .c(TM1),
    .y(_01568_)
  );
  al_nand2 _06479_ (
    .a(_01568_),
    .b(_01567_),
    .y(_01569_)
  );
  al_aoi21ttf _06480_ (
    .a(TM0),
    .b(\DFF_394.Q ),
    .c(TM1),
    .y(_01570_)
  );
  al_and2 _06481_ (
    .a(_01570_),
    .b(_01100_),
    .y(_01571_)
  );
  al_nor3fft _06482_ (
    .a(RESET),
    .b(_01569_),
    .c(_01571_),
    .y(\DFF_426.D )
  );
  al_or2 _06483_ (
    .a(TM1),
    .b(\DFF_683.Q ),
    .y(_01572_)
  );
  al_nand2 _06484_ (
    .a(TM1),
    .b(\DFF_683.Q ),
    .y(_01573_)
  );
  al_nand3 _06485_ (
    .a(\DFF_715.Q ),
    .b(_01572_),
    .c(_01573_),
    .y(_01574_)
  );
  al_nand2ft _06486_ (
    .a(TM1),
    .b(\DFF_683.Q ),
    .y(_01575_)
  );
  al_and2ft _06487_ (
    .a(\DFF_683.Q ),
    .b(TM1),
    .y(_01576_)
  );
  al_and3fft _06488_ (
    .a(\DFF_715.Q ),
    .b(_01576_),
    .c(_01575_),
    .y(_01577_)
  );
  al_and2ft _06489_ (
    .a(\DFF_651.Q ),
    .b(\DFF_619.Q ),
    .y(_01578_)
  );
  al_nand2ft _06490_ (
    .a(\DFF_619.Q ),
    .b(\DFF_651.Q ),
    .y(_01579_)
  );
  al_nand2ft _06491_ (
    .a(_01578_),
    .b(_01579_),
    .y(_01580_)
  );
  al_oai21ftf _06492_ (
    .a(_01574_),
    .b(_01577_),
    .c(_01580_),
    .y(_01581_)
  );
  al_nand3ftt _06493_ (
    .a(_01577_),
    .b(_01574_),
    .c(_01580_),
    .y(_01582_)
  );
  al_nand3 _06494_ (
    .a(_00448_),
    .b(_01581_),
    .c(_01582_),
    .y(_01583_)
  );
  al_aoi21 _06495_ (
    .a(TM0),
    .b(\DFF_564.Q ),
    .c(TM1),
    .y(_01584_)
  );
  al_nand2 _06496_ (
    .a(_01584_),
    .b(_01583_),
    .y(_01585_)
  );
  al_aoi21ttf _06497_ (
    .a(TM0),
    .b(\DFF_395.Q ),
    .c(TM1),
    .y(_01586_)
  );
  al_and2 _06498_ (
    .a(_01586_),
    .b(_01115_),
    .y(_01587_)
  );
  al_nor3fft _06499_ (
    .a(RESET),
    .b(_01585_),
    .c(_01587_),
    .y(\DFF_427.D )
  );
  al_or2 _06500_ (
    .a(TM1),
    .b(\DFF_684.Q ),
    .y(_01588_)
  );
  al_nand2 _06501_ (
    .a(TM1),
    .b(\DFF_684.Q ),
    .y(_01589_)
  );
  al_nand3 _06502_ (
    .a(\DFF_716.Q ),
    .b(_01588_),
    .c(_01589_),
    .y(_01590_)
  );
  al_nand2ft _06503_ (
    .a(TM1),
    .b(\DFF_684.Q ),
    .y(_01591_)
  );
  al_and2ft _06504_ (
    .a(\DFF_684.Q ),
    .b(TM1),
    .y(_01592_)
  );
  al_and3fft _06505_ (
    .a(\DFF_716.Q ),
    .b(_01592_),
    .c(_01591_),
    .y(_01593_)
  );
  al_and2ft _06506_ (
    .a(\DFF_652.Q ),
    .b(\DFF_620.Q ),
    .y(_01594_)
  );
  al_nand2ft _06507_ (
    .a(\DFF_620.Q ),
    .b(\DFF_652.Q ),
    .y(_01595_)
  );
  al_nand2ft _06508_ (
    .a(_01594_),
    .b(_01595_),
    .y(_01596_)
  );
  al_oai21ftf _06509_ (
    .a(_01590_),
    .b(_01593_),
    .c(_01596_),
    .y(_01597_)
  );
  al_nand3ftt _06510_ (
    .a(_01593_),
    .b(_01590_),
    .c(_01596_),
    .y(_01598_)
  );
  al_nand3 _06511_ (
    .a(_00448_),
    .b(_01597_),
    .c(_01598_),
    .y(_01599_)
  );
  al_aoi21 _06512_ (
    .a(TM0),
    .b(\DFF_563.Q ),
    .c(TM1),
    .y(_01600_)
  );
  al_nand2 _06513_ (
    .a(_01600_),
    .b(_01599_),
    .y(_01601_)
  );
  al_aoi21ttf _06514_ (
    .a(TM0),
    .b(\DFF_396.Q ),
    .c(TM1),
    .y(_01602_)
  );
  al_and2 _06515_ (
    .a(_01602_),
    .b(_01130_),
    .y(_01603_)
  );
  al_nor3fft _06516_ (
    .a(RESET),
    .b(_01601_),
    .c(_01603_),
    .y(\DFF_428.D )
  );
  al_or2 _06517_ (
    .a(TM1),
    .b(\DFF_685.Q ),
    .y(_01604_)
  );
  al_nand2 _06518_ (
    .a(TM1),
    .b(\DFF_685.Q ),
    .y(_01605_)
  );
  al_nand3 _06519_ (
    .a(\DFF_717.Q ),
    .b(_01604_),
    .c(_01605_),
    .y(_01606_)
  );
  al_nand2ft _06520_ (
    .a(TM1),
    .b(\DFF_685.Q ),
    .y(_01607_)
  );
  al_and2ft _06521_ (
    .a(\DFF_685.Q ),
    .b(TM1),
    .y(_01608_)
  );
  al_and3fft _06522_ (
    .a(\DFF_717.Q ),
    .b(_01608_),
    .c(_01607_),
    .y(_01609_)
  );
  al_and2ft _06523_ (
    .a(\DFF_653.Q ),
    .b(\DFF_621.Q ),
    .y(_01610_)
  );
  al_nand2ft _06524_ (
    .a(\DFF_621.Q ),
    .b(\DFF_653.Q ),
    .y(_01611_)
  );
  al_nand2ft _06525_ (
    .a(_01610_),
    .b(_01611_),
    .y(_01612_)
  );
  al_oai21ftf _06526_ (
    .a(_01606_),
    .b(_01609_),
    .c(_01612_),
    .y(_01613_)
  );
  al_nand3ftt _06527_ (
    .a(_01609_),
    .b(_01606_),
    .c(_01612_),
    .y(_01614_)
  );
  al_nand3 _06528_ (
    .a(_00448_),
    .b(_01613_),
    .c(_01614_),
    .y(_01615_)
  );
  al_aoi21 _06529_ (
    .a(TM0),
    .b(\DFF_562.Q ),
    .c(TM1),
    .y(_01616_)
  );
  al_nand2 _06530_ (
    .a(_01616_),
    .b(_01615_),
    .y(_01617_)
  );
  al_aoi21ttf _06531_ (
    .a(TM0),
    .b(\DFF_397.Q ),
    .c(TM1),
    .y(_01618_)
  );
  al_and2 _06532_ (
    .a(_01618_),
    .b(_01145_),
    .y(_01619_)
  );
  al_nor3fft _06533_ (
    .a(RESET),
    .b(_01617_),
    .c(_01619_),
    .y(\DFF_429.D )
  );
  al_or2 _06534_ (
    .a(TM1),
    .b(\DFF_686.Q ),
    .y(_01620_)
  );
  al_nand2 _06535_ (
    .a(TM1),
    .b(\DFF_686.Q ),
    .y(_01621_)
  );
  al_nand3 _06536_ (
    .a(\DFF_718.Q ),
    .b(_01620_),
    .c(_01621_),
    .y(_01622_)
  );
  al_nand2ft _06537_ (
    .a(TM1),
    .b(\DFF_686.Q ),
    .y(_01623_)
  );
  al_and2ft _06538_ (
    .a(\DFF_686.Q ),
    .b(TM1),
    .y(_01624_)
  );
  al_and3fft _06539_ (
    .a(\DFF_718.Q ),
    .b(_01624_),
    .c(_01623_),
    .y(_01625_)
  );
  al_and2ft _06540_ (
    .a(\DFF_654.Q ),
    .b(\DFF_622.Q ),
    .y(_01626_)
  );
  al_nand2ft _06541_ (
    .a(\DFF_622.Q ),
    .b(\DFF_654.Q ),
    .y(_01627_)
  );
  al_nand2ft _06542_ (
    .a(_01626_),
    .b(_01627_),
    .y(_01628_)
  );
  al_oai21ftf _06543_ (
    .a(_01622_),
    .b(_01625_),
    .c(_01628_),
    .y(_01629_)
  );
  al_nand3ftt _06544_ (
    .a(_01625_),
    .b(_01622_),
    .c(_01628_),
    .y(_01630_)
  );
  al_nand3 _06545_ (
    .a(_00448_),
    .b(_01629_),
    .c(_01630_),
    .y(_01631_)
  );
  al_aoi21 _06546_ (
    .a(TM0),
    .b(\DFF_561.Q ),
    .c(TM1),
    .y(_01632_)
  );
  al_nand2 _06547_ (
    .a(_01632_),
    .b(_01631_),
    .y(_01633_)
  );
  al_aoi21ttf _06548_ (
    .a(TM0),
    .b(\DFF_398.Q ),
    .c(TM1),
    .y(_01634_)
  );
  al_and2 _06549_ (
    .a(_01634_),
    .b(_01160_),
    .y(_01635_)
  );
  al_nor3fft _06550_ (
    .a(RESET),
    .b(_01633_),
    .c(_01635_),
    .y(\DFF_430.D )
  );
  al_or2 _06551_ (
    .a(TM1),
    .b(\DFF_687.Q ),
    .y(_01636_)
  );
  al_nand2 _06552_ (
    .a(TM1),
    .b(\DFF_687.Q ),
    .y(_01637_)
  );
  al_nand3 _06553_ (
    .a(\DFF_719.Q ),
    .b(_01636_),
    .c(_01637_),
    .y(_01638_)
  );
  al_nand2ft _06554_ (
    .a(TM1),
    .b(\DFF_687.Q ),
    .y(_01639_)
  );
  al_and2ft _06555_ (
    .a(\DFF_687.Q ),
    .b(TM1),
    .y(_01640_)
  );
  al_and3fft _06556_ (
    .a(\DFF_719.Q ),
    .b(_01640_),
    .c(_01639_),
    .y(_01641_)
  );
  al_and2ft _06557_ (
    .a(\DFF_655.Q ),
    .b(\DFF_623.Q ),
    .y(_01642_)
  );
  al_nand2ft _06558_ (
    .a(\DFF_623.Q ),
    .b(\DFF_655.Q ),
    .y(_01643_)
  );
  al_nand2ft _06559_ (
    .a(_01642_),
    .b(_01643_),
    .y(_01644_)
  );
  al_oai21ftf _06560_ (
    .a(_01638_),
    .b(_01641_),
    .c(_01644_),
    .y(_01645_)
  );
  al_nand3ftt _06561_ (
    .a(_01641_),
    .b(_01638_),
    .c(_01644_),
    .y(_01646_)
  );
  al_nand3 _06562_ (
    .a(_00448_),
    .b(_01645_),
    .c(_01646_),
    .y(_01647_)
  );
  al_aoi21 _06563_ (
    .a(TM0),
    .b(\DFF_560.Q ),
    .c(TM1),
    .y(_01648_)
  );
  al_nand2 _06564_ (
    .a(_01648_),
    .b(_01647_),
    .y(_01649_)
  );
  al_aoi21ttf _06565_ (
    .a(TM0),
    .b(\DFF_399.Q ),
    .c(TM1),
    .y(_01650_)
  );
  al_and2 _06566_ (
    .a(_01650_),
    .b(_01175_),
    .y(_01651_)
  );
  al_nor3fft _06567_ (
    .a(RESET),
    .b(_01649_),
    .c(_01651_),
    .y(\DFF_431.D )
  );
  al_inv _06568_ (
    .a(TM1),
    .y(_01652_)
  );
  al_nor2 _06569_ (
    .a(\DFF_656.Q ),
    .b(\DFF_688.Q ),
    .y(_01653_)
  );
  al_and2 _06570_ (
    .a(\DFF_656.Q ),
    .b(\DFF_688.Q ),
    .y(_01654_)
  );
  al_and2ft _06571_ (
    .a(\DFF_624.Q ),
    .b(\DFF_720.Q ),
    .y(_01655_)
  );
  al_nand2ft _06572_ (
    .a(\DFF_720.Q ),
    .b(\DFF_624.Q ),
    .y(_01656_)
  );
  al_nand2ft _06573_ (
    .a(_01655_),
    .b(_01656_),
    .y(_01657_)
  );
  al_oa21ttf _06574_ (
    .a(_01653_),
    .b(_01654_),
    .c(_01657_),
    .y(_01658_)
  );
  al_nand3fft _06575_ (
    .a(_01653_),
    .b(_01654_),
    .c(_01657_),
    .y(_01659_)
  );
  al_and3fft _06576_ (
    .a(TM0),
    .b(_01658_),
    .c(_01659_),
    .y(_01660_)
  );
  al_nand2 _06577_ (
    .a(TM0),
    .b(\DFF_559.Q ),
    .y(_01661_)
  );
  al_or3fft _06578_ (
    .a(_01652_),
    .b(_01661_),
    .c(_01660_),
    .y(_01662_)
  );
  al_and2 _06579_ (
    .a(TM0),
    .b(\DFF_400.Q ),
    .y(_01663_)
  );
  al_and3fft _06580_ (
    .a(_01663_),
    .b(_01186_),
    .c(TM1),
    .y(_01664_)
  );
  al_nor3fft _06581_ (
    .a(RESET),
    .b(_01662_),
    .c(_01664_),
    .y(\DFF_432.D )
  );
  al_nor2 _06582_ (
    .a(\DFF_657.Q ),
    .b(\DFF_689.Q ),
    .y(_01665_)
  );
  al_and2 _06583_ (
    .a(\DFF_657.Q ),
    .b(\DFF_689.Q ),
    .y(_01666_)
  );
  al_and2ft _06584_ (
    .a(\DFF_625.Q ),
    .b(\DFF_721.Q ),
    .y(_01667_)
  );
  al_nand2ft _06585_ (
    .a(\DFF_721.Q ),
    .b(\DFF_625.Q ),
    .y(_01668_)
  );
  al_nand2ft _06586_ (
    .a(_01667_),
    .b(_01668_),
    .y(_01669_)
  );
  al_oa21ttf _06587_ (
    .a(_01665_),
    .b(_01666_),
    .c(_01669_),
    .y(_01670_)
  );
  al_nand3fft _06588_ (
    .a(_01665_),
    .b(_01666_),
    .c(_01669_),
    .y(_01671_)
  );
  al_and3fft _06589_ (
    .a(TM0),
    .b(_01670_),
    .c(_01671_),
    .y(_01672_)
  );
  al_nand2 _06590_ (
    .a(TM0),
    .b(\DFF_558.Q ),
    .y(_01673_)
  );
  al_or3fft _06591_ (
    .a(_01652_),
    .b(_01673_),
    .c(_01672_),
    .y(_01674_)
  );
  al_and2 _06592_ (
    .a(TM0),
    .b(\DFF_401.Q ),
    .y(_01675_)
  );
  al_and3fft _06593_ (
    .a(_01675_),
    .b(_01197_),
    .c(TM1),
    .y(_01676_)
  );
  al_nor3fft _06594_ (
    .a(RESET),
    .b(_01674_),
    .c(_01676_),
    .y(\DFF_433.D )
  );
  al_nor2 _06595_ (
    .a(\DFF_658.Q ),
    .b(\DFF_690.Q ),
    .y(_01677_)
  );
  al_and2 _06596_ (
    .a(\DFF_658.Q ),
    .b(\DFF_690.Q ),
    .y(_01678_)
  );
  al_and2ft _06597_ (
    .a(\DFF_626.Q ),
    .b(\DFF_722.Q ),
    .y(_01679_)
  );
  al_nand2ft _06598_ (
    .a(\DFF_722.Q ),
    .b(\DFF_626.Q ),
    .y(_01680_)
  );
  al_nand2ft _06599_ (
    .a(_01679_),
    .b(_01680_),
    .y(_01681_)
  );
  al_oa21ttf _06600_ (
    .a(_01677_),
    .b(_01678_),
    .c(_01681_),
    .y(_01682_)
  );
  al_nand3fft _06601_ (
    .a(_01677_),
    .b(_01678_),
    .c(_01681_),
    .y(_01683_)
  );
  al_and3fft _06602_ (
    .a(TM0),
    .b(_01682_),
    .c(_01683_),
    .y(_01684_)
  );
  al_nand2 _06603_ (
    .a(TM0),
    .b(\DFF_557.Q ),
    .y(_01685_)
  );
  al_or3fft _06604_ (
    .a(_01652_),
    .b(_01685_),
    .c(_01684_),
    .y(_01686_)
  );
  al_and2 _06605_ (
    .a(TM0),
    .b(\DFF_402.Q ),
    .y(_01687_)
  );
  al_and3fft _06606_ (
    .a(_01687_),
    .b(_01208_),
    .c(TM1),
    .y(_01688_)
  );
  al_nor3fft _06607_ (
    .a(RESET),
    .b(_01686_),
    .c(_01688_),
    .y(\DFF_434.D )
  );
  al_nor2 _06608_ (
    .a(\DFF_659.Q ),
    .b(\DFF_691.Q ),
    .y(_01689_)
  );
  al_and2 _06609_ (
    .a(\DFF_659.Q ),
    .b(\DFF_691.Q ),
    .y(_01690_)
  );
  al_and2ft _06610_ (
    .a(\DFF_627.Q ),
    .b(\DFF_723.Q ),
    .y(_01691_)
  );
  al_nand2ft _06611_ (
    .a(\DFF_723.Q ),
    .b(\DFF_627.Q ),
    .y(_01692_)
  );
  al_nand2ft _06612_ (
    .a(_01691_),
    .b(_01692_),
    .y(_01693_)
  );
  al_oa21ttf _06613_ (
    .a(_01689_),
    .b(_01690_),
    .c(_01693_),
    .y(_01694_)
  );
  al_nand3fft _06614_ (
    .a(_01689_),
    .b(_01690_),
    .c(_01693_),
    .y(_01695_)
  );
  al_and3fft _06615_ (
    .a(TM0),
    .b(_01694_),
    .c(_01695_),
    .y(_01696_)
  );
  al_nand2 _06616_ (
    .a(TM0),
    .b(\DFF_556.Q ),
    .y(_01697_)
  );
  al_or3fft _06617_ (
    .a(_01652_),
    .b(_01697_),
    .c(_01696_),
    .y(_01698_)
  );
  al_and2 _06618_ (
    .a(TM0),
    .b(\DFF_403.Q ),
    .y(_01699_)
  );
  al_and3fft _06619_ (
    .a(_01699_),
    .b(_01219_),
    .c(TM1),
    .y(_01700_)
  );
  al_nor3fft _06620_ (
    .a(RESET),
    .b(_01698_),
    .c(_01700_),
    .y(\DFF_435.D )
  );
  al_nor2 _06621_ (
    .a(\DFF_660.Q ),
    .b(\DFF_692.Q ),
    .y(_01701_)
  );
  al_and2 _06622_ (
    .a(\DFF_660.Q ),
    .b(\DFF_692.Q ),
    .y(_01702_)
  );
  al_and2ft _06623_ (
    .a(\DFF_628.Q ),
    .b(\DFF_724.Q ),
    .y(_01703_)
  );
  al_nand2ft _06624_ (
    .a(\DFF_724.Q ),
    .b(\DFF_628.Q ),
    .y(_01704_)
  );
  al_nand2ft _06625_ (
    .a(_01703_),
    .b(_01704_),
    .y(_01705_)
  );
  al_oa21ttf _06626_ (
    .a(_01701_),
    .b(_01702_),
    .c(_01705_),
    .y(_01706_)
  );
  al_nand3fft _06627_ (
    .a(_01701_),
    .b(_01702_),
    .c(_01705_),
    .y(_01707_)
  );
  al_and3fft _06628_ (
    .a(TM0),
    .b(_01706_),
    .c(_01707_),
    .y(_01708_)
  );
  al_nand2 _06629_ (
    .a(TM0),
    .b(\DFF_555.Q ),
    .y(_01709_)
  );
  al_or3fft _06630_ (
    .a(_01652_),
    .b(_01709_),
    .c(_01708_),
    .y(_01710_)
  );
  al_and2 _06631_ (
    .a(TM0),
    .b(\DFF_404.Q ),
    .y(_01711_)
  );
  al_and3fft _06632_ (
    .a(_01711_),
    .b(_01230_),
    .c(TM1),
    .y(_01712_)
  );
  al_nor3fft _06633_ (
    .a(RESET),
    .b(_01710_),
    .c(_01712_),
    .y(\DFF_436.D )
  );
  al_nor2 _06634_ (
    .a(\DFF_661.Q ),
    .b(\DFF_693.Q ),
    .y(_01713_)
  );
  al_and2 _06635_ (
    .a(\DFF_661.Q ),
    .b(\DFF_693.Q ),
    .y(_01714_)
  );
  al_and2ft _06636_ (
    .a(\DFF_629.Q ),
    .b(\DFF_725.Q ),
    .y(_01715_)
  );
  al_nand2ft _06637_ (
    .a(\DFF_725.Q ),
    .b(\DFF_629.Q ),
    .y(_01716_)
  );
  al_nand2ft _06638_ (
    .a(_01715_),
    .b(_01716_),
    .y(_01717_)
  );
  al_oa21ttf _06639_ (
    .a(_01713_),
    .b(_01714_),
    .c(_01717_),
    .y(_01718_)
  );
  al_nand3fft _06640_ (
    .a(_01713_),
    .b(_01714_),
    .c(_01717_),
    .y(_01719_)
  );
  al_and3fft _06641_ (
    .a(TM0),
    .b(_01718_),
    .c(_01719_),
    .y(_01720_)
  );
  al_nand2 _06642_ (
    .a(TM0),
    .b(\DFF_554.Q ),
    .y(_01721_)
  );
  al_or3fft _06643_ (
    .a(_01652_),
    .b(_01721_),
    .c(_01720_),
    .y(_01722_)
  );
  al_and2 _06644_ (
    .a(TM0),
    .b(\DFF_405.Q ),
    .y(_01723_)
  );
  al_and3fft _06645_ (
    .a(_01723_),
    .b(_01241_),
    .c(TM1),
    .y(_01724_)
  );
  al_nor3fft _06646_ (
    .a(RESET),
    .b(_01722_),
    .c(_01724_),
    .y(\DFF_437.D )
  );
  al_nor2 _06647_ (
    .a(\DFF_662.Q ),
    .b(\DFF_694.Q ),
    .y(_01725_)
  );
  al_and2 _06648_ (
    .a(\DFF_662.Q ),
    .b(\DFF_694.Q ),
    .y(_01726_)
  );
  al_and2ft _06649_ (
    .a(\DFF_630.Q ),
    .b(\DFF_726.Q ),
    .y(_01727_)
  );
  al_nand2ft _06650_ (
    .a(\DFF_726.Q ),
    .b(\DFF_630.Q ),
    .y(_01728_)
  );
  al_nand2ft _06651_ (
    .a(_01727_),
    .b(_01728_),
    .y(_01729_)
  );
  al_oa21ttf _06652_ (
    .a(_01725_),
    .b(_01726_),
    .c(_01729_),
    .y(_01730_)
  );
  al_nand3fft _06653_ (
    .a(_01725_),
    .b(_01726_),
    .c(_01729_),
    .y(_01731_)
  );
  al_and3fft _06654_ (
    .a(TM0),
    .b(_01730_),
    .c(_01731_),
    .y(_01732_)
  );
  al_nand2 _06655_ (
    .a(TM0),
    .b(\DFF_553.Q ),
    .y(_01733_)
  );
  al_or3fft _06656_ (
    .a(_01652_),
    .b(_01733_),
    .c(_01732_),
    .y(_01734_)
  );
  al_and2 _06657_ (
    .a(TM0),
    .b(\DFF_406.Q ),
    .y(_01735_)
  );
  al_and3fft _06658_ (
    .a(_01735_),
    .b(_01252_),
    .c(TM1),
    .y(_01736_)
  );
  al_nor3fft _06659_ (
    .a(RESET),
    .b(_01734_),
    .c(_01736_),
    .y(\DFF_438.D )
  );
  al_nor2 _06660_ (
    .a(\DFF_663.Q ),
    .b(\DFF_695.Q ),
    .y(_01737_)
  );
  al_and2 _06661_ (
    .a(\DFF_663.Q ),
    .b(\DFF_695.Q ),
    .y(_01738_)
  );
  al_and2ft _06662_ (
    .a(\DFF_631.Q ),
    .b(\DFF_727.Q ),
    .y(_01739_)
  );
  al_nand2ft _06663_ (
    .a(\DFF_727.Q ),
    .b(\DFF_631.Q ),
    .y(_01740_)
  );
  al_nand2ft _06664_ (
    .a(_01739_),
    .b(_01740_),
    .y(_01741_)
  );
  al_oa21ttf _06665_ (
    .a(_01737_),
    .b(_01738_),
    .c(_01741_),
    .y(_01742_)
  );
  al_nand3fft _06666_ (
    .a(_01737_),
    .b(_01738_),
    .c(_01741_),
    .y(_01743_)
  );
  al_and3fft _06667_ (
    .a(TM0),
    .b(_01742_),
    .c(_01743_),
    .y(_01744_)
  );
  al_nand2 _06668_ (
    .a(TM0),
    .b(\DFF_552.Q ),
    .y(_01745_)
  );
  al_or3fft _06669_ (
    .a(_01652_),
    .b(_01745_),
    .c(_01744_),
    .y(_01746_)
  );
  al_and2 _06670_ (
    .a(TM0),
    .b(\DFF_407.Q ),
    .y(_01747_)
  );
  al_and3fft _06671_ (
    .a(_01747_),
    .b(_01263_),
    .c(TM1),
    .y(_01748_)
  );
  al_nor3fft _06672_ (
    .a(RESET),
    .b(_01746_),
    .c(_01748_),
    .y(\DFF_439.D )
  );
  al_nor2 _06673_ (
    .a(\DFF_664.Q ),
    .b(\DFF_696.Q ),
    .y(_01749_)
  );
  al_and2 _06674_ (
    .a(\DFF_664.Q ),
    .b(\DFF_696.Q ),
    .y(_01750_)
  );
  al_and2ft _06675_ (
    .a(\DFF_632.Q ),
    .b(\DFF_728.Q ),
    .y(_01751_)
  );
  al_nand2ft _06676_ (
    .a(\DFF_728.Q ),
    .b(\DFF_632.Q ),
    .y(_01752_)
  );
  al_nand2ft _06677_ (
    .a(_01751_),
    .b(_01752_),
    .y(_01753_)
  );
  al_oa21ttf _06678_ (
    .a(_01749_),
    .b(_01750_),
    .c(_01753_),
    .y(_01754_)
  );
  al_nand3fft _06679_ (
    .a(_01749_),
    .b(_01750_),
    .c(_01753_),
    .y(_01755_)
  );
  al_and3fft _06680_ (
    .a(TM0),
    .b(_01754_),
    .c(_01755_),
    .y(_01756_)
  );
  al_nand2 _06681_ (
    .a(TM0),
    .b(\DFF_551.Q ),
    .y(_01757_)
  );
  al_or3fft _06682_ (
    .a(_01652_),
    .b(_01757_),
    .c(_01756_),
    .y(_01758_)
  );
  al_and2 _06683_ (
    .a(TM0),
    .b(\DFF_408.Q ),
    .y(_01759_)
  );
  al_and3fft _06684_ (
    .a(_01759_),
    .b(_01274_),
    .c(TM1),
    .y(_01760_)
  );
  al_nor3fft _06685_ (
    .a(RESET),
    .b(_01758_),
    .c(_01760_),
    .y(\DFF_440.D )
  );
  al_nor2 _06686_ (
    .a(\DFF_665.Q ),
    .b(\DFF_697.Q ),
    .y(_01761_)
  );
  al_and2 _06687_ (
    .a(\DFF_665.Q ),
    .b(\DFF_697.Q ),
    .y(_01762_)
  );
  al_and2ft _06688_ (
    .a(\DFF_633.Q ),
    .b(\DFF_729.Q ),
    .y(_01763_)
  );
  al_nand2ft _06689_ (
    .a(\DFF_729.Q ),
    .b(\DFF_633.Q ),
    .y(_01764_)
  );
  al_nand2ft _06690_ (
    .a(_01763_),
    .b(_01764_),
    .y(_01765_)
  );
  al_oa21ttf _06691_ (
    .a(_01761_),
    .b(_01762_),
    .c(_01765_),
    .y(_01766_)
  );
  al_nand3fft _06692_ (
    .a(_01761_),
    .b(_01762_),
    .c(_01765_),
    .y(_01767_)
  );
  al_and3fft _06693_ (
    .a(TM0),
    .b(_01766_),
    .c(_01767_),
    .y(_01768_)
  );
  al_nand2 _06694_ (
    .a(TM0),
    .b(\DFF_550.Q ),
    .y(_01769_)
  );
  al_or3fft _06695_ (
    .a(_01652_),
    .b(_01769_),
    .c(_01768_),
    .y(_01770_)
  );
  al_and2 _06696_ (
    .a(TM0),
    .b(\DFF_409.Q ),
    .y(_01771_)
  );
  al_and3fft _06697_ (
    .a(_01771_),
    .b(_01285_),
    .c(TM1),
    .y(_01772_)
  );
  al_nor3fft _06698_ (
    .a(RESET),
    .b(_01770_),
    .c(_01772_),
    .y(\DFF_441.D )
  );
  al_nor2 _06699_ (
    .a(\DFF_666.Q ),
    .b(\DFF_698.Q ),
    .y(_01773_)
  );
  al_and2 _06700_ (
    .a(\DFF_666.Q ),
    .b(\DFF_698.Q ),
    .y(_01774_)
  );
  al_and2ft _06701_ (
    .a(\DFF_634.Q ),
    .b(\DFF_730.Q ),
    .y(_01775_)
  );
  al_nand2ft _06702_ (
    .a(\DFF_730.Q ),
    .b(\DFF_634.Q ),
    .y(_01776_)
  );
  al_nand2ft _06703_ (
    .a(_01775_),
    .b(_01776_),
    .y(_01777_)
  );
  al_oa21ttf _06704_ (
    .a(_01773_),
    .b(_01774_),
    .c(_01777_),
    .y(_01778_)
  );
  al_nand3fft _06705_ (
    .a(_01773_),
    .b(_01774_),
    .c(_01777_),
    .y(_01779_)
  );
  al_and3fft _06706_ (
    .a(TM0),
    .b(_01778_),
    .c(_01779_),
    .y(_01780_)
  );
  al_nand2 _06707_ (
    .a(TM0),
    .b(\DFF_549.Q ),
    .y(_01781_)
  );
  al_or3fft _06708_ (
    .a(_01652_),
    .b(_01781_),
    .c(_01780_),
    .y(_01782_)
  );
  al_and2 _06709_ (
    .a(TM0),
    .b(\DFF_410.Q ),
    .y(_01783_)
  );
  al_and3fft _06710_ (
    .a(_01783_),
    .b(_01296_),
    .c(TM1),
    .y(_01784_)
  );
  al_nor3fft _06711_ (
    .a(RESET),
    .b(_01782_),
    .c(_01784_),
    .y(\DFF_442.D )
  );
  al_nor2 _06712_ (
    .a(\DFF_667.Q ),
    .b(\DFF_699.Q ),
    .y(_01785_)
  );
  al_and2 _06713_ (
    .a(\DFF_667.Q ),
    .b(\DFF_699.Q ),
    .y(_01786_)
  );
  al_and2ft _06714_ (
    .a(\DFF_635.Q ),
    .b(\DFF_731.Q ),
    .y(_01787_)
  );
  al_nand2ft _06715_ (
    .a(\DFF_731.Q ),
    .b(\DFF_635.Q ),
    .y(_01788_)
  );
  al_nand2ft _06716_ (
    .a(_01787_),
    .b(_01788_),
    .y(_01789_)
  );
  al_oa21ttf _06717_ (
    .a(_01785_),
    .b(_01786_),
    .c(_01789_),
    .y(_01790_)
  );
  al_nand3fft _06718_ (
    .a(_01785_),
    .b(_01786_),
    .c(_01789_),
    .y(_01791_)
  );
  al_and3fft _06719_ (
    .a(TM0),
    .b(_01790_),
    .c(_01791_),
    .y(_01792_)
  );
  al_nand2 _06720_ (
    .a(TM0),
    .b(\DFF_548.Q ),
    .y(_01793_)
  );
  al_or3fft _06721_ (
    .a(_01652_),
    .b(_01793_),
    .c(_01792_),
    .y(_01794_)
  );
  al_and2 _06722_ (
    .a(TM0),
    .b(\DFF_411.Q ),
    .y(_01795_)
  );
  al_and3fft _06723_ (
    .a(_01795_),
    .b(_01307_),
    .c(TM1),
    .y(_01796_)
  );
  al_nor3fft _06724_ (
    .a(RESET),
    .b(_01794_),
    .c(_01796_),
    .y(\DFF_443.D )
  );
  al_nor2 _06725_ (
    .a(\DFF_668.Q ),
    .b(\DFF_700.Q ),
    .y(_01797_)
  );
  al_and2 _06726_ (
    .a(\DFF_668.Q ),
    .b(\DFF_700.Q ),
    .y(_01798_)
  );
  al_and2ft _06727_ (
    .a(\DFF_636.Q ),
    .b(\DFF_732.Q ),
    .y(_01799_)
  );
  al_nand2ft _06728_ (
    .a(\DFF_732.Q ),
    .b(\DFF_636.Q ),
    .y(_01800_)
  );
  al_nand2ft _06729_ (
    .a(_01799_),
    .b(_01800_),
    .y(_01801_)
  );
  al_oa21ttf _06730_ (
    .a(_01797_),
    .b(_01798_),
    .c(_01801_),
    .y(_01802_)
  );
  al_nand3fft _06731_ (
    .a(_01797_),
    .b(_01798_),
    .c(_01801_),
    .y(_01803_)
  );
  al_and3fft _06732_ (
    .a(TM0),
    .b(_01802_),
    .c(_01803_),
    .y(_01804_)
  );
  al_nand2 _06733_ (
    .a(TM0),
    .b(\DFF_547.Q ),
    .y(_01805_)
  );
  al_or3fft _06734_ (
    .a(_01652_),
    .b(_01805_),
    .c(_01804_),
    .y(_01806_)
  );
  al_and2 _06735_ (
    .a(TM0),
    .b(\DFF_412.Q ),
    .y(_01807_)
  );
  al_and3fft _06736_ (
    .a(_01807_),
    .b(_01318_),
    .c(TM1),
    .y(_01808_)
  );
  al_nor3fft _06737_ (
    .a(RESET),
    .b(_01806_),
    .c(_01808_),
    .y(\DFF_444.D )
  );
  al_nor2 _06738_ (
    .a(\DFF_669.Q ),
    .b(\DFF_701.Q ),
    .y(_01809_)
  );
  al_and2 _06739_ (
    .a(\DFF_669.Q ),
    .b(\DFF_701.Q ),
    .y(_01810_)
  );
  al_and2ft _06740_ (
    .a(\DFF_637.Q ),
    .b(\DFF_733.Q ),
    .y(_01811_)
  );
  al_nand2ft _06741_ (
    .a(\DFF_733.Q ),
    .b(\DFF_637.Q ),
    .y(_01812_)
  );
  al_nand2ft _06742_ (
    .a(_01811_),
    .b(_01812_),
    .y(_01813_)
  );
  al_oa21ttf _06743_ (
    .a(_01809_),
    .b(_01810_),
    .c(_01813_),
    .y(_01814_)
  );
  al_nand3fft _06744_ (
    .a(_01809_),
    .b(_01810_),
    .c(_01813_),
    .y(_01815_)
  );
  al_and3fft _06745_ (
    .a(TM0),
    .b(_01814_),
    .c(_01815_),
    .y(_01816_)
  );
  al_nand2 _06746_ (
    .a(TM0),
    .b(\DFF_546.Q ),
    .y(_01817_)
  );
  al_or3fft _06747_ (
    .a(_01652_),
    .b(_01817_),
    .c(_01816_),
    .y(_01818_)
  );
  al_and2 _06748_ (
    .a(TM0),
    .b(\DFF_413.Q ),
    .y(_01819_)
  );
  al_and3fft _06749_ (
    .a(_01819_),
    .b(_01329_),
    .c(TM1),
    .y(_01820_)
  );
  al_nor3fft _06750_ (
    .a(RESET),
    .b(_01818_),
    .c(_01820_),
    .y(\DFF_445.D )
  );
  al_nor2 _06751_ (
    .a(\DFF_670.Q ),
    .b(\DFF_702.Q ),
    .y(_01821_)
  );
  al_and2 _06752_ (
    .a(\DFF_670.Q ),
    .b(\DFF_702.Q ),
    .y(_01822_)
  );
  al_and2ft _06753_ (
    .a(\DFF_638.Q ),
    .b(\DFF_734.Q ),
    .y(_01823_)
  );
  al_nand2ft _06754_ (
    .a(\DFF_734.Q ),
    .b(\DFF_638.Q ),
    .y(_01824_)
  );
  al_nand2ft _06755_ (
    .a(_01823_),
    .b(_01824_),
    .y(_01825_)
  );
  al_oa21ttf _06756_ (
    .a(_01821_),
    .b(_01822_),
    .c(_01825_),
    .y(_01826_)
  );
  al_nand3fft _06757_ (
    .a(_01821_),
    .b(_01822_),
    .c(_01825_),
    .y(_01827_)
  );
  al_and3fft _06758_ (
    .a(TM0),
    .b(_01826_),
    .c(_01827_),
    .y(_01828_)
  );
  al_nand2 _06759_ (
    .a(TM0),
    .b(\DFF_545.Q ),
    .y(_01829_)
  );
  al_or3fft _06760_ (
    .a(_01652_),
    .b(_01829_),
    .c(_01828_),
    .y(_01830_)
  );
  al_and2 _06761_ (
    .a(TM0),
    .b(\DFF_414.Q ),
    .y(_01831_)
  );
  al_and3fft _06762_ (
    .a(_01831_),
    .b(_01340_),
    .c(TM1),
    .y(_01832_)
  );
  al_nor3fft _06763_ (
    .a(RESET),
    .b(_01830_),
    .c(_01832_),
    .y(\DFF_446.D )
  );
  al_nor2 _06764_ (
    .a(\DFF_671.Q ),
    .b(\DFF_703.Q ),
    .y(_01833_)
  );
  al_and2 _06765_ (
    .a(\DFF_671.Q ),
    .b(\DFF_703.Q ),
    .y(_01834_)
  );
  al_and2ft _06766_ (
    .a(\DFF_639.Q ),
    .b(\DFF_735.Q ),
    .y(_01835_)
  );
  al_nand2ft _06767_ (
    .a(\DFF_735.Q ),
    .b(\DFF_639.Q ),
    .y(_01836_)
  );
  al_nand2ft _06768_ (
    .a(_01835_),
    .b(_01836_),
    .y(_01837_)
  );
  al_oa21ttf _06769_ (
    .a(_01833_),
    .b(_01834_),
    .c(_01837_),
    .y(_01838_)
  );
  al_nand3fft _06770_ (
    .a(_01833_),
    .b(_01834_),
    .c(_01837_),
    .y(_01839_)
  );
  al_and3fft _06771_ (
    .a(TM0),
    .b(_01838_),
    .c(_01839_),
    .y(_01840_)
  );
  al_nand2 _06772_ (
    .a(TM0),
    .b(\DFF_544.Q ),
    .y(_01841_)
  );
  al_or3fft _06773_ (
    .a(_01652_),
    .b(_01841_),
    .c(_01840_),
    .y(_01842_)
  );
  al_and2 _06774_ (
    .a(TM0),
    .b(\DFF_415.Q ),
    .y(_01843_)
  );
  al_and3fft _06775_ (
    .a(_01843_),
    .b(_01351_),
    .c(TM1),
    .y(_01844_)
  );
  al_nor3fft _06776_ (
    .a(RESET),
    .b(_01842_),
    .c(_01844_),
    .y(\DFF_447.D )
  );
  al_and2 _06777_ (
    .a(RESET),
    .b(\DFF_416.Q ),
    .y(\DFF_448.D )
  );
  al_and2 _06778_ (
    .a(RESET),
    .b(\DFF_417.Q ),
    .y(\DFF_449.D )
  );
  al_and2 _06779_ (
    .a(RESET),
    .b(\DFF_418.Q ),
    .y(\DFF_450.D )
  );
  al_and2 _06780_ (
    .a(RESET),
    .b(\DFF_419.Q ),
    .y(\DFF_451.D )
  );
  al_and2 _06781_ (
    .a(RESET),
    .b(\DFF_420.Q ),
    .y(\DFF_452.D )
  );
  al_and2 _06782_ (
    .a(RESET),
    .b(\DFF_421.Q ),
    .y(\DFF_453.D )
  );
  al_and2 _06783_ (
    .a(RESET),
    .b(\DFF_422.Q ),
    .y(\DFF_454.D )
  );
  al_and2 _06784_ (
    .a(RESET),
    .b(\DFF_423.Q ),
    .y(\DFF_455.D )
  );
  al_and2 _06785_ (
    .a(RESET),
    .b(\DFF_424.Q ),
    .y(\DFF_456.D )
  );
  al_and2 _06786_ (
    .a(RESET),
    .b(\DFF_425.Q ),
    .y(\DFF_457.D )
  );
  al_and2 _06787_ (
    .a(RESET),
    .b(\DFF_426.Q ),
    .y(\DFF_458.D )
  );
  al_and2 _06788_ (
    .a(RESET),
    .b(\DFF_427.Q ),
    .y(\DFF_459.D )
  );
  al_and2 _06789_ (
    .a(RESET),
    .b(\DFF_428.Q ),
    .y(\DFF_460.D )
  );
  al_and2 _06790_ (
    .a(RESET),
    .b(\DFF_429.Q ),
    .y(\DFF_461.D )
  );
  al_and2 _06791_ (
    .a(RESET),
    .b(\DFF_430.Q ),
    .y(\DFF_462.D )
  );
  al_and2 _06792_ (
    .a(RESET),
    .b(\DFF_431.Q ),
    .y(\DFF_463.D )
  );
  al_and2 _06793_ (
    .a(RESET),
    .b(\DFF_432.Q ),
    .y(\DFF_464.D )
  );
  al_and2 _06794_ (
    .a(RESET),
    .b(\DFF_433.Q ),
    .y(\DFF_465.D )
  );
  al_and2 _06795_ (
    .a(RESET),
    .b(\DFF_434.Q ),
    .y(\DFF_466.D )
  );
  al_and2 _06796_ (
    .a(RESET),
    .b(\DFF_435.Q ),
    .y(\DFF_467.D )
  );
  al_and2 _06797_ (
    .a(RESET),
    .b(\DFF_436.Q ),
    .y(\DFF_468.D )
  );
  al_and2 _06798_ (
    .a(RESET),
    .b(\DFF_437.Q ),
    .y(\DFF_469.D )
  );
  al_and2 _06799_ (
    .a(RESET),
    .b(\DFF_438.Q ),
    .y(\DFF_470.D )
  );
  al_and2 _06800_ (
    .a(RESET),
    .b(\DFF_439.Q ),
    .y(\DFF_471.D )
  );
  al_and2 _06801_ (
    .a(RESET),
    .b(\DFF_440.Q ),
    .y(\DFF_472.D )
  );
  al_and2 _06802_ (
    .a(RESET),
    .b(\DFF_441.Q ),
    .y(\DFF_473.D )
  );
  al_and2 _06803_ (
    .a(RESET),
    .b(\DFF_442.Q ),
    .y(\DFF_474.D )
  );
  al_and2 _06804_ (
    .a(RESET),
    .b(\DFF_443.Q ),
    .y(\DFF_475.D )
  );
  al_and2 _06805_ (
    .a(RESET),
    .b(\DFF_444.Q ),
    .y(\DFF_476.D )
  );
  al_and2 _06806_ (
    .a(RESET),
    .b(\DFF_445.Q ),
    .y(\DFF_477.D )
  );
  al_and2 _06807_ (
    .a(RESET),
    .b(\DFF_446.Q ),
    .y(\DFF_478.D )
  );
  al_and2 _06808_ (
    .a(RESET),
    .b(\DFF_447.Q ),
    .y(\DFF_479.D )
  );
  al_and2 _06809_ (
    .a(RESET),
    .b(\DFF_448.Q ),
    .y(\DFF_480.D )
  );
  al_and2 _06810_ (
    .a(RESET),
    .b(\DFF_449.Q ),
    .y(\DFF_481.D )
  );
  al_and2 _06811_ (
    .a(RESET),
    .b(\DFF_450.Q ),
    .y(\DFF_482.D )
  );
  al_and2 _06812_ (
    .a(RESET),
    .b(\DFF_451.Q ),
    .y(\DFF_483.D )
  );
  al_and2 _06813_ (
    .a(RESET),
    .b(\DFF_452.Q ),
    .y(\DFF_484.D )
  );
  al_and2 _06814_ (
    .a(RESET),
    .b(\DFF_453.Q ),
    .y(\DFF_485.D )
  );
  al_and2 _06815_ (
    .a(RESET),
    .b(\DFF_454.Q ),
    .y(\DFF_486.D )
  );
  al_and2 _06816_ (
    .a(RESET),
    .b(\DFF_455.Q ),
    .y(\DFF_487.D )
  );
  al_and2 _06817_ (
    .a(RESET),
    .b(\DFF_456.Q ),
    .y(\DFF_488.D )
  );
  al_and2 _06818_ (
    .a(RESET),
    .b(\DFF_457.Q ),
    .y(\DFF_489.D )
  );
  al_and2 _06819_ (
    .a(RESET),
    .b(\DFF_458.Q ),
    .y(\DFF_490.D )
  );
  al_and2 _06820_ (
    .a(RESET),
    .b(\DFF_459.Q ),
    .y(\DFF_491.D )
  );
  al_and2 _06821_ (
    .a(RESET),
    .b(\DFF_460.Q ),
    .y(\DFF_492.D )
  );
  al_and2 _06822_ (
    .a(RESET),
    .b(\DFF_461.Q ),
    .y(\DFF_493.D )
  );
  al_and2 _06823_ (
    .a(RESET),
    .b(\DFF_462.Q ),
    .y(\DFF_494.D )
  );
  al_and2 _06824_ (
    .a(RESET),
    .b(\DFF_463.Q ),
    .y(\DFF_495.D )
  );
  al_and2 _06825_ (
    .a(RESET),
    .b(\DFF_464.Q ),
    .y(\DFF_496.D )
  );
  al_and2 _06826_ (
    .a(RESET),
    .b(\DFF_465.Q ),
    .y(\DFF_497.D )
  );
  al_and2 _06827_ (
    .a(RESET),
    .b(\DFF_466.Q ),
    .y(\DFF_498.D )
  );
  al_and2 _06828_ (
    .a(RESET),
    .b(\DFF_467.Q ),
    .y(\DFF_499.D )
  );
  al_and2 _06829_ (
    .a(RESET),
    .b(\DFF_468.Q ),
    .y(\DFF_500.D )
  );
  al_and2 _06830_ (
    .a(RESET),
    .b(\DFF_469.Q ),
    .y(\DFF_501.D )
  );
  al_and2 _06831_ (
    .a(RESET),
    .b(\DFF_470.Q ),
    .y(\DFF_502.D )
  );
  al_and2 _06832_ (
    .a(RESET),
    .b(\DFF_471.Q ),
    .y(\DFF_503.D )
  );
  al_and2 _06833_ (
    .a(RESET),
    .b(\DFF_472.Q ),
    .y(\DFF_504.D )
  );
  al_and2 _06834_ (
    .a(RESET),
    .b(\DFF_473.Q ),
    .y(\DFF_505.D )
  );
  al_and2 _06835_ (
    .a(RESET),
    .b(\DFF_474.Q ),
    .y(\DFF_506.D )
  );
  al_and2 _06836_ (
    .a(RESET),
    .b(\DFF_475.Q ),
    .y(\DFF_507.D )
  );
  al_and2 _06837_ (
    .a(RESET),
    .b(\DFF_476.Q ),
    .y(\DFF_508.D )
  );
  al_and2 _06838_ (
    .a(RESET),
    .b(\DFF_477.Q ),
    .y(\DFF_509.D )
  );
  al_and2 _06839_ (
    .a(RESET),
    .b(\DFF_478.Q ),
    .y(\DFF_510.D )
  );
  al_and2 _06840_ (
    .a(RESET),
    .b(\DFF_479.Q ),
    .y(\DFF_511.D )
  );
  al_and2 _06841_ (
    .a(RESET),
    .b(\DFF_480.Q ),
    .y(\DFF_512.D )
  );
  al_and2 _06842_ (
    .a(RESET),
    .b(\DFF_481.Q ),
    .y(\DFF_513.D )
  );
  al_and2 _06843_ (
    .a(RESET),
    .b(\DFF_482.Q ),
    .y(\DFF_514.D )
  );
  al_and2 _06844_ (
    .a(RESET),
    .b(\DFF_483.Q ),
    .y(\DFF_515.D )
  );
  al_and2 _06845_ (
    .a(RESET),
    .b(\DFF_484.Q ),
    .y(\DFF_516.D )
  );
  al_and2 _06846_ (
    .a(RESET),
    .b(\DFF_485.Q ),
    .y(\DFF_517.D )
  );
  al_and2 _06847_ (
    .a(RESET),
    .b(\DFF_486.Q ),
    .y(\DFF_518.D )
  );
  al_and2 _06848_ (
    .a(RESET),
    .b(\DFF_487.Q ),
    .y(\DFF_519.D )
  );
  al_and2 _06849_ (
    .a(RESET),
    .b(\DFF_488.Q ),
    .y(\DFF_520.D )
  );
  al_and2 _06850_ (
    .a(RESET),
    .b(\DFF_489.Q ),
    .y(\DFF_521.D )
  );
  al_and2 _06851_ (
    .a(RESET),
    .b(\DFF_490.Q ),
    .y(\DFF_522.D )
  );
  al_and2 _06852_ (
    .a(RESET),
    .b(\DFF_491.Q ),
    .y(\DFF_523.D )
  );
  al_and2 _06853_ (
    .a(RESET),
    .b(\DFF_492.Q ),
    .y(\DFF_524.D )
  );
  al_and2 _06854_ (
    .a(RESET),
    .b(\DFF_493.Q ),
    .y(\DFF_525.D )
  );
  al_and2 _06855_ (
    .a(RESET),
    .b(\DFF_494.Q ),
    .y(\DFF_526.D )
  );
  al_and2 _06856_ (
    .a(RESET),
    .b(\DFF_495.Q ),
    .y(\DFF_527.D )
  );
  al_and2 _06857_ (
    .a(RESET),
    .b(\DFF_496.Q ),
    .y(\DFF_528.D )
  );
  al_and2 _06858_ (
    .a(RESET),
    .b(\DFF_497.Q ),
    .y(\DFF_529.D )
  );
  al_and2 _06859_ (
    .a(RESET),
    .b(\DFF_498.Q ),
    .y(\DFF_530.D )
  );
  al_and2 _06860_ (
    .a(RESET),
    .b(\DFF_499.Q ),
    .y(\DFF_531.D )
  );
  al_and2 _06861_ (
    .a(RESET),
    .b(\DFF_500.Q ),
    .y(\DFF_532.D )
  );
  al_and2 _06862_ (
    .a(RESET),
    .b(\DFF_501.Q ),
    .y(\DFF_533.D )
  );
  al_and2 _06863_ (
    .a(RESET),
    .b(\DFF_502.Q ),
    .y(\DFF_534.D )
  );
  al_and2 _06864_ (
    .a(RESET),
    .b(\DFF_503.Q ),
    .y(\DFF_535.D )
  );
  al_and2 _06865_ (
    .a(RESET),
    .b(\DFF_504.Q ),
    .y(\DFF_536.D )
  );
  al_and2 _06866_ (
    .a(RESET),
    .b(\DFF_505.Q ),
    .y(\DFF_537.D )
  );
  al_and2 _06867_ (
    .a(RESET),
    .b(\DFF_506.Q ),
    .y(\DFF_538.D )
  );
  al_and2 _06868_ (
    .a(RESET),
    .b(\DFF_507.Q ),
    .y(\DFF_539.D )
  );
  al_and2 _06869_ (
    .a(RESET),
    .b(\DFF_508.Q ),
    .y(\DFF_540.D )
  );
  al_and2 _06870_ (
    .a(RESET),
    .b(\DFF_509.Q ),
    .y(\DFF_541.D )
  );
  al_and2 _06871_ (
    .a(RESET),
    .b(\DFF_510.Q ),
    .y(\DFF_542.D )
  );
  al_and2 _06872_ (
    .a(RESET),
    .b(\DFF_511.Q ),
    .y(\DFF_543.D )
  );
  al_oa21ftt _06873_ (
    .a(\DFF_543.Q ),
    .b(\DFF_575.Q ),
    .c(RESET),
    .y(_01845_)
  );
  al_aoi21ftf _06874_ (
    .a(\DFF_543.Q ),
    .b(\DFF_575.Q ),
    .c(_01845_),
    .y(\DFF_544.D )
  );
  al_oa21ftt _06875_ (
    .a(\DFF_542.Q ),
    .b(\DFF_544.Q ),
    .c(RESET),
    .y(_01846_)
  );
  al_aoi21ftf _06876_ (
    .a(\DFF_542.Q ),
    .b(\DFF_544.Q ),
    .c(_01846_),
    .y(\DFF_545.D )
  );
  al_oa21ftt _06877_ (
    .a(\DFF_541.Q ),
    .b(\DFF_545.Q ),
    .c(RESET),
    .y(_01847_)
  );
  al_aoi21ftf _06878_ (
    .a(\DFF_541.Q ),
    .b(\DFF_545.Q ),
    .c(_01847_),
    .y(\DFF_546.D )
  );
  al_oa21ftt _06879_ (
    .a(\DFF_540.Q ),
    .b(\DFF_546.Q ),
    .c(RESET),
    .y(_01848_)
  );
  al_aoi21ftf _06880_ (
    .a(\DFF_540.Q ),
    .b(\DFF_546.Q ),
    .c(_01848_),
    .y(\DFF_547.D )
  );
  al_nand2ft _06881_ (
    .a(\DFF_539.Q ),
    .b(\DFF_547.Q ),
    .y(_01849_)
  );
  al_nand2ft _06882_ (
    .a(\DFF_547.Q ),
    .b(\DFF_539.Q ),
    .y(_01850_)
  );
  al_ao21ttf _06883_ (
    .a(_01849_),
    .b(_01850_),
    .c(\DFF_575.Q ),
    .y(_01851_)
  );
  al_nand3ftt _06884_ (
    .a(\DFF_575.Q ),
    .b(_01849_),
    .c(_01850_),
    .y(_01852_)
  );
  al_aoi21 _06885_ (
    .a(_01852_),
    .b(_01851_),
    .c(_00451_),
    .y(\DFF_548.D )
  );
  al_oa21ftt _06886_ (
    .a(\DFF_538.Q ),
    .b(\DFF_548.Q ),
    .c(RESET),
    .y(_01853_)
  );
  al_aoi21ftf _06887_ (
    .a(\DFF_538.Q ),
    .b(\DFF_548.Q ),
    .c(_01853_),
    .y(\DFF_549.D )
  );
  al_oa21ftt _06888_ (
    .a(\DFF_537.Q ),
    .b(\DFF_549.Q ),
    .c(RESET),
    .y(_01854_)
  );
  al_aoi21ftf _06889_ (
    .a(\DFF_537.Q ),
    .b(\DFF_549.Q ),
    .c(_01854_),
    .y(\DFF_550.D )
  );
  al_oa21ftt _06890_ (
    .a(\DFF_536.Q ),
    .b(\DFF_550.Q ),
    .c(RESET),
    .y(_01855_)
  );
  al_aoi21ftf _06891_ (
    .a(\DFF_536.Q ),
    .b(\DFF_550.Q ),
    .c(_01855_),
    .y(\DFF_551.D )
  );
  al_oa21ftt _06892_ (
    .a(\DFF_535.Q ),
    .b(\DFF_551.Q ),
    .c(RESET),
    .y(_01856_)
  );
  al_aoi21ftf _06893_ (
    .a(\DFF_535.Q ),
    .b(\DFF_551.Q ),
    .c(_01856_),
    .y(\DFF_552.D )
  );
  al_oa21ftt _06894_ (
    .a(\DFF_534.Q ),
    .b(\DFF_552.Q ),
    .c(RESET),
    .y(_01857_)
  );
  al_aoi21ftf _06895_ (
    .a(\DFF_534.Q ),
    .b(\DFF_552.Q ),
    .c(_01857_),
    .y(\DFF_553.D )
  );
  al_oa21ftt _06896_ (
    .a(\DFF_533.Q ),
    .b(\DFF_553.Q ),
    .c(RESET),
    .y(_01858_)
  );
  al_aoi21ftf _06897_ (
    .a(\DFF_533.Q ),
    .b(\DFF_553.Q ),
    .c(_01858_),
    .y(\DFF_554.D )
  );
  al_nand2ft _06898_ (
    .a(\DFF_532.Q ),
    .b(\DFF_554.Q ),
    .y(_01859_)
  );
  al_nand2ft _06899_ (
    .a(\DFF_554.Q ),
    .b(\DFF_532.Q ),
    .y(_01860_)
  );
  al_ao21ttf _06900_ (
    .a(_01859_),
    .b(_01860_),
    .c(\DFF_575.Q ),
    .y(_01861_)
  );
  al_nand3ftt _06901_ (
    .a(\DFF_575.Q ),
    .b(_01859_),
    .c(_01860_),
    .y(_01862_)
  );
  al_aoi21 _06902_ (
    .a(_01862_),
    .b(_01861_),
    .c(_00451_),
    .y(\DFF_555.D )
  );
  al_oa21ftt _06903_ (
    .a(\DFF_531.Q ),
    .b(\DFF_555.Q ),
    .c(RESET),
    .y(_01863_)
  );
  al_aoi21ftf _06904_ (
    .a(\DFF_531.Q ),
    .b(\DFF_555.Q ),
    .c(_01863_),
    .y(\DFF_556.D )
  );
  al_oa21ftt _06905_ (
    .a(\DFF_530.Q ),
    .b(\DFF_556.Q ),
    .c(RESET),
    .y(_01864_)
  );
  al_aoi21ftf _06906_ (
    .a(\DFF_530.Q ),
    .b(\DFF_556.Q ),
    .c(_01864_),
    .y(\DFF_557.D )
  );
  al_oa21ftt _06907_ (
    .a(\DFF_529.Q ),
    .b(\DFF_557.Q ),
    .c(RESET),
    .y(_01865_)
  );
  al_aoi21ftf _06908_ (
    .a(\DFF_529.Q ),
    .b(\DFF_557.Q ),
    .c(_01865_),
    .y(\DFF_558.D )
  );
  al_oa21ftt _06909_ (
    .a(\DFF_528.Q ),
    .b(\DFF_558.Q ),
    .c(RESET),
    .y(_01866_)
  );
  al_aoi21ftf _06910_ (
    .a(\DFF_528.Q ),
    .b(\DFF_558.Q ),
    .c(_01866_),
    .y(\DFF_559.D )
  );
  al_nand2ft _06911_ (
    .a(\DFF_527.Q ),
    .b(\DFF_559.Q ),
    .y(_01867_)
  );
  al_nand2ft _06912_ (
    .a(\DFF_559.Q ),
    .b(\DFF_527.Q ),
    .y(_01868_)
  );
  al_ao21ttf _06913_ (
    .a(_01867_),
    .b(_01868_),
    .c(\DFF_575.Q ),
    .y(_01869_)
  );
  al_nand3ftt _06914_ (
    .a(\DFF_575.Q ),
    .b(_01867_),
    .c(_01868_),
    .y(_01870_)
  );
  al_aoi21 _06915_ (
    .a(_01870_),
    .b(_01869_),
    .c(_00451_),
    .y(\DFF_560.D )
  );
  al_oa21ftt _06916_ (
    .a(\DFF_526.Q ),
    .b(\DFF_560.Q ),
    .c(RESET),
    .y(_01871_)
  );
  al_aoi21ftf _06917_ (
    .a(\DFF_526.Q ),
    .b(\DFF_560.Q ),
    .c(_01871_),
    .y(\DFF_561.D )
  );
  al_oa21ftt _06918_ (
    .a(\DFF_525.Q ),
    .b(\DFF_561.Q ),
    .c(RESET),
    .y(_01872_)
  );
  al_aoi21ftf _06919_ (
    .a(\DFF_525.Q ),
    .b(\DFF_561.Q ),
    .c(_01872_),
    .y(\DFF_562.D )
  );
  al_oa21ftt _06920_ (
    .a(\DFF_524.Q ),
    .b(\DFF_562.Q ),
    .c(RESET),
    .y(_01873_)
  );
  al_aoi21ftf _06921_ (
    .a(\DFF_524.Q ),
    .b(\DFF_562.Q ),
    .c(_01873_),
    .y(\DFF_563.D )
  );
  al_oa21ftt _06922_ (
    .a(\DFF_523.Q ),
    .b(\DFF_563.Q ),
    .c(RESET),
    .y(_01874_)
  );
  al_aoi21ftf _06923_ (
    .a(\DFF_523.Q ),
    .b(\DFF_563.Q ),
    .c(_01874_),
    .y(\DFF_564.D )
  );
  al_oa21ftt _06924_ (
    .a(\DFF_522.Q ),
    .b(\DFF_564.Q ),
    .c(RESET),
    .y(_01875_)
  );
  al_aoi21ftf _06925_ (
    .a(\DFF_522.Q ),
    .b(\DFF_564.Q ),
    .c(_01875_),
    .y(\DFF_565.D )
  );
  al_oa21ftt _06926_ (
    .a(\DFF_521.Q ),
    .b(\DFF_565.Q ),
    .c(RESET),
    .y(_01876_)
  );
  al_aoi21ftf _06927_ (
    .a(\DFF_521.Q ),
    .b(\DFF_565.Q ),
    .c(_01876_),
    .y(\DFF_566.D )
  );
  al_oa21ftt _06928_ (
    .a(\DFF_520.Q ),
    .b(\DFF_566.Q ),
    .c(RESET),
    .y(_01877_)
  );
  al_aoi21ftf _06929_ (
    .a(\DFF_520.Q ),
    .b(\DFF_566.Q ),
    .c(_01877_),
    .y(\DFF_567.D )
  );
  al_oa21ftt _06930_ (
    .a(\DFF_519.Q ),
    .b(\DFF_567.Q ),
    .c(RESET),
    .y(_01878_)
  );
  al_aoi21ftf _06931_ (
    .a(\DFF_519.Q ),
    .b(\DFF_567.Q ),
    .c(_01878_),
    .y(\DFF_568.D )
  );
  al_oa21ftt _06932_ (
    .a(\DFF_518.Q ),
    .b(\DFF_568.Q ),
    .c(RESET),
    .y(_01879_)
  );
  al_aoi21ftf _06933_ (
    .a(\DFF_518.Q ),
    .b(\DFF_568.Q ),
    .c(_01879_),
    .y(\DFF_569.D )
  );
  al_oa21ftt _06934_ (
    .a(\DFF_517.Q ),
    .b(\DFF_569.Q ),
    .c(RESET),
    .y(_01880_)
  );
  al_aoi21ftf _06935_ (
    .a(\DFF_517.Q ),
    .b(\DFF_569.Q ),
    .c(_01880_),
    .y(\DFF_570.D )
  );
  al_oa21ftt _06936_ (
    .a(\DFF_516.Q ),
    .b(\DFF_570.Q ),
    .c(RESET),
    .y(_01881_)
  );
  al_aoi21ftf _06937_ (
    .a(\DFF_516.Q ),
    .b(\DFF_570.Q ),
    .c(_01881_),
    .y(\DFF_571.D )
  );
  al_oa21ftt _06938_ (
    .a(\DFF_515.Q ),
    .b(\DFF_571.Q ),
    .c(RESET),
    .y(_01882_)
  );
  al_aoi21ftf _06939_ (
    .a(\DFF_515.Q ),
    .b(\DFF_571.Q ),
    .c(_01882_),
    .y(\DFF_572.D )
  );
  al_oa21ftt _06940_ (
    .a(\DFF_514.Q ),
    .b(\DFF_572.Q ),
    .c(RESET),
    .y(_01883_)
  );
  al_aoi21ftf _06941_ (
    .a(\DFF_514.Q ),
    .b(\DFF_572.Q ),
    .c(_01883_),
    .y(\DFF_573.D )
  );
  al_oa21ftt _06942_ (
    .a(\DFF_513.Q ),
    .b(\DFF_573.Q ),
    .c(RESET),
    .y(_01884_)
  );
  al_aoi21ftf _06943_ (
    .a(\DFF_513.Q ),
    .b(\DFF_573.Q ),
    .c(_01884_),
    .y(\DFF_574.D )
  );
  al_oa21ftt _06944_ (
    .a(\DFF_512.Q ),
    .b(\DFF_574.Q ),
    .c(RESET),
    .y(_01885_)
  );
  al_aoi21ftf _06945_ (
    .a(\DFF_512.Q ),
    .b(\DFF_574.Q ),
    .c(_01885_),
    .y(\DFF_575.D )
  );
  al_and2 _06946_ (
    .a(RESET),
    .b(\DFF_577.Q ),
    .y(\DFF_576.D )
  );
  al_and2 _06947_ (
    .a(RESET),
    .b(\DFF_578.Q ),
    .y(\DFF_577.D )
  );
  al_and2 _06948_ (
    .a(RESET),
    .b(\DFF_579.Q ),
    .y(\DFF_578.D )
  );
  al_and2 _06949_ (
    .a(RESET),
    .b(\DFF_580.Q ),
    .y(\DFF_579.D )
  );
  al_and2 _06950_ (
    .a(RESET),
    .b(\DFF_581.Q ),
    .y(\DFF_580.D )
  );
  al_and2 _06951_ (
    .a(RESET),
    .b(\DFF_582.Q ),
    .y(\DFF_581.D )
  );
  al_and2 _06952_ (
    .a(RESET),
    .b(\DFF_583.Q ),
    .y(\DFF_582.D )
  );
  al_and2 _06953_ (
    .a(RESET),
    .b(\DFF_584.Q ),
    .y(\DFF_583.D )
  );
  al_and2 _06954_ (
    .a(RESET),
    .b(\DFF_585.Q ),
    .y(\DFF_584.D )
  );
  al_and2 _06955_ (
    .a(RESET),
    .b(\DFF_586.Q ),
    .y(\DFF_585.D )
  );
  al_and2 _06956_ (
    .a(RESET),
    .b(\DFF_587.Q ),
    .y(\DFF_586.D )
  );
  al_and2 _06957_ (
    .a(RESET),
    .b(\DFF_588.Q ),
    .y(\DFF_587.D )
  );
  al_and2 _06958_ (
    .a(RESET),
    .b(\DFF_589.Q ),
    .y(\DFF_588.D )
  );
  al_and2 _06959_ (
    .a(RESET),
    .b(\DFF_590.Q ),
    .y(\DFF_589.D )
  );
  al_and2 _06960_ (
    .a(RESET),
    .b(\DFF_591.Q ),
    .y(\DFF_590.D )
  );
  al_and2 _06961_ (
    .a(RESET),
    .b(\DFF_592.Q ),
    .y(\DFF_591.D )
  );
  al_and2 _06962_ (
    .a(RESET),
    .b(\DFF_593.Q ),
    .y(\DFF_592.D )
  );
  al_and2 _06963_ (
    .a(RESET),
    .b(\DFF_594.Q ),
    .y(\DFF_593.D )
  );
  al_and2 _06964_ (
    .a(RESET),
    .b(\DFF_595.Q ),
    .y(\DFF_594.D )
  );
  al_and2 _06965_ (
    .a(RESET),
    .b(\DFF_596.Q ),
    .y(\DFF_595.D )
  );
  al_and2 _06966_ (
    .a(RESET),
    .b(\DFF_597.Q ),
    .y(\DFF_596.D )
  );
  al_and2 _06967_ (
    .a(RESET),
    .b(\DFF_598.Q ),
    .y(\DFF_597.D )
  );
  al_and2 _06968_ (
    .a(RESET),
    .b(\DFF_599.Q ),
    .y(\DFF_598.D )
  );
  al_and2 _06969_ (
    .a(RESET),
    .b(\DFF_600.Q ),
    .y(\DFF_599.D )
  );
  al_and2 _06970_ (
    .a(RESET),
    .b(\DFF_601.Q ),
    .y(\DFF_600.D )
  );
  al_and2 _06971_ (
    .a(RESET),
    .b(\DFF_602.Q ),
    .y(\DFF_601.D )
  );
  al_and2 _06972_ (
    .a(RESET),
    .b(\DFF_603.Q ),
    .y(\DFF_602.D )
  );
  al_and2 _06973_ (
    .a(RESET),
    .b(\DFF_604.Q ),
    .y(\DFF_603.D )
  );
  al_and2 _06974_ (
    .a(RESET),
    .b(\DFF_605.Q ),
    .y(\DFF_604.D )
  );
  al_and2 _06975_ (
    .a(RESET),
    .b(\DFF_606.Q ),
    .y(\DFF_605.D )
  );
  al_and2 _06976_ (
    .a(RESET),
    .b(\DFF_607.Q ),
    .y(\DFF_606.D )
  );
  al_and2ft _06977_ (
    .a(\DFF_576.Q ),
    .b(RESET),
    .y(\DFF_607.D )
  );
  al_or2 _06978_ (
    .a(TM1),
    .b(\DFF_864.Q ),
    .y(_01886_)
  );
  al_nand2 _06979_ (
    .a(TM1),
    .b(\DFF_864.Q ),
    .y(_01887_)
  );
  al_nand3 _06980_ (
    .a(\DFF_896.Q ),
    .b(_01886_),
    .c(_01887_),
    .y(_01888_)
  );
  al_nand2ft _06981_ (
    .a(TM1),
    .b(\DFF_864.Q ),
    .y(_01889_)
  );
  al_and2ft _06982_ (
    .a(\DFF_864.Q ),
    .b(TM1),
    .y(_01890_)
  );
  al_and3fft _06983_ (
    .a(\DFF_896.Q ),
    .b(_01890_),
    .c(_01889_),
    .y(_01891_)
  );
  al_and2ft _06984_ (
    .a(\DFF_832.Q ),
    .b(\DFF_800.Q ),
    .y(_01892_)
  );
  al_nand2ft _06985_ (
    .a(\DFF_800.Q ),
    .b(\DFF_832.Q ),
    .y(_01893_)
  );
  al_nand2ft _06986_ (
    .a(_01892_),
    .b(_01893_),
    .y(_01894_)
  );
  al_oai21ftf _06987_ (
    .a(_01888_),
    .b(_01891_),
    .c(_01894_),
    .y(_01895_)
  );
  al_nand3ftt _06988_ (
    .a(_01891_),
    .b(_01888_),
    .c(_01894_),
    .y(_01896_)
  );
  al_nand3 _06989_ (
    .a(_00448_),
    .b(_01895_),
    .c(_01896_),
    .y(_01897_)
  );
  al_aoi21 _06990_ (
    .a(TM0),
    .b(\DFF_767.Q ),
    .c(TM1),
    .y(_01898_)
  );
  al_nand2 _06991_ (
    .a(_01898_),
    .b(_01897_),
    .y(_01899_)
  );
  al_aoi21ttf _06992_ (
    .a(\DFF_576.Q ),
    .b(TM0),
    .c(TM1),
    .y(_01900_)
  );
  al_and2 _06993_ (
    .a(_01900_),
    .b(_01407_),
    .y(_01901_)
  );
  al_nor3fft _06994_ (
    .a(RESET),
    .b(_01899_),
    .c(_01901_),
    .y(\DFF_608.D )
  );
  al_or2 _06995_ (
    .a(TM1),
    .b(\DFF_865.Q ),
    .y(_01902_)
  );
  al_nand2 _06996_ (
    .a(TM1),
    .b(\DFF_865.Q ),
    .y(_01903_)
  );
  al_nand3 _06997_ (
    .a(\DFF_897.Q ),
    .b(_01902_),
    .c(_01903_),
    .y(_01904_)
  );
  al_nand2ft _06998_ (
    .a(TM1),
    .b(\DFF_865.Q ),
    .y(_01905_)
  );
  al_and2ft _06999_ (
    .a(\DFF_865.Q ),
    .b(TM1),
    .y(_01906_)
  );
  al_and3fft _07000_ (
    .a(\DFF_897.Q ),
    .b(_01906_),
    .c(_01905_),
    .y(_01907_)
  );
  al_and2ft _07001_ (
    .a(\DFF_833.Q ),
    .b(\DFF_801.Q ),
    .y(_01908_)
  );
  al_nand2ft _07002_ (
    .a(\DFF_801.Q ),
    .b(\DFF_833.Q ),
    .y(_01909_)
  );
  al_nand2ft _07003_ (
    .a(_01908_),
    .b(_01909_),
    .y(_01910_)
  );
  al_oai21ftf _07004_ (
    .a(_01904_),
    .b(_01907_),
    .c(_01910_),
    .y(_01911_)
  );
  al_nand3ftt _07005_ (
    .a(_01907_),
    .b(_01904_),
    .c(_01910_),
    .y(_01912_)
  );
  al_nand3 _07006_ (
    .a(_00448_),
    .b(_01911_),
    .c(_01912_),
    .y(_01913_)
  );
  al_aoi21 _07007_ (
    .a(TM0),
    .b(\DFF_766.Q ),
    .c(TM1),
    .y(_01914_)
  );
  al_nand2 _07008_ (
    .a(_01914_),
    .b(_01913_),
    .y(_01915_)
  );
  al_aoi21ttf _07009_ (
    .a(TM0),
    .b(\DFF_577.Q ),
    .c(TM1),
    .y(_01916_)
  );
  al_and2 _07010_ (
    .a(_01916_),
    .b(_01423_),
    .y(_01917_)
  );
  al_nor3fft _07011_ (
    .a(RESET),
    .b(_01915_),
    .c(_01917_),
    .y(\DFF_609.D )
  );
  al_or2 _07012_ (
    .a(TM1),
    .b(\DFF_866.Q ),
    .y(_01918_)
  );
  al_nand2 _07013_ (
    .a(TM1),
    .b(\DFF_866.Q ),
    .y(_01919_)
  );
  al_nand3 _07014_ (
    .a(\DFF_898.Q ),
    .b(_01918_),
    .c(_01919_),
    .y(_01920_)
  );
  al_nand2ft _07015_ (
    .a(TM1),
    .b(\DFF_866.Q ),
    .y(_01921_)
  );
  al_and2ft _07016_ (
    .a(\DFF_866.Q ),
    .b(TM1),
    .y(_01922_)
  );
  al_and3fft _07017_ (
    .a(\DFF_898.Q ),
    .b(_01922_),
    .c(_01921_),
    .y(_01923_)
  );
  al_and2ft _07018_ (
    .a(\DFF_834.Q ),
    .b(\DFF_802.Q ),
    .y(_01924_)
  );
  al_nand2ft _07019_ (
    .a(\DFF_802.Q ),
    .b(\DFF_834.Q ),
    .y(_01925_)
  );
  al_nand2ft _07020_ (
    .a(_01924_),
    .b(_01925_),
    .y(_01926_)
  );
  al_oai21ftf _07021_ (
    .a(_01920_),
    .b(_01923_),
    .c(_01926_),
    .y(_01927_)
  );
  al_nand3ftt _07022_ (
    .a(_01923_),
    .b(_01920_),
    .c(_01926_),
    .y(_01928_)
  );
  al_nand3 _07023_ (
    .a(_00448_),
    .b(_01927_),
    .c(_01928_),
    .y(_01929_)
  );
  al_aoi21 _07024_ (
    .a(TM0),
    .b(\DFF_765.Q ),
    .c(TM1),
    .y(_01930_)
  );
  al_nand2 _07025_ (
    .a(_01930_),
    .b(_01929_),
    .y(_01931_)
  );
  al_aoi21ttf _07026_ (
    .a(TM0),
    .b(\DFF_578.Q ),
    .c(TM1),
    .y(_01932_)
  );
  al_and2 _07027_ (
    .a(_01932_),
    .b(_01439_),
    .y(_01933_)
  );
  al_nor3fft _07028_ (
    .a(RESET),
    .b(_01931_),
    .c(_01933_),
    .y(\DFF_610.D )
  );
  al_or2 _07029_ (
    .a(TM1),
    .b(\DFF_867.Q ),
    .y(_01934_)
  );
  al_nand2 _07030_ (
    .a(TM1),
    .b(\DFF_867.Q ),
    .y(_01935_)
  );
  al_nand3 _07031_ (
    .a(\DFF_899.Q ),
    .b(_01934_),
    .c(_01935_),
    .y(_01936_)
  );
  al_nand2ft _07032_ (
    .a(TM1),
    .b(\DFF_867.Q ),
    .y(_01937_)
  );
  al_and2ft _07033_ (
    .a(\DFF_867.Q ),
    .b(TM1),
    .y(_01938_)
  );
  al_and3fft _07034_ (
    .a(\DFF_899.Q ),
    .b(_01938_),
    .c(_01937_),
    .y(_01939_)
  );
  al_and2ft _07035_ (
    .a(\DFF_835.Q ),
    .b(\DFF_803.Q ),
    .y(_01940_)
  );
  al_nand2ft _07036_ (
    .a(\DFF_803.Q ),
    .b(\DFF_835.Q ),
    .y(_01941_)
  );
  al_nand2ft _07037_ (
    .a(_01940_),
    .b(_01941_),
    .y(_01942_)
  );
  al_oai21ftf _07038_ (
    .a(_01936_),
    .b(_01939_),
    .c(_01942_),
    .y(_01943_)
  );
  al_nand3ftt _07039_ (
    .a(_01939_),
    .b(_01936_),
    .c(_01942_),
    .y(_01944_)
  );
  al_nand3 _07040_ (
    .a(_00448_),
    .b(_01943_),
    .c(_01944_),
    .y(_01945_)
  );
  al_aoi21 _07041_ (
    .a(TM0),
    .b(\DFF_764.Q ),
    .c(TM1),
    .y(_01946_)
  );
  al_nand2 _07042_ (
    .a(_01946_),
    .b(_01945_),
    .y(_01947_)
  );
  al_aoi21ttf _07043_ (
    .a(TM0),
    .b(\DFF_579.Q ),
    .c(TM1),
    .y(_01948_)
  );
  al_and2 _07044_ (
    .a(_01948_),
    .b(_01455_),
    .y(_01949_)
  );
  al_nor3fft _07045_ (
    .a(RESET),
    .b(_01947_),
    .c(_01949_),
    .y(\DFF_611.D )
  );
  al_or2 _07046_ (
    .a(TM1),
    .b(\DFF_868.Q ),
    .y(_01950_)
  );
  al_nand2 _07047_ (
    .a(TM1),
    .b(\DFF_868.Q ),
    .y(_01951_)
  );
  al_nand3 _07048_ (
    .a(\DFF_900.Q ),
    .b(_01950_),
    .c(_01951_),
    .y(_01952_)
  );
  al_nand2ft _07049_ (
    .a(TM1),
    .b(\DFF_868.Q ),
    .y(_01953_)
  );
  al_and2ft _07050_ (
    .a(\DFF_868.Q ),
    .b(TM1),
    .y(_01954_)
  );
  al_and3fft _07051_ (
    .a(\DFF_900.Q ),
    .b(_01954_),
    .c(_01953_),
    .y(_01955_)
  );
  al_and2ft _07052_ (
    .a(\DFF_836.Q ),
    .b(\DFF_804.Q ),
    .y(_01956_)
  );
  al_nand2ft _07053_ (
    .a(\DFF_804.Q ),
    .b(\DFF_836.Q ),
    .y(_01957_)
  );
  al_nand2ft _07054_ (
    .a(_01956_),
    .b(_01957_),
    .y(_01958_)
  );
  al_oai21ftf _07055_ (
    .a(_01952_),
    .b(_01955_),
    .c(_01958_),
    .y(_01959_)
  );
  al_nand3ftt _07056_ (
    .a(_01955_),
    .b(_01952_),
    .c(_01958_),
    .y(_01960_)
  );
  al_nand3 _07057_ (
    .a(_00448_),
    .b(_01959_),
    .c(_01960_),
    .y(_01961_)
  );
  al_aoi21 _07058_ (
    .a(TM0),
    .b(\DFF_763.Q ),
    .c(TM1),
    .y(_01962_)
  );
  al_nand2 _07059_ (
    .a(_01962_),
    .b(_01961_),
    .y(_01963_)
  );
  al_aoi21ttf _07060_ (
    .a(TM0),
    .b(\DFF_580.Q ),
    .c(TM1),
    .y(_01964_)
  );
  al_and2 _07061_ (
    .a(_01964_),
    .b(_01471_),
    .y(_01965_)
  );
  al_nor3fft _07062_ (
    .a(RESET),
    .b(_01963_),
    .c(_01965_),
    .y(\DFF_612.D )
  );
  al_or2 _07063_ (
    .a(TM1),
    .b(\DFF_869.Q ),
    .y(_01966_)
  );
  al_nand2 _07064_ (
    .a(TM1),
    .b(\DFF_869.Q ),
    .y(_01967_)
  );
  al_nand3 _07065_ (
    .a(\DFF_901.Q ),
    .b(_01966_),
    .c(_01967_),
    .y(_01968_)
  );
  al_nand2ft _07066_ (
    .a(TM1),
    .b(\DFF_869.Q ),
    .y(_01969_)
  );
  al_and2ft _07067_ (
    .a(\DFF_869.Q ),
    .b(TM1),
    .y(_01970_)
  );
  al_and3fft _07068_ (
    .a(\DFF_901.Q ),
    .b(_01970_),
    .c(_01969_),
    .y(_01971_)
  );
  al_and2ft _07069_ (
    .a(\DFF_837.Q ),
    .b(\DFF_805.Q ),
    .y(_01972_)
  );
  al_nand2ft _07070_ (
    .a(\DFF_805.Q ),
    .b(\DFF_837.Q ),
    .y(_01973_)
  );
  al_nand2ft _07071_ (
    .a(_01972_),
    .b(_01973_),
    .y(_01974_)
  );
  al_oai21ftf _07072_ (
    .a(_01968_),
    .b(_01971_),
    .c(_01974_),
    .y(_01975_)
  );
  al_nand3ftt _07073_ (
    .a(_01971_),
    .b(_01968_),
    .c(_01974_),
    .y(_01976_)
  );
  al_nand3 _07074_ (
    .a(_00448_),
    .b(_01975_),
    .c(_01976_),
    .y(_01977_)
  );
  al_aoi21 _07075_ (
    .a(TM0),
    .b(\DFF_762.Q ),
    .c(TM1),
    .y(_01978_)
  );
  al_nand2 _07076_ (
    .a(_01978_),
    .b(_01977_),
    .y(_01979_)
  );
  al_aoi21ttf _07077_ (
    .a(TM0),
    .b(\DFF_581.Q ),
    .c(TM1),
    .y(_01980_)
  );
  al_and2 _07078_ (
    .a(_01980_),
    .b(_01487_),
    .y(_01981_)
  );
  al_nor3fft _07079_ (
    .a(RESET),
    .b(_01979_),
    .c(_01981_),
    .y(\DFF_613.D )
  );
  al_or2 _07080_ (
    .a(TM1),
    .b(\DFF_870.Q ),
    .y(_01982_)
  );
  al_nand2 _07081_ (
    .a(TM1),
    .b(\DFF_870.Q ),
    .y(_01983_)
  );
  al_nand3 _07082_ (
    .a(\DFF_902.Q ),
    .b(_01982_),
    .c(_01983_),
    .y(_01984_)
  );
  al_nand2ft _07083_ (
    .a(TM1),
    .b(\DFF_870.Q ),
    .y(_01985_)
  );
  al_and2ft _07084_ (
    .a(\DFF_870.Q ),
    .b(TM1),
    .y(_01986_)
  );
  al_and3fft _07085_ (
    .a(\DFF_902.Q ),
    .b(_01986_),
    .c(_01985_),
    .y(_01987_)
  );
  al_and2ft _07086_ (
    .a(\DFF_838.Q ),
    .b(\DFF_806.Q ),
    .y(_01988_)
  );
  al_nand2ft _07087_ (
    .a(\DFF_806.Q ),
    .b(\DFF_838.Q ),
    .y(_01989_)
  );
  al_nand2ft _07088_ (
    .a(_01988_),
    .b(_01989_),
    .y(_01990_)
  );
  al_oai21ftf _07089_ (
    .a(_01984_),
    .b(_01987_),
    .c(_01990_),
    .y(_01991_)
  );
  al_nand3ftt _07090_ (
    .a(_01987_),
    .b(_01984_),
    .c(_01990_),
    .y(_01992_)
  );
  al_nand3 _07091_ (
    .a(_00448_),
    .b(_01991_),
    .c(_01992_),
    .y(_01993_)
  );
  al_aoi21 _07092_ (
    .a(TM0),
    .b(\DFF_761.Q ),
    .c(TM1),
    .y(_01994_)
  );
  al_nand2 _07093_ (
    .a(_01994_),
    .b(_01993_),
    .y(_01995_)
  );
  al_aoi21ttf _07094_ (
    .a(TM0),
    .b(\DFF_582.Q ),
    .c(TM1),
    .y(_01996_)
  );
  al_and2 _07095_ (
    .a(_01996_),
    .b(_01503_),
    .y(_01997_)
  );
  al_nor3fft _07096_ (
    .a(RESET),
    .b(_01995_),
    .c(_01997_),
    .y(\DFF_614.D )
  );
  al_or2 _07097_ (
    .a(TM1),
    .b(\DFF_871.Q ),
    .y(_01998_)
  );
  al_nand2 _07098_ (
    .a(TM1),
    .b(\DFF_871.Q ),
    .y(_01999_)
  );
  al_nand3 _07099_ (
    .a(\DFF_903.Q ),
    .b(_01998_),
    .c(_01999_),
    .y(_02000_)
  );
  al_nand2ft _07100_ (
    .a(TM1),
    .b(\DFF_871.Q ),
    .y(_02001_)
  );
  al_and2ft _07101_ (
    .a(\DFF_871.Q ),
    .b(TM1),
    .y(_02002_)
  );
  al_and3fft _07102_ (
    .a(\DFF_903.Q ),
    .b(_02002_),
    .c(_02001_),
    .y(_02003_)
  );
  al_and2ft _07103_ (
    .a(\DFF_839.Q ),
    .b(\DFF_807.Q ),
    .y(_02004_)
  );
  al_nand2ft _07104_ (
    .a(\DFF_807.Q ),
    .b(\DFF_839.Q ),
    .y(_02005_)
  );
  al_nand2ft _07105_ (
    .a(_02004_),
    .b(_02005_),
    .y(_02006_)
  );
  al_oai21ftf _07106_ (
    .a(_02000_),
    .b(_02003_),
    .c(_02006_),
    .y(_02007_)
  );
  al_nand3ftt _07107_ (
    .a(_02003_),
    .b(_02000_),
    .c(_02006_),
    .y(_02008_)
  );
  al_nand3 _07108_ (
    .a(_00448_),
    .b(_02007_),
    .c(_02008_),
    .y(_02009_)
  );
  al_aoi21 _07109_ (
    .a(TM0),
    .b(\DFF_760.Q ),
    .c(TM1),
    .y(_02010_)
  );
  al_nand2 _07110_ (
    .a(_02010_),
    .b(_02009_),
    .y(_02011_)
  );
  al_aoi21ttf _07111_ (
    .a(TM0),
    .b(\DFF_583.Q ),
    .c(TM1),
    .y(_02012_)
  );
  al_and2 _07112_ (
    .a(_02012_),
    .b(_01519_),
    .y(_02013_)
  );
  al_nor3fft _07113_ (
    .a(RESET),
    .b(_02011_),
    .c(_02013_),
    .y(\DFF_615.D )
  );
  al_or2 _07114_ (
    .a(TM1),
    .b(\DFF_872.Q ),
    .y(_02014_)
  );
  al_nand2 _07115_ (
    .a(TM1),
    .b(\DFF_872.Q ),
    .y(_02015_)
  );
  al_nand3 _07116_ (
    .a(\DFF_904.Q ),
    .b(_02014_),
    .c(_02015_),
    .y(_02016_)
  );
  al_nand2ft _07117_ (
    .a(TM1),
    .b(\DFF_872.Q ),
    .y(_02017_)
  );
  al_and2ft _07118_ (
    .a(\DFF_872.Q ),
    .b(TM1),
    .y(_02018_)
  );
  al_and3fft _07119_ (
    .a(\DFF_904.Q ),
    .b(_02018_),
    .c(_02017_),
    .y(_02019_)
  );
  al_and2ft _07120_ (
    .a(\DFF_840.Q ),
    .b(\DFF_808.Q ),
    .y(_02020_)
  );
  al_nand2ft _07121_ (
    .a(\DFF_808.Q ),
    .b(\DFF_840.Q ),
    .y(_02021_)
  );
  al_nand2ft _07122_ (
    .a(_02020_),
    .b(_02021_),
    .y(_02022_)
  );
  al_oai21ftf _07123_ (
    .a(_02016_),
    .b(_02019_),
    .c(_02022_),
    .y(_02023_)
  );
  al_nand3ftt _07124_ (
    .a(_02019_),
    .b(_02016_),
    .c(_02022_),
    .y(_02024_)
  );
  al_nand3 _07125_ (
    .a(_00448_),
    .b(_02023_),
    .c(_02024_),
    .y(_02025_)
  );
  al_aoi21 _07126_ (
    .a(TM0),
    .b(\DFF_759.Q ),
    .c(TM1),
    .y(_02026_)
  );
  al_nand2 _07127_ (
    .a(_02026_),
    .b(_02025_),
    .y(_02027_)
  );
  al_aoi21ttf _07128_ (
    .a(TM0),
    .b(\DFF_584.Q ),
    .c(TM1),
    .y(_02028_)
  );
  al_and2 _07129_ (
    .a(_02028_),
    .b(_01535_),
    .y(_02029_)
  );
  al_nor3fft _07130_ (
    .a(RESET),
    .b(_02027_),
    .c(_02029_),
    .y(\DFF_616.D )
  );
  al_or2 _07131_ (
    .a(TM1),
    .b(\DFF_873.Q ),
    .y(_02030_)
  );
  al_nand2 _07132_ (
    .a(TM1),
    .b(\DFF_873.Q ),
    .y(_02031_)
  );
  al_nand3 _07133_ (
    .a(\DFF_905.Q ),
    .b(_02030_),
    .c(_02031_),
    .y(_02032_)
  );
  al_nand2ft _07134_ (
    .a(TM1),
    .b(\DFF_873.Q ),
    .y(_02033_)
  );
  al_and2ft _07135_ (
    .a(\DFF_873.Q ),
    .b(TM1),
    .y(_02034_)
  );
  al_and3fft _07136_ (
    .a(\DFF_905.Q ),
    .b(_02034_),
    .c(_02033_),
    .y(_02035_)
  );
  al_and2ft _07137_ (
    .a(\DFF_841.Q ),
    .b(\DFF_809.Q ),
    .y(_02036_)
  );
  al_nand2ft _07138_ (
    .a(\DFF_809.Q ),
    .b(\DFF_841.Q ),
    .y(_02037_)
  );
  al_nand2ft _07139_ (
    .a(_02036_),
    .b(_02037_),
    .y(_02038_)
  );
  al_oai21ftf _07140_ (
    .a(_02032_),
    .b(_02035_),
    .c(_02038_),
    .y(_02039_)
  );
  al_nand3ftt _07141_ (
    .a(_02035_),
    .b(_02032_),
    .c(_02038_),
    .y(_02040_)
  );
  al_nand3 _07142_ (
    .a(_00448_),
    .b(_02039_),
    .c(_02040_),
    .y(_02041_)
  );
  al_aoi21 _07143_ (
    .a(TM0),
    .b(\DFF_758.Q ),
    .c(TM1),
    .y(_02042_)
  );
  al_nand2 _07144_ (
    .a(_02042_),
    .b(_02041_),
    .y(_02043_)
  );
  al_aoi21ttf _07145_ (
    .a(TM0),
    .b(\DFF_585.Q ),
    .c(TM1),
    .y(_02044_)
  );
  al_and2 _07146_ (
    .a(_02044_),
    .b(_01551_),
    .y(_02045_)
  );
  al_nor3fft _07147_ (
    .a(RESET),
    .b(_02043_),
    .c(_02045_),
    .y(\DFF_617.D )
  );
  al_or2 _07148_ (
    .a(TM1),
    .b(\DFF_874.Q ),
    .y(_02046_)
  );
  al_nand2 _07149_ (
    .a(TM1),
    .b(\DFF_874.Q ),
    .y(_02047_)
  );
  al_nand3 _07150_ (
    .a(\DFF_906.Q ),
    .b(_02046_),
    .c(_02047_),
    .y(_02048_)
  );
  al_nand2ft _07151_ (
    .a(TM1),
    .b(\DFF_874.Q ),
    .y(_02049_)
  );
  al_and2ft _07152_ (
    .a(\DFF_874.Q ),
    .b(TM1),
    .y(_02050_)
  );
  al_and3fft _07153_ (
    .a(\DFF_906.Q ),
    .b(_02050_),
    .c(_02049_),
    .y(_02051_)
  );
  al_and2ft _07154_ (
    .a(\DFF_842.Q ),
    .b(\DFF_810.Q ),
    .y(_02052_)
  );
  al_nand2ft _07155_ (
    .a(\DFF_810.Q ),
    .b(\DFF_842.Q ),
    .y(_02053_)
  );
  al_nand2ft _07156_ (
    .a(_02052_),
    .b(_02053_),
    .y(_02054_)
  );
  al_oai21ftf _07157_ (
    .a(_02048_),
    .b(_02051_),
    .c(_02054_),
    .y(_02055_)
  );
  al_nand3ftt _07158_ (
    .a(_02051_),
    .b(_02048_),
    .c(_02054_),
    .y(_02056_)
  );
  al_nand3 _07159_ (
    .a(_00448_),
    .b(_02055_),
    .c(_02056_),
    .y(_02057_)
  );
  al_aoi21 _07160_ (
    .a(TM0),
    .b(\DFF_757.Q ),
    .c(TM1),
    .y(_02058_)
  );
  al_nand2 _07161_ (
    .a(_02058_),
    .b(_02057_),
    .y(_02059_)
  );
  al_aoi21ttf _07162_ (
    .a(TM0),
    .b(\DFF_586.Q ),
    .c(TM1),
    .y(_02060_)
  );
  al_and2 _07163_ (
    .a(_02060_),
    .b(_01567_),
    .y(_02061_)
  );
  al_nor3fft _07164_ (
    .a(RESET),
    .b(_02059_),
    .c(_02061_),
    .y(\DFF_618.D )
  );
  al_or2 _07165_ (
    .a(TM1),
    .b(\DFF_875.Q ),
    .y(_02062_)
  );
  al_nand2 _07166_ (
    .a(TM1),
    .b(\DFF_875.Q ),
    .y(_02063_)
  );
  al_nand3 _07167_ (
    .a(\DFF_907.Q ),
    .b(_02062_),
    .c(_02063_),
    .y(_02064_)
  );
  al_nand2ft _07168_ (
    .a(TM1),
    .b(\DFF_875.Q ),
    .y(_02065_)
  );
  al_and2ft _07169_ (
    .a(\DFF_875.Q ),
    .b(TM1),
    .y(_02066_)
  );
  al_and3fft _07170_ (
    .a(\DFF_907.Q ),
    .b(_02066_),
    .c(_02065_),
    .y(_02067_)
  );
  al_and2ft _07171_ (
    .a(\DFF_843.Q ),
    .b(\DFF_811.Q ),
    .y(_02068_)
  );
  al_nand2ft _07172_ (
    .a(\DFF_811.Q ),
    .b(\DFF_843.Q ),
    .y(_02069_)
  );
  al_nand2ft _07173_ (
    .a(_02068_),
    .b(_02069_),
    .y(_02070_)
  );
  al_oai21ftf _07174_ (
    .a(_02064_),
    .b(_02067_),
    .c(_02070_),
    .y(_02071_)
  );
  al_nand3ftt _07175_ (
    .a(_02067_),
    .b(_02064_),
    .c(_02070_),
    .y(_02072_)
  );
  al_nand3 _07176_ (
    .a(_00448_),
    .b(_02071_),
    .c(_02072_),
    .y(_02073_)
  );
  al_aoi21 _07177_ (
    .a(TM0),
    .b(\DFF_756.Q ),
    .c(TM1),
    .y(_02074_)
  );
  al_nand2 _07178_ (
    .a(_02074_),
    .b(_02073_),
    .y(_02075_)
  );
  al_aoi21ttf _07179_ (
    .a(TM0),
    .b(\DFF_587.Q ),
    .c(TM1),
    .y(_02076_)
  );
  al_and2 _07180_ (
    .a(_02076_),
    .b(_01583_),
    .y(_02077_)
  );
  al_nor3fft _07181_ (
    .a(RESET),
    .b(_02075_),
    .c(_02077_),
    .y(\DFF_619.D )
  );
  al_or2 _07182_ (
    .a(TM1),
    .b(\DFF_876.Q ),
    .y(_02078_)
  );
  al_nand2 _07183_ (
    .a(TM1),
    .b(\DFF_876.Q ),
    .y(_02079_)
  );
  al_nand3 _07184_ (
    .a(\DFF_908.Q ),
    .b(_02078_),
    .c(_02079_),
    .y(_02080_)
  );
  al_nand2ft _07185_ (
    .a(TM1),
    .b(\DFF_876.Q ),
    .y(_02081_)
  );
  al_and2ft _07186_ (
    .a(\DFF_876.Q ),
    .b(TM1),
    .y(_02082_)
  );
  al_and3fft _07187_ (
    .a(\DFF_908.Q ),
    .b(_02082_),
    .c(_02081_),
    .y(_02083_)
  );
  al_and2ft _07188_ (
    .a(\DFF_844.Q ),
    .b(\DFF_812.Q ),
    .y(_02084_)
  );
  al_nand2ft _07189_ (
    .a(\DFF_812.Q ),
    .b(\DFF_844.Q ),
    .y(_02085_)
  );
  al_nand2ft _07190_ (
    .a(_02084_),
    .b(_02085_),
    .y(_02086_)
  );
  al_oai21ftf _07191_ (
    .a(_02080_),
    .b(_02083_),
    .c(_02086_),
    .y(_02087_)
  );
  al_nand3ftt _07192_ (
    .a(_02083_),
    .b(_02080_),
    .c(_02086_),
    .y(_02088_)
  );
  al_nand3 _07193_ (
    .a(_00448_),
    .b(_02087_),
    .c(_02088_),
    .y(_02089_)
  );
  al_aoi21 _07194_ (
    .a(TM0),
    .b(\DFF_755.Q ),
    .c(TM1),
    .y(_02090_)
  );
  al_nand2 _07195_ (
    .a(_02090_),
    .b(_02089_),
    .y(_02091_)
  );
  al_aoi21ttf _07196_ (
    .a(TM0),
    .b(\DFF_588.Q ),
    .c(TM1),
    .y(_02092_)
  );
  al_and2 _07197_ (
    .a(_02092_),
    .b(_01599_),
    .y(_02093_)
  );
  al_nor3fft _07198_ (
    .a(RESET),
    .b(_02091_),
    .c(_02093_),
    .y(\DFF_620.D )
  );
  al_or2 _07199_ (
    .a(TM1),
    .b(\DFF_877.Q ),
    .y(_02094_)
  );
  al_nand2 _07200_ (
    .a(TM1),
    .b(\DFF_877.Q ),
    .y(_02095_)
  );
  al_nand3 _07201_ (
    .a(\DFF_909.Q ),
    .b(_02094_),
    .c(_02095_),
    .y(_02096_)
  );
  al_nand2ft _07202_ (
    .a(TM1),
    .b(\DFF_877.Q ),
    .y(_02097_)
  );
  al_and2ft _07203_ (
    .a(\DFF_877.Q ),
    .b(TM1),
    .y(_02098_)
  );
  al_and3fft _07204_ (
    .a(\DFF_909.Q ),
    .b(_02098_),
    .c(_02097_),
    .y(_02099_)
  );
  al_and2ft _07205_ (
    .a(\DFF_845.Q ),
    .b(\DFF_813.Q ),
    .y(_02100_)
  );
  al_nand2ft _07206_ (
    .a(\DFF_813.Q ),
    .b(\DFF_845.Q ),
    .y(_02101_)
  );
  al_nand2ft _07207_ (
    .a(_02100_),
    .b(_02101_),
    .y(_02102_)
  );
  al_oai21ftf _07208_ (
    .a(_02096_),
    .b(_02099_),
    .c(_02102_),
    .y(_02103_)
  );
  al_nand3ftt _07209_ (
    .a(_02099_),
    .b(_02096_),
    .c(_02102_),
    .y(_02104_)
  );
  al_nand3 _07210_ (
    .a(_00448_),
    .b(_02103_),
    .c(_02104_),
    .y(_02105_)
  );
  al_aoi21 _07211_ (
    .a(TM0),
    .b(\DFF_754.Q ),
    .c(TM1),
    .y(_02106_)
  );
  al_nand2 _07212_ (
    .a(_02106_),
    .b(_02105_),
    .y(_02107_)
  );
  al_aoi21ttf _07213_ (
    .a(TM0),
    .b(\DFF_589.Q ),
    .c(TM1),
    .y(_02108_)
  );
  al_and2 _07214_ (
    .a(_02108_),
    .b(_01615_),
    .y(_02109_)
  );
  al_nor3fft _07215_ (
    .a(RESET),
    .b(_02107_),
    .c(_02109_),
    .y(\DFF_621.D )
  );
  al_or2 _07216_ (
    .a(TM1),
    .b(\DFF_878.Q ),
    .y(_02110_)
  );
  al_nand2 _07217_ (
    .a(TM1),
    .b(\DFF_878.Q ),
    .y(_02111_)
  );
  al_nand3 _07218_ (
    .a(\DFF_910.Q ),
    .b(_02110_),
    .c(_02111_),
    .y(_02112_)
  );
  al_nand2ft _07219_ (
    .a(TM1),
    .b(\DFF_878.Q ),
    .y(_02113_)
  );
  al_and2ft _07220_ (
    .a(\DFF_878.Q ),
    .b(TM1),
    .y(_02114_)
  );
  al_and3fft _07221_ (
    .a(\DFF_910.Q ),
    .b(_02114_),
    .c(_02113_),
    .y(_02115_)
  );
  al_and2ft _07222_ (
    .a(\DFF_846.Q ),
    .b(\DFF_814.Q ),
    .y(_02116_)
  );
  al_nand2ft _07223_ (
    .a(\DFF_814.Q ),
    .b(\DFF_846.Q ),
    .y(_02117_)
  );
  al_nand2ft _07224_ (
    .a(_02116_),
    .b(_02117_),
    .y(_02118_)
  );
  al_oai21ftf _07225_ (
    .a(_02112_),
    .b(_02115_),
    .c(_02118_),
    .y(_02119_)
  );
  al_nand3ftt _07226_ (
    .a(_02115_),
    .b(_02112_),
    .c(_02118_),
    .y(_02120_)
  );
  al_nand3 _07227_ (
    .a(_00448_),
    .b(_02119_),
    .c(_02120_),
    .y(_02121_)
  );
  al_aoi21 _07228_ (
    .a(TM0),
    .b(\DFF_753.Q ),
    .c(TM1),
    .y(_02122_)
  );
  al_nand2 _07229_ (
    .a(_02122_),
    .b(_02121_),
    .y(_02123_)
  );
  al_aoi21ttf _07230_ (
    .a(TM0),
    .b(\DFF_590.Q ),
    .c(TM1),
    .y(_02124_)
  );
  al_and2 _07231_ (
    .a(_02124_),
    .b(_01631_),
    .y(_02125_)
  );
  al_nor3fft _07232_ (
    .a(RESET),
    .b(_02123_),
    .c(_02125_),
    .y(\DFF_622.D )
  );
  al_or2 _07233_ (
    .a(TM1),
    .b(\DFF_879.Q ),
    .y(_02126_)
  );
  al_nand2 _07234_ (
    .a(TM1),
    .b(\DFF_879.Q ),
    .y(_02127_)
  );
  al_nand3 _07235_ (
    .a(\DFF_911.Q ),
    .b(_02126_),
    .c(_02127_),
    .y(_02128_)
  );
  al_nand2ft _07236_ (
    .a(TM1),
    .b(\DFF_879.Q ),
    .y(_02129_)
  );
  al_and2ft _07237_ (
    .a(\DFF_879.Q ),
    .b(TM1),
    .y(_02130_)
  );
  al_and3fft _07238_ (
    .a(\DFF_911.Q ),
    .b(_02130_),
    .c(_02129_),
    .y(_02131_)
  );
  al_and2ft _07239_ (
    .a(\DFF_847.Q ),
    .b(\DFF_815.Q ),
    .y(_02132_)
  );
  al_nand2ft _07240_ (
    .a(\DFF_815.Q ),
    .b(\DFF_847.Q ),
    .y(_02133_)
  );
  al_nand2ft _07241_ (
    .a(_02132_),
    .b(_02133_),
    .y(_02134_)
  );
  al_oai21ftf _07242_ (
    .a(_02128_),
    .b(_02131_),
    .c(_02134_),
    .y(_02135_)
  );
  al_nand3ftt _07243_ (
    .a(_02131_),
    .b(_02128_),
    .c(_02134_),
    .y(_02136_)
  );
  al_nand3 _07244_ (
    .a(_00448_),
    .b(_02135_),
    .c(_02136_),
    .y(_02137_)
  );
  al_aoi21 _07245_ (
    .a(TM0),
    .b(\DFF_752.Q ),
    .c(TM1),
    .y(_02138_)
  );
  al_nand2 _07246_ (
    .a(_02138_),
    .b(_02137_),
    .y(_02139_)
  );
  al_aoi21ttf _07247_ (
    .a(TM0),
    .b(\DFF_591.Q ),
    .c(TM1),
    .y(_02140_)
  );
  al_and2 _07248_ (
    .a(_02140_),
    .b(_01647_),
    .y(_02141_)
  );
  al_nor3fft _07249_ (
    .a(RESET),
    .b(_02139_),
    .c(_02141_),
    .y(\DFF_623.D )
  );
  al_nor2 _07250_ (
    .a(\DFF_848.Q ),
    .b(\DFF_880.Q ),
    .y(_02142_)
  );
  al_and2 _07251_ (
    .a(\DFF_848.Q ),
    .b(\DFF_880.Q ),
    .y(_02143_)
  );
  al_and2ft _07252_ (
    .a(\DFF_816.Q ),
    .b(\DFF_912.Q ),
    .y(_02144_)
  );
  al_nand2ft _07253_ (
    .a(\DFF_912.Q ),
    .b(\DFF_816.Q ),
    .y(_02145_)
  );
  al_nand2ft _07254_ (
    .a(_02144_),
    .b(_02145_),
    .y(_02146_)
  );
  al_oa21ttf _07255_ (
    .a(_02142_),
    .b(_02143_),
    .c(_02146_),
    .y(_02147_)
  );
  al_nand3fft _07256_ (
    .a(_02142_),
    .b(_02143_),
    .c(_02146_),
    .y(_02148_)
  );
  al_and3fft _07257_ (
    .a(TM0),
    .b(_02147_),
    .c(_02148_),
    .y(_02149_)
  );
  al_nand2 _07258_ (
    .a(TM0),
    .b(\DFF_751.Q ),
    .y(_02150_)
  );
  al_or3fft _07259_ (
    .a(_01652_),
    .b(_02150_),
    .c(_02149_),
    .y(_02151_)
  );
  al_and2 _07260_ (
    .a(TM0),
    .b(\DFF_592.Q ),
    .y(_02152_)
  );
  al_and3fft _07261_ (
    .a(_02152_),
    .b(_01660_),
    .c(TM1),
    .y(_02153_)
  );
  al_nor3fft _07262_ (
    .a(RESET),
    .b(_02151_),
    .c(_02153_),
    .y(\DFF_624.D )
  );
  al_nor2 _07263_ (
    .a(\DFF_849.Q ),
    .b(\DFF_881.Q ),
    .y(_02154_)
  );
  al_and2 _07264_ (
    .a(\DFF_849.Q ),
    .b(\DFF_881.Q ),
    .y(_02155_)
  );
  al_and2ft _07265_ (
    .a(\DFF_817.Q ),
    .b(\DFF_913.Q ),
    .y(_02156_)
  );
  al_nand2ft _07266_ (
    .a(\DFF_913.Q ),
    .b(\DFF_817.Q ),
    .y(_02157_)
  );
  al_nand2ft _07267_ (
    .a(_02156_),
    .b(_02157_),
    .y(_02158_)
  );
  al_oa21ttf _07268_ (
    .a(_02154_),
    .b(_02155_),
    .c(_02158_),
    .y(_02159_)
  );
  al_nand3fft _07269_ (
    .a(_02154_),
    .b(_02155_),
    .c(_02158_),
    .y(_02160_)
  );
  al_and3fft _07270_ (
    .a(TM0),
    .b(_02159_),
    .c(_02160_),
    .y(_02161_)
  );
  al_nand2 _07271_ (
    .a(TM0),
    .b(\DFF_750.Q ),
    .y(_02162_)
  );
  al_or3fft _07272_ (
    .a(_01652_),
    .b(_02162_),
    .c(_02161_),
    .y(_02163_)
  );
  al_and2 _07273_ (
    .a(TM0),
    .b(\DFF_593.Q ),
    .y(_02164_)
  );
  al_and3fft _07274_ (
    .a(_02164_),
    .b(_01672_),
    .c(TM1),
    .y(_02165_)
  );
  al_nor3fft _07275_ (
    .a(RESET),
    .b(_02163_),
    .c(_02165_),
    .y(\DFF_625.D )
  );
  al_nor2 _07276_ (
    .a(\DFF_850.Q ),
    .b(\DFF_882.Q ),
    .y(_02166_)
  );
  al_and2 _07277_ (
    .a(\DFF_850.Q ),
    .b(\DFF_882.Q ),
    .y(_02167_)
  );
  al_and2ft _07278_ (
    .a(\DFF_818.Q ),
    .b(\DFF_914.Q ),
    .y(_02168_)
  );
  al_nand2ft _07279_ (
    .a(\DFF_914.Q ),
    .b(\DFF_818.Q ),
    .y(_02169_)
  );
  al_nand2ft _07280_ (
    .a(_02168_),
    .b(_02169_),
    .y(_02170_)
  );
  al_oa21ttf _07281_ (
    .a(_02166_),
    .b(_02167_),
    .c(_02170_),
    .y(_02171_)
  );
  al_nand3fft _07282_ (
    .a(_02166_),
    .b(_02167_),
    .c(_02170_),
    .y(_02172_)
  );
  al_and3fft _07283_ (
    .a(TM0),
    .b(_02171_),
    .c(_02172_),
    .y(_02173_)
  );
  al_nand2 _07284_ (
    .a(TM0),
    .b(\DFF_749.Q ),
    .y(_02174_)
  );
  al_or3fft _07285_ (
    .a(_01652_),
    .b(_02174_),
    .c(_02173_),
    .y(_02175_)
  );
  al_and2 _07286_ (
    .a(TM0),
    .b(\DFF_594.Q ),
    .y(_02176_)
  );
  al_and3fft _07287_ (
    .a(_02176_),
    .b(_01684_),
    .c(TM1),
    .y(_02177_)
  );
  al_nor3fft _07288_ (
    .a(RESET),
    .b(_02175_),
    .c(_02177_),
    .y(\DFF_626.D )
  );
  al_nor2 _07289_ (
    .a(\DFF_851.Q ),
    .b(\DFF_883.Q ),
    .y(_02178_)
  );
  al_and2 _07290_ (
    .a(\DFF_851.Q ),
    .b(\DFF_883.Q ),
    .y(_02179_)
  );
  al_and2ft _07291_ (
    .a(\DFF_819.Q ),
    .b(\DFF_915.Q ),
    .y(_02180_)
  );
  al_nand2ft _07292_ (
    .a(\DFF_915.Q ),
    .b(\DFF_819.Q ),
    .y(_02181_)
  );
  al_nand2ft _07293_ (
    .a(_02180_),
    .b(_02181_),
    .y(_02182_)
  );
  al_oa21ttf _07294_ (
    .a(_02178_),
    .b(_02179_),
    .c(_02182_),
    .y(_02183_)
  );
  al_nand3fft _07295_ (
    .a(_02178_),
    .b(_02179_),
    .c(_02182_),
    .y(_02184_)
  );
  al_and3fft _07296_ (
    .a(TM0),
    .b(_02183_),
    .c(_02184_),
    .y(_02185_)
  );
  al_nand2 _07297_ (
    .a(TM0),
    .b(\DFF_748.Q ),
    .y(_02186_)
  );
  al_or3fft _07298_ (
    .a(_01652_),
    .b(_02186_),
    .c(_02185_),
    .y(_02187_)
  );
  al_and2 _07299_ (
    .a(TM0),
    .b(\DFF_595.Q ),
    .y(_02188_)
  );
  al_and3fft _07300_ (
    .a(_02188_),
    .b(_01696_),
    .c(TM1),
    .y(_02189_)
  );
  al_nor3fft _07301_ (
    .a(RESET),
    .b(_02187_),
    .c(_02189_),
    .y(\DFF_627.D )
  );
  al_nor2 _07302_ (
    .a(\DFF_852.Q ),
    .b(\DFF_884.Q ),
    .y(_02190_)
  );
  al_and2 _07303_ (
    .a(\DFF_852.Q ),
    .b(\DFF_884.Q ),
    .y(_02191_)
  );
  al_and2ft _07304_ (
    .a(\DFF_820.Q ),
    .b(\DFF_916.Q ),
    .y(_02192_)
  );
  al_nand2ft _07305_ (
    .a(\DFF_916.Q ),
    .b(\DFF_820.Q ),
    .y(_02193_)
  );
  al_nand2ft _07306_ (
    .a(_02192_),
    .b(_02193_),
    .y(_02194_)
  );
  al_oa21ttf _07307_ (
    .a(_02190_),
    .b(_02191_),
    .c(_02194_),
    .y(_02195_)
  );
  al_nand3fft _07308_ (
    .a(_02190_),
    .b(_02191_),
    .c(_02194_),
    .y(_02196_)
  );
  al_and3fft _07309_ (
    .a(TM0),
    .b(_02195_),
    .c(_02196_),
    .y(_02197_)
  );
  al_nand2 _07310_ (
    .a(TM0),
    .b(\DFF_747.Q ),
    .y(_02198_)
  );
  al_or3fft _07311_ (
    .a(_01652_),
    .b(_02198_),
    .c(_02197_),
    .y(_02199_)
  );
  al_and2 _07312_ (
    .a(TM0),
    .b(\DFF_596.Q ),
    .y(_02200_)
  );
  al_and3fft _07313_ (
    .a(_02200_),
    .b(_01708_),
    .c(TM1),
    .y(_02201_)
  );
  al_nor3fft _07314_ (
    .a(RESET),
    .b(_02199_),
    .c(_02201_),
    .y(\DFF_628.D )
  );
  al_nor2 _07315_ (
    .a(\DFF_853.Q ),
    .b(\DFF_885.Q ),
    .y(_02202_)
  );
  al_and2 _07316_ (
    .a(\DFF_853.Q ),
    .b(\DFF_885.Q ),
    .y(_02203_)
  );
  al_and2ft _07317_ (
    .a(\DFF_821.Q ),
    .b(\DFF_917.Q ),
    .y(_02204_)
  );
  al_nand2ft _07318_ (
    .a(\DFF_917.Q ),
    .b(\DFF_821.Q ),
    .y(_02205_)
  );
  al_nand2ft _07319_ (
    .a(_02204_),
    .b(_02205_),
    .y(_02206_)
  );
  al_oa21ttf _07320_ (
    .a(_02202_),
    .b(_02203_),
    .c(_02206_),
    .y(_02207_)
  );
  al_nand3fft _07321_ (
    .a(_02202_),
    .b(_02203_),
    .c(_02206_),
    .y(_02208_)
  );
  al_and3fft _07322_ (
    .a(TM0),
    .b(_02207_),
    .c(_02208_),
    .y(_02209_)
  );
  al_nand2 _07323_ (
    .a(TM0),
    .b(\DFF_746.Q ),
    .y(_02210_)
  );
  al_or3fft _07324_ (
    .a(_01652_),
    .b(_02210_),
    .c(_02209_),
    .y(_02211_)
  );
  al_and2 _07325_ (
    .a(TM0),
    .b(\DFF_597.Q ),
    .y(_02212_)
  );
  al_and3fft _07326_ (
    .a(_02212_),
    .b(_01720_),
    .c(TM1),
    .y(_02213_)
  );
  al_nor3fft _07327_ (
    .a(RESET),
    .b(_02211_),
    .c(_02213_),
    .y(\DFF_629.D )
  );
  al_nor2 _07328_ (
    .a(\DFF_854.Q ),
    .b(\DFF_886.Q ),
    .y(_02214_)
  );
  al_and2 _07329_ (
    .a(\DFF_854.Q ),
    .b(\DFF_886.Q ),
    .y(_02215_)
  );
  al_and2ft _07330_ (
    .a(\DFF_822.Q ),
    .b(\DFF_918.Q ),
    .y(_02216_)
  );
  al_nand2ft _07331_ (
    .a(\DFF_918.Q ),
    .b(\DFF_822.Q ),
    .y(_02217_)
  );
  al_nand2ft _07332_ (
    .a(_02216_),
    .b(_02217_),
    .y(_02218_)
  );
  al_oa21ttf _07333_ (
    .a(_02214_),
    .b(_02215_),
    .c(_02218_),
    .y(_02219_)
  );
  al_nand3fft _07334_ (
    .a(_02214_),
    .b(_02215_),
    .c(_02218_),
    .y(_02220_)
  );
  al_and3fft _07335_ (
    .a(TM0),
    .b(_02219_),
    .c(_02220_),
    .y(_02221_)
  );
  al_nand2 _07336_ (
    .a(TM0),
    .b(\DFF_745.Q ),
    .y(_02222_)
  );
  al_or3fft _07337_ (
    .a(_01652_),
    .b(_02222_),
    .c(_02221_),
    .y(_02223_)
  );
  al_and2 _07338_ (
    .a(TM0),
    .b(\DFF_598.Q ),
    .y(_02224_)
  );
  al_and3fft _07339_ (
    .a(_02224_),
    .b(_01732_),
    .c(TM1),
    .y(_02225_)
  );
  al_nor3fft _07340_ (
    .a(RESET),
    .b(_02223_),
    .c(_02225_),
    .y(\DFF_630.D )
  );
  al_nor2 _07341_ (
    .a(\DFF_855.Q ),
    .b(\DFF_887.Q ),
    .y(_02226_)
  );
  al_and2 _07342_ (
    .a(\DFF_855.Q ),
    .b(\DFF_887.Q ),
    .y(_02227_)
  );
  al_and2ft _07343_ (
    .a(\DFF_823.Q ),
    .b(\DFF_919.Q ),
    .y(_02228_)
  );
  al_nand2ft _07344_ (
    .a(\DFF_919.Q ),
    .b(\DFF_823.Q ),
    .y(_02229_)
  );
  al_nand2ft _07345_ (
    .a(_02228_),
    .b(_02229_),
    .y(_02230_)
  );
  al_oa21ttf _07346_ (
    .a(_02226_),
    .b(_02227_),
    .c(_02230_),
    .y(_02231_)
  );
  al_nand3fft _07347_ (
    .a(_02226_),
    .b(_02227_),
    .c(_02230_),
    .y(_02232_)
  );
  al_and3fft _07348_ (
    .a(TM0),
    .b(_02231_),
    .c(_02232_),
    .y(_02233_)
  );
  al_nand2 _07349_ (
    .a(TM0),
    .b(\DFF_744.Q ),
    .y(_02234_)
  );
  al_or3fft _07350_ (
    .a(_01652_),
    .b(_02234_),
    .c(_02233_),
    .y(_02235_)
  );
  al_and2 _07351_ (
    .a(TM0),
    .b(\DFF_599.Q ),
    .y(_02236_)
  );
  al_and3fft _07352_ (
    .a(_02236_),
    .b(_01744_),
    .c(TM1),
    .y(_02237_)
  );
  al_nor3fft _07353_ (
    .a(RESET),
    .b(_02235_),
    .c(_02237_),
    .y(\DFF_631.D )
  );
  al_nor2 _07354_ (
    .a(\DFF_856.Q ),
    .b(\DFF_888.Q ),
    .y(_02238_)
  );
  al_and2 _07355_ (
    .a(\DFF_856.Q ),
    .b(\DFF_888.Q ),
    .y(_02239_)
  );
  al_and2ft _07356_ (
    .a(\DFF_824.Q ),
    .b(\DFF_920.Q ),
    .y(_02240_)
  );
  al_nand2ft _07357_ (
    .a(\DFF_920.Q ),
    .b(\DFF_824.Q ),
    .y(_02241_)
  );
  al_nand2ft _07358_ (
    .a(_02240_),
    .b(_02241_),
    .y(_02242_)
  );
  al_oa21ttf _07359_ (
    .a(_02238_),
    .b(_02239_),
    .c(_02242_),
    .y(_02243_)
  );
  al_nand3fft _07360_ (
    .a(_02238_),
    .b(_02239_),
    .c(_02242_),
    .y(_02244_)
  );
  al_and3fft _07361_ (
    .a(TM0),
    .b(_02243_),
    .c(_02244_),
    .y(_02245_)
  );
  al_nand2 _07362_ (
    .a(TM0),
    .b(\DFF_743.Q ),
    .y(_02246_)
  );
  al_or3fft _07363_ (
    .a(_01652_),
    .b(_02246_),
    .c(_02245_),
    .y(_02247_)
  );
  al_and2 _07364_ (
    .a(TM0),
    .b(\DFF_600.Q ),
    .y(_02248_)
  );
  al_and3fft _07365_ (
    .a(_02248_),
    .b(_01756_),
    .c(TM1),
    .y(_02249_)
  );
  al_nor3fft _07366_ (
    .a(RESET),
    .b(_02247_),
    .c(_02249_),
    .y(\DFF_632.D )
  );
  al_nor2 _07367_ (
    .a(\DFF_857.Q ),
    .b(\DFF_889.Q ),
    .y(_02250_)
  );
  al_and2 _07368_ (
    .a(\DFF_857.Q ),
    .b(\DFF_889.Q ),
    .y(_02251_)
  );
  al_and2ft _07369_ (
    .a(\DFF_825.Q ),
    .b(\DFF_921.Q ),
    .y(_02252_)
  );
  al_nand2ft _07370_ (
    .a(\DFF_921.Q ),
    .b(\DFF_825.Q ),
    .y(_02253_)
  );
  al_nand2ft _07371_ (
    .a(_02252_),
    .b(_02253_),
    .y(_02254_)
  );
  al_oa21ttf _07372_ (
    .a(_02250_),
    .b(_02251_),
    .c(_02254_),
    .y(_02255_)
  );
  al_nand3fft _07373_ (
    .a(_02250_),
    .b(_02251_),
    .c(_02254_),
    .y(_02256_)
  );
  al_and3fft _07374_ (
    .a(TM0),
    .b(_02255_),
    .c(_02256_),
    .y(_02257_)
  );
  al_nand2 _07375_ (
    .a(TM0),
    .b(\DFF_742.Q ),
    .y(_02258_)
  );
  al_or3fft _07376_ (
    .a(_01652_),
    .b(_02258_),
    .c(_02257_),
    .y(_02259_)
  );
  al_and2 _07377_ (
    .a(TM0),
    .b(\DFF_601.Q ),
    .y(_02260_)
  );
  al_and3fft _07378_ (
    .a(_02260_),
    .b(_01768_),
    .c(TM1),
    .y(_02261_)
  );
  al_nor3fft _07379_ (
    .a(RESET),
    .b(_02259_),
    .c(_02261_),
    .y(\DFF_633.D )
  );
  al_nor2 _07380_ (
    .a(\DFF_858.Q ),
    .b(\DFF_890.Q ),
    .y(_02262_)
  );
  al_and2 _07381_ (
    .a(\DFF_858.Q ),
    .b(\DFF_890.Q ),
    .y(_02263_)
  );
  al_and2ft _07382_ (
    .a(\DFF_826.Q ),
    .b(\DFF_922.Q ),
    .y(_02264_)
  );
  al_nand2ft _07383_ (
    .a(\DFF_922.Q ),
    .b(\DFF_826.Q ),
    .y(_02265_)
  );
  al_nand2ft _07384_ (
    .a(_02264_),
    .b(_02265_),
    .y(_02266_)
  );
  al_oa21ttf _07385_ (
    .a(_02262_),
    .b(_02263_),
    .c(_02266_),
    .y(_02267_)
  );
  al_nand3fft _07386_ (
    .a(_02262_),
    .b(_02263_),
    .c(_02266_),
    .y(_02268_)
  );
  al_and3fft _07387_ (
    .a(TM0),
    .b(_02267_),
    .c(_02268_),
    .y(_02269_)
  );
  al_nand2 _07388_ (
    .a(TM0),
    .b(\DFF_741.Q ),
    .y(_02270_)
  );
  al_or3fft _07389_ (
    .a(_01652_),
    .b(_02270_),
    .c(_02269_),
    .y(_02271_)
  );
  al_and2 _07390_ (
    .a(TM0),
    .b(\DFF_602.Q ),
    .y(_02272_)
  );
  al_and3fft _07391_ (
    .a(_02272_),
    .b(_01780_),
    .c(TM1),
    .y(_02273_)
  );
  al_nor3fft _07392_ (
    .a(RESET),
    .b(_02271_),
    .c(_02273_),
    .y(\DFF_634.D )
  );
  al_nor2 _07393_ (
    .a(\DFF_859.Q ),
    .b(\DFF_891.Q ),
    .y(_02274_)
  );
  al_and2 _07394_ (
    .a(\DFF_859.Q ),
    .b(\DFF_891.Q ),
    .y(_02275_)
  );
  al_and2ft _07395_ (
    .a(\DFF_827.Q ),
    .b(\DFF_923.Q ),
    .y(_02276_)
  );
  al_nand2ft _07396_ (
    .a(\DFF_923.Q ),
    .b(\DFF_827.Q ),
    .y(_02277_)
  );
  al_nand2ft _07397_ (
    .a(_02276_),
    .b(_02277_),
    .y(_02278_)
  );
  al_oa21ttf _07398_ (
    .a(_02274_),
    .b(_02275_),
    .c(_02278_),
    .y(_02279_)
  );
  al_nand3fft _07399_ (
    .a(_02274_),
    .b(_02275_),
    .c(_02278_),
    .y(_02280_)
  );
  al_and3fft _07400_ (
    .a(TM0),
    .b(_02279_),
    .c(_02280_),
    .y(_02281_)
  );
  al_nand2 _07401_ (
    .a(TM0),
    .b(\DFF_740.Q ),
    .y(_02282_)
  );
  al_or3fft _07402_ (
    .a(_01652_),
    .b(_02282_),
    .c(_02281_),
    .y(_02283_)
  );
  al_and2 _07403_ (
    .a(TM0),
    .b(\DFF_603.Q ),
    .y(_02284_)
  );
  al_and3fft _07404_ (
    .a(_02284_),
    .b(_01792_),
    .c(TM1),
    .y(_02285_)
  );
  al_nor3fft _07405_ (
    .a(RESET),
    .b(_02283_),
    .c(_02285_),
    .y(\DFF_635.D )
  );
  al_nor2 _07406_ (
    .a(\DFF_860.Q ),
    .b(\DFF_892.Q ),
    .y(_02286_)
  );
  al_and2 _07407_ (
    .a(\DFF_860.Q ),
    .b(\DFF_892.Q ),
    .y(_02287_)
  );
  al_and2ft _07408_ (
    .a(\DFF_828.Q ),
    .b(\DFF_924.Q ),
    .y(_02288_)
  );
  al_nand2ft _07409_ (
    .a(\DFF_924.Q ),
    .b(\DFF_828.Q ),
    .y(_02289_)
  );
  al_nand2ft _07410_ (
    .a(_02288_),
    .b(_02289_),
    .y(_02290_)
  );
  al_oa21ttf _07411_ (
    .a(_02286_),
    .b(_02287_),
    .c(_02290_),
    .y(_02291_)
  );
  al_nand3fft _07412_ (
    .a(_02286_),
    .b(_02287_),
    .c(_02290_),
    .y(_02292_)
  );
  al_and3fft _07413_ (
    .a(TM0),
    .b(_02291_),
    .c(_02292_),
    .y(_02293_)
  );
  al_nand2 _07414_ (
    .a(TM0),
    .b(\DFF_739.Q ),
    .y(_02294_)
  );
  al_or3fft _07415_ (
    .a(_01652_),
    .b(_02294_),
    .c(_02293_),
    .y(_02295_)
  );
  al_and2 _07416_ (
    .a(TM0),
    .b(\DFF_604.Q ),
    .y(_02296_)
  );
  al_and3fft _07417_ (
    .a(_02296_),
    .b(_01804_),
    .c(TM1),
    .y(_02297_)
  );
  al_nor3fft _07418_ (
    .a(RESET),
    .b(_02295_),
    .c(_02297_),
    .y(\DFF_636.D )
  );
  al_nor2 _07419_ (
    .a(\DFF_861.Q ),
    .b(\DFF_893.Q ),
    .y(_02298_)
  );
  al_and2 _07420_ (
    .a(\DFF_861.Q ),
    .b(\DFF_893.Q ),
    .y(_02299_)
  );
  al_and2ft _07421_ (
    .a(\DFF_829.Q ),
    .b(\DFF_925.Q ),
    .y(_02300_)
  );
  al_nand2ft _07422_ (
    .a(\DFF_925.Q ),
    .b(\DFF_829.Q ),
    .y(_02301_)
  );
  al_nand2ft _07423_ (
    .a(_02300_),
    .b(_02301_),
    .y(_02302_)
  );
  al_oa21ttf _07424_ (
    .a(_02298_),
    .b(_02299_),
    .c(_02302_),
    .y(_02303_)
  );
  al_nand3fft _07425_ (
    .a(_02298_),
    .b(_02299_),
    .c(_02302_),
    .y(_02304_)
  );
  al_and3fft _07426_ (
    .a(TM0),
    .b(_02303_),
    .c(_02304_),
    .y(_02305_)
  );
  al_nand2 _07427_ (
    .a(TM0),
    .b(\DFF_738.Q ),
    .y(_02306_)
  );
  al_or3fft _07428_ (
    .a(_01652_),
    .b(_02306_),
    .c(_02305_),
    .y(_02307_)
  );
  al_and2 _07429_ (
    .a(TM0),
    .b(\DFF_605.Q ),
    .y(_02308_)
  );
  al_and3fft _07430_ (
    .a(_02308_),
    .b(_01816_),
    .c(TM1),
    .y(_02309_)
  );
  al_nor3fft _07431_ (
    .a(RESET),
    .b(_02307_),
    .c(_02309_),
    .y(\DFF_637.D )
  );
  al_nor2 _07432_ (
    .a(\DFF_862.Q ),
    .b(\DFF_894.Q ),
    .y(_02310_)
  );
  al_and2 _07433_ (
    .a(\DFF_862.Q ),
    .b(\DFF_894.Q ),
    .y(_02311_)
  );
  al_and2ft _07434_ (
    .a(\DFF_830.Q ),
    .b(\DFF_926.Q ),
    .y(_02312_)
  );
  al_nand2ft _07435_ (
    .a(\DFF_926.Q ),
    .b(\DFF_830.Q ),
    .y(_02313_)
  );
  al_nand2ft _07436_ (
    .a(_02312_),
    .b(_02313_),
    .y(_02314_)
  );
  al_oa21ttf _07437_ (
    .a(_02310_),
    .b(_02311_),
    .c(_02314_),
    .y(_02315_)
  );
  al_nand3fft _07438_ (
    .a(_02310_),
    .b(_02311_),
    .c(_02314_),
    .y(_02316_)
  );
  al_and3fft _07439_ (
    .a(TM0),
    .b(_02315_),
    .c(_02316_),
    .y(_02317_)
  );
  al_nand2 _07440_ (
    .a(TM0),
    .b(\DFF_737.Q ),
    .y(_02318_)
  );
  al_or3fft _07441_ (
    .a(_01652_),
    .b(_02318_),
    .c(_02317_),
    .y(_02319_)
  );
  al_and2 _07442_ (
    .a(TM0),
    .b(\DFF_606.Q ),
    .y(_02320_)
  );
  al_and3fft _07443_ (
    .a(_02320_),
    .b(_01828_),
    .c(TM1),
    .y(_02321_)
  );
  al_nor3fft _07444_ (
    .a(RESET),
    .b(_02319_),
    .c(_02321_),
    .y(\DFF_638.D )
  );
  al_nor2 _07445_ (
    .a(\DFF_863.Q ),
    .b(\DFF_895.Q ),
    .y(_02322_)
  );
  al_and2 _07446_ (
    .a(\DFF_863.Q ),
    .b(\DFF_895.Q ),
    .y(_02323_)
  );
  al_and2ft _07447_ (
    .a(\DFF_831.Q ),
    .b(\DFF_927.Q ),
    .y(_02324_)
  );
  al_nand2ft _07448_ (
    .a(\DFF_927.Q ),
    .b(\DFF_831.Q ),
    .y(_02325_)
  );
  al_nand2ft _07449_ (
    .a(_02324_),
    .b(_02325_),
    .y(_02326_)
  );
  al_oa21ttf _07450_ (
    .a(_02322_),
    .b(_02323_),
    .c(_02326_),
    .y(_02327_)
  );
  al_nand3fft _07451_ (
    .a(_02322_),
    .b(_02323_),
    .c(_02326_),
    .y(_02328_)
  );
  al_and3fft _07452_ (
    .a(TM0),
    .b(_02327_),
    .c(_02328_),
    .y(_02329_)
  );
  al_nand2 _07453_ (
    .a(TM0),
    .b(\DFF_736.Q ),
    .y(_02330_)
  );
  al_or3fft _07454_ (
    .a(_01652_),
    .b(_02330_),
    .c(_02329_),
    .y(_02331_)
  );
  al_and2 _07455_ (
    .a(TM0),
    .b(\DFF_607.Q ),
    .y(_02332_)
  );
  al_and3fft _07456_ (
    .a(_02332_),
    .b(_01840_),
    .c(TM1),
    .y(_02333_)
  );
  al_nor3fft _07457_ (
    .a(RESET),
    .b(_02331_),
    .c(_02333_),
    .y(\DFF_639.D )
  );
  al_and2 _07458_ (
    .a(RESET),
    .b(\DFF_608.Q ),
    .y(\DFF_640.D )
  );
  al_and2 _07459_ (
    .a(RESET),
    .b(\DFF_609.Q ),
    .y(\DFF_641.D )
  );
  al_and2 _07460_ (
    .a(RESET),
    .b(\DFF_610.Q ),
    .y(\DFF_642.D )
  );
  al_and2 _07461_ (
    .a(RESET),
    .b(\DFF_611.Q ),
    .y(\DFF_643.D )
  );
  al_and2 _07462_ (
    .a(RESET),
    .b(\DFF_612.Q ),
    .y(\DFF_644.D )
  );
  al_and2 _07463_ (
    .a(RESET),
    .b(\DFF_613.Q ),
    .y(\DFF_645.D )
  );
  al_and2 _07464_ (
    .a(RESET),
    .b(\DFF_614.Q ),
    .y(\DFF_646.D )
  );
  al_and2 _07465_ (
    .a(RESET),
    .b(\DFF_615.Q ),
    .y(\DFF_647.D )
  );
  al_and2 _07466_ (
    .a(RESET),
    .b(\DFF_616.Q ),
    .y(\DFF_648.D )
  );
  al_and2 _07467_ (
    .a(RESET),
    .b(\DFF_617.Q ),
    .y(\DFF_649.D )
  );
  al_and2 _07468_ (
    .a(RESET),
    .b(\DFF_618.Q ),
    .y(\DFF_650.D )
  );
  al_and2 _07469_ (
    .a(RESET),
    .b(\DFF_619.Q ),
    .y(\DFF_651.D )
  );
  al_and2 _07470_ (
    .a(RESET),
    .b(\DFF_620.Q ),
    .y(\DFF_652.D )
  );
  al_and2 _07471_ (
    .a(RESET),
    .b(\DFF_621.Q ),
    .y(\DFF_653.D )
  );
  al_and2 _07472_ (
    .a(RESET),
    .b(\DFF_622.Q ),
    .y(\DFF_654.D )
  );
  al_and2 _07473_ (
    .a(RESET),
    .b(\DFF_623.Q ),
    .y(\DFF_655.D )
  );
  al_and2 _07474_ (
    .a(RESET),
    .b(\DFF_624.Q ),
    .y(\DFF_656.D )
  );
  al_and2 _07475_ (
    .a(RESET),
    .b(\DFF_625.Q ),
    .y(\DFF_657.D )
  );
  al_and2 _07476_ (
    .a(RESET),
    .b(\DFF_626.Q ),
    .y(\DFF_658.D )
  );
  al_and2 _07477_ (
    .a(RESET),
    .b(\DFF_627.Q ),
    .y(\DFF_659.D )
  );
  al_and2 _07478_ (
    .a(RESET),
    .b(\DFF_628.Q ),
    .y(\DFF_660.D )
  );
  al_and2 _07479_ (
    .a(RESET),
    .b(\DFF_629.Q ),
    .y(\DFF_661.D )
  );
  al_and2 _07480_ (
    .a(RESET),
    .b(\DFF_630.Q ),
    .y(\DFF_662.D )
  );
  al_and2 _07481_ (
    .a(RESET),
    .b(\DFF_631.Q ),
    .y(\DFF_663.D )
  );
  al_and2 _07482_ (
    .a(RESET),
    .b(\DFF_632.Q ),
    .y(\DFF_664.D )
  );
  al_and2 _07483_ (
    .a(RESET),
    .b(\DFF_633.Q ),
    .y(\DFF_665.D )
  );
  al_and2 _07484_ (
    .a(RESET),
    .b(\DFF_634.Q ),
    .y(\DFF_666.D )
  );
  al_and2 _07485_ (
    .a(RESET),
    .b(\DFF_635.Q ),
    .y(\DFF_667.D )
  );
  al_and2 _07486_ (
    .a(RESET),
    .b(\DFF_636.Q ),
    .y(\DFF_668.D )
  );
  al_and2 _07487_ (
    .a(RESET),
    .b(\DFF_637.Q ),
    .y(\DFF_669.D )
  );
  al_and2 _07488_ (
    .a(RESET),
    .b(\DFF_638.Q ),
    .y(\DFF_670.D )
  );
  al_and2 _07489_ (
    .a(RESET),
    .b(\DFF_639.Q ),
    .y(\DFF_671.D )
  );
  al_and2 _07490_ (
    .a(RESET),
    .b(\DFF_640.Q ),
    .y(\DFF_672.D )
  );
  al_and2 _07491_ (
    .a(RESET),
    .b(\DFF_641.Q ),
    .y(\DFF_673.D )
  );
  al_and2 _07492_ (
    .a(RESET),
    .b(\DFF_642.Q ),
    .y(\DFF_674.D )
  );
  al_and2 _07493_ (
    .a(RESET),
    .b(\DFF_643.Q ),
    .y(\DFF_675.D )
  );
  al_and2 _07494_ (
    .a(RESET),
    .b(\DFF_644.Q ),
    .y(\DFF_676.D )
  );
  al_and2 _07495_ (
    .a(RESET),
    .b(\DFF_645.Q ),
    .y(\DFF_677.D )
  );
  al_and2 _07496_ (
    .a(RESET),
    .b(\DFF_646.Q ),
    .y(\DFF_678.D )
  );
  al_and2 _07497_ (
    .a(RESET),
    .b(\DFF_647.Q ),
    .y(\DFF_679.D )
  );
  al_and2 _07498_ (
    .a(RESET),
    .b(\DFF_648.Q ),
    .y(\DFF_680.D )
  );
  al_and2 _07499_ (
    .a(RESET),
    .b(\DFF_649.Q ),
    .y(\DFF_681.D )
  );
  al_and2 _07500_ (
    .a(RESET),
    .b(\DFF_650.Q ),
    .y(\DFF_682.D )
  );
  al_and2 _07501_ (
    .a(RESET),
    .b(\DFF_651.Q ),
    .y(\DFF_683.D )
  );
  al_and2 _07502_ (
    .a(RESET),
    .b(\DFF_652.Q ),
    .y(\DFF_684.D )
  );
  al_and2 _07503_ (
    .a(RESET),
    .b(\DFF_653.Q ),
    .y(\DFF_685.D )
  );
  al_and2 _07504_ (
    .a(RESET),
    .b(\DFF_654.Q ),
    .y(\DFF_686.D )
  );
  al_and2 _07505_ (
    .a(RESET),
    .b(\DFF_655.Q ),
    .y(\DFF_687.D )
  );
  al_and2 _07506_ (
    .a(RESET),
    .b(\DFF_656.Q ),
    .y(\DFF_688.D )
  );
  al_and2 _07507_ (
    .a(RESET),
    .b(\DFF_657.Q ),
    .y(\DFF_689.D )
  );
  al_and2 _07508_ (
    .a(RESET),
    .b(\DFF_658.Q ),
    .y(\DFF_690.D )
  );
  al_and2 _07509_ (
    .a(RESET),
    .b(\DFF_659.Q ),
    .y(\DFF_691.D )
  );
  al_and2 _07510_ (
    .a(RESET),
    .b(\DFF_660.Q ),
    .y(\DFF_692.D )
  );
  al_and2 _07511_ (
    .a(RESET),
    .b(\DFF_661.Q ),
    .y(\DFF_693.D )
  );
  al_and2 _07512_ (
    .a(RESET),
    .b(\DFF_662.Q ),
    .y(\DFF_694.D )
  );
  al_and2 _07513_ (
    .a(RESET),
    .b(\DFF_663.Q ),
    .y(\DFF_695.D )
  );
  al_and2 _07514_ (
    .a(RESET),
    .b(\DFF_664.Q ),
    .y(\DFF_696.D )
  );
  al_and2 _07515_ (
    .a(RESET),
    .b(\DFF_665.Q ),
    .y(\DFF_697.D )
  );
  al_and2 _07516_ (
    .a(RESET),
    .b(\DFF_666.Q ),
    .y(\DFF_698.D )
  );
  al_and2 _07517_ (
    .a(RESET),
    .b(\DFF_667.Q ),
    .y(\DFF_699.D )
  );
  al_and2 _07518_ (
    .a(RESET),
    .b(\DFF_668.Q ),
    .y(\DFF_700.D )
  );
  al_and2 _07519_ (
    .a(RESET),
    .b(\DFF_669.Q ),
    .y(\DFF_701.D )
  );
  al_and2 _07520_ (
    .a(RESET),
    .b(\DFF_670.Q ),
    .y(\DFF_702.D )
  );
  al_and2 _07521_ (
    .a(RESET),
    .b(\DFF_671.Q ),
    .y(\DFF_703.D )
  );
  al_and2 _07522_ (
    .a(RESET),
    .b(\DFF_672.Q ),
    .y(\DFF_704.D )
  );
  al_and2 _07523_ (
    .a(RESET),
    .b(\DFF_673.Q ),
    .y(\DFF_705.D )
  );
  al_and2 _07524_ (
    .a(RESET),
    .b(\DFF_674.Q ),
    .y(\DFF_706.D )
  );
  al_and2 _07525_ (
    .a(RESET),
    .b(\DFF_675.Q ),
    .y(\DFF_707.D )
  );
  al_and2 _07526_ (
    .a(RESET),
    .b(\DFF_676.Q ),
    .y(\DFF_708.D )
  );
  al_and2 _07527_ (
    .a(RESET),
    .b(\DFF_677.Q ),
    .y(\DFF_709.D )
  );
  al_and2 _07528_ (
    .a(RESET),
    .b(\DFF_678.Q ),
    .y(\DFF_710.D )
  );
  al_and2 _07529_ (
    .a(RESET),
    .b(\DFF_679.Q ),
    .y(\DFF_711.D )
  );
  al_and2 _07530_ (
    .a(RESET),
    .b(\DFF_680.Q ),
    .y(\DFF_712.D )
  );
  al_and2 _07531_ (
    .a(RESET),
    .b(\DFF_681.Q ),
    .y(\DFF_713.D )
  );
  al_and2 _07532_ (
    .a(RESET),
    .b(\DFF_682.Q ),
    .y(\DFF_714.D )
  );
  al_and2 _07533_ (
    .a(RESET),
    .b(\DFF_683.Q ),
    .y(\DFF_715.D )
  );
  al_and2 _07534_ (
    .a(RESET),
    .b(\DFF_684.Q ),
    .y(\DFF_716.D )
  );
  al_and2 _07535_ (
    .a(RESET),
    .b(\DFF_685.Q ),
    .y(\DFF_717.D )
  );
  al_and2 _07536_ (
    .a(RESET),
    .b(\DFF_686.Q ),
    .y(\DFF_718.D )
  );
  al_and2 _07537_ (
    .a(RESET),
    .b(\DFF_687.Q ),
    .y(\DFF_719.D )
  );
  al_and2 _07538_ (
    .a(RESET),
    .b(\DFF_688.Q ),
    .y(\DFF_720.D )
  );
  al_and2 _07539_ (
    .a(RESET),
    .b(\DFF_689.Q ),
    .y(\DFF_721.D )
  );
  al_and2 _07540_ (
    .a(RESET),
    .b(\DFF_690.Q ),
    .y(\DFF_722.D )
  );
  al_and2 _07541_ (
    .a(RESET),
    .b(\DFF_691.Q ),
    .y(\DFF_723.D )
  );
  al_and2 _07542_ (
    .a(RESET),
    .b(\DFF_692.Q ),
    .y(\DFF_724.D )
  );
  al_and2 _07543_ (
    .a(RESET),
    .b(\DFF_693.Q ),
    .y(\DFF_725.D )
  );
  al_and2 _07544_ (
    .a(RESET),
    .b(\DFF_694.Q ),
    .y(\DFF_726.D )
  );
  al_and2 _07545_ (
    .a(RESET),
    .b(\DFF_695.Q ),
    .y(\DFF_727.D )
  );
  al_and2 _07546_ (
    .a(RESET),
    .b(\DFF_696.Q ),
    .y(\DFF_728.D )
  );
  al_and2 _07547_ (
    .a(RESET),
    .b(\DFF_697.Q ),
    .y(\DFF_729.D )
  );
  al_and2 _07548_ (
    .a(RESET),
    .b(\DFF_698.Q ),
    .y(\DFF_730.D )
  );
  al_and2 _07549_ (
    .a(RESET),
    .b(\DFF_699.Q ),
    .y(\DFF_731.D )
  );
  al_and2 _07550_ (
    .a(RESET),
    .b(\DFF_700.Q ),
    .y(\DFF_732.D )
  );
  al_and2 _07551_ (
    .a(RESET),
    .b(\DFF_701.Q ),
    .y(\DFF_733.D )
  );
  al_and2 _07552_ (
    .a(RESET),
    .b(\DFF_702.Q ),
    .y(\DFF_734.D )
  );
  al_and2 _07553_ (
    .a(RESET),
    .b(\DFF_703.Q ),
    .y(\DFF_735.D )
  );
  al_oa21ftt _07554_ (
    .a(\DFF_735.Q ),
    .b(\DFF_767.Q ),
    .c(RESET),
    .y(_02334_)
  );
  al_aoi21ftf _07555_ (
    .a(\DFF_735.Q ),
    .b(\DFF_767.Q ),
    .c(_02334_),
    .y(\DFF_736.D )
  );
  al_oa21ftt _07556_ (
    .a(\DFF_734.Q ),
    .b(\DFF_736.Q ),
    .c(RESET),
    .y(_02335_)
  );
  al_aoi21ftf _07557_ (
    .a(\DFF_734.Q ),
    .b(\DFF_736.Q ),
    .c(_02335_),
    .y(\DFF_737.D )
  );
  al_oa21ftt _07558_ (
    .a(\DFF_733.Q ),
    .b(\DFF_737.Q ),
    .c(RESET),
    .y(_02336_)
  );
  al_aoi21ftf _07559_ (
    .a(\DFF_733.Q ),
    .b(\DFF_737.Q ),
    .c(_02336_),
    .y(\DFF_738.D )
  );
  al_oa21ftt _07560_ (
    .a(\DFF_732.Q ),
    .b(\DFF_738.Q ),
    .c(RESET),
    .y(_02337_)
  );
  al_aoi21ftf _07561_ (
    .a(\DFF_732.Q ),
    .b(\DFF_738.Q ),
    .c(_02337_),
    .y(\DFF_739.D )
  );
  al_nand2ft _07562_ (
    .a(\DFF_731.Q ),
    .b(\DFF_739.Q ),
    .y(_02338_)
  );
  al_nand2ft _07563_ (
    .a(\DFF_739.Q ),
    .b(\DFF_731.Q ),
    .y(_02339_)
  );
  al_ao21ttf _07564_ (
    .a(_02338_),
    .b(_02339_),
    .c(\DFF_767.Q ),
    .y(_02340_)
  );
  al_nand3ftt _07565_ (
    .a(\DFF_767.Q ),
    .b(_02338_),
    .c(_02339_),
    .y(_02341_)
  );
  al_aoi21 _07566_ (
    .a(_02341_),
    .b(_02340_),
    .c(_00451_),
    .y(\DFF_740.D )
  );
  al_oa21ftt _07567_ (
    .a(\DFF_730.Q ),
    .b(\DFF_740.Q ),
    .c(RESET),
    .y(_02342_)
  );
  al_aoi21ftf _07568_ (
    .a(\DFF_730.Q ),
    .b(\DFF_740.Q ),
    .c(_02342_),
    .y(\DFF_741.D )
  );
  al_oa21ftt _07569_ (
    .a(\DFF_729.Q ),
    .b(\DFF_741.Q ),
    .c(RESET),
    .y(_02343_)
  );
  al_aoi21ftf _07570_ (
    .a(\DFF_729.Q ),
    .b(\DFF_741.Q ),
    .c(_02343_),
    .y(\DFF_742.D )
  );
  al_oa21ftt _07571_ (
    .a(\DFF_728.Q ),
    .b(\DFF_742.Q ),
    .c(RESET),
    .y(_02344_)
  );
  al_aoi21ftf _07572_ (
    .a(\DFF_728.Q ),
    .b(\DFF_742.Q ),
    .c(_02344_),
    .y(\DFF_743.D )
  );
  al_oa21ftt _07573_ (
    .a(\DFF_727.Q ),
    .b(\DFF_743.Q ),
    .c(RESET),
    .y(_02345_)
  );
  al_aoi21ftf _07574_ (
    .a(\DFF_727.Q ),
    .b(\DFF_743.Q ),
    .c(_02345_),
    .y(\DFF_744.D )
  );
  al_oa21ftt _07575_ (
    .a(\DFF_726.Q ),
    .b(\DFF_744.Q ),
    .c(RESET),
    .y(_02346_)
  );
  al_aoi21ftf _07576_ (
    .a(\DFF_726.Q ),
    .b(\DFF_744.Q ),
    .c(_02346_),
    .y(\DFF_745.D )
  );
  al_oa21ftt _07577_ (
    .a(\DFF_725.Q ),
    .b(\DFF_745.Q ),
    .c(RESET),
    .y(_02347_)
  );
  al_aoi21ftf _07578_ (
    .a(\DFF_725.Q ),
    .b(\DFF_745.Q ),
    .c(_02347_),
    .y(\DFF_746.D )
  );
  al_nand2ft _07579_ (
    .a(\DFF_724.Q ),
    .b(\DFF_746.Q ),
    .y(_02348_)
  );
  al_nand2ft _07580_ (
    .a(\DFF_746.Q ),
    .b(\DFF_724.Q ),
    .y(_02349_)
  );
  al_ao21ttf _07581_ (
    .a(_02348_),
    .b(_02349_),
    .c(\DFF_767.Q ),
    .y(_02350_)
  );
  al_nand3ftt _07582_ (
    .a(\DFF_767.Q ),
    .b(_02348_),
    .c(_02349_),
    .y(_02351_)
  );
  al_aoi21 _07583_ (
    .a(_02351_),
    .b(_02350_),
    .c(_00451_),
    .y(\DFF_747.D )
  );
  al_oa21ftt _07584_ (
    .a(\DFF_723.Q ),
    .b(\DFF_747.Q ),
    .c(RESET),
    .y(_02352_)
  );
  al_aoi21ftf _07585_ (
    .a(\DFF_723.Q ),
    .b(\DFF_747.Q ),
    .c(_02352_),
    .y(\DFF_748.D )
  );
  al_oa21ftt _07586_ (
    .a(\DFF_722.Q ),
    .b(\DFF_748.Q ),
    .c(RESET),
    .y(_02353_)
  );
  al_aoi21ftf _07587_ (
    .a(\DFF_722.Q ),
    .b(\DFF_748.Q ),
    .c(_02353_),
    .y(\DFF_749.D )
  );
  al_oa21ftt _07588_ (
    .a(\DFF_721.Q ),
    .b(\DFF_749.Q ),
    .c(RESET),
    .y(_02354_)
  );
  al_aoi21ftf _07589_ (
    .a(\DFF_721.Q ),
    .b(\DFF_749.Q ),
    .c(_02354_),
    .y(\DFF_750.D )
  );
  al_oa21ftt _07590_ (
    .a(\DFF_720.Q ),
    .b(\DFF_750.Q ),
    .c(RESET),
    .y(_02355_)
  );
  al_aoi21ftf _07591_ (
    .a(\DFF_720.Q ),
    .b(\DFF_750.Q ),
    .c(_02355_),
    .y(\DFF_751.D )
  );
  al_nand2ft _07592_ (
    .a(\DFF_719.Q ),
    .b(\DFF_751.Q ),
    .y(_02356_)
  );
  al_nand2ft _07593_ (
    .a(\DFF_751.Q ),
    .b(\DFF_719.Q ),
    .y(_02357_)
  );
  al_ao21ttf _07594_ (
    .a(_02356_),
    .b(_02357_),
    .c(\DFF_767.Q ),
    .y(_02358_)
  );
  al_nand3ftt _07595_ (
    .a(\DFF_767.Q ),
    .b(_02356_),
    .c(_02357_),
    .y(_02359_)
  );
  al_aoi21 _07596_ (
    .a(_02359_),
    .b(_02358_),
    .c(_00451_),
    .y(\DFF_752.D )
  );
  al_oa21ftt _07597_ (
    .a(\DFF_718.Q ),
    .b(\DFF_752.Q ),
    .c(RESET),
    .y(_02360_)
  );
  al_aoi21ftf _07598_ (
    .a(\DFF_718.Q ),
    .b(\DFF_752.Q ),
    .c(_02360_),
    .y(\DFF_753.D )
  );
  al_oa21ftt _07599_ (
    .a(\DFF_717.Q ),
    .b(\DFF_753.Q ),
    .c(RESET),
    .y(_02361_)
  );
  al_aoi21ftf _07600_ (
    .a(\DFF_717.Q ),
    .b(\DFF_753.Q ),
    .c(_02361_),
    .y(\DFF_754.D )
  );
  al_oa21ftt _07601_ (
    .a(\DFF_716.Q ),
    .b(\DFF_754.Q ),
    .c(RESET),
    .y(_02362_)
  );
  al_aoi21ftf _07602_ (
    .a(\DFF_716.Q ),
    .b(\DFF_754.Q ),
    .c(_02362_),
    .y(\DFF_755.D )
  );
  al_oa21ftt _07603_ (
    .a(\DFF_715.Q ),
    .b(\DFF_755.Q ),
    .c(RESET),
    .y(_02363_)
  );
  al_aoi21ftf _07604_ (
    .a(\DFF_715.Q ),
    .b(\DFF_755.Q ),
    .c(_02363_),
    .y(\DFF_756.D )
  );
  al_oa21ftt _07605_ (
    .a(\DFF_714.Q ),
    .b(\DFF_756.Q ),
    .c(RESET),
    .y(_02364_)
  );
  al_aoi21ftf _07606_ (
    .a(\DFF_714.Q ),
    .b(\DFF_756.Q ),
    .c(_02364_),
    .y(\DFF_757.D )
  );
  al_oa21ftt _07607_ (
    .a(\DFF_713.Q ),
    .b(\DFF_757.Q ),
    .c(RESET),
    .y(_02365_)
  );
  al_aoi21ftf _07608_ (
    .a(\DFF_713.Q ),
    .b(\DFF_757.Q ),
    .c(_02365_),
    .y(\DFF_758.D )
  );
  al_oa21ftt _07609_ (
    .a(\DFF_712.Q ),
    .b(\DFF_758.Q ),
    .c(RESET),
    .y(_02366_)
  );
  al_aoi21ftf _07610_ (
    .a(\DFF_712.Q ),
    .b(\DFF_758.Q ),
    .c(_02366_),
    .y(\DFF_759.D )
  );
  al_oa21ftt _07611_ (
    .a(\DFF_711.Q ),
    .b(\DFF_759.Q ),
    .c(RESET),
    .y(_02367_)
  );
  al_aoi21ftf _07612_ (
    .a(\DFF_711.Q ),
    .b(\DFF_759.Q ),
    .c(_02367_),
    .y(\DFF_760.D )
  );
  al_oa21ftt _07613_ (
    .a(\DFF_710.Q ),
    .b(\DFF_760.Q ),
    .c(RESET),
    .y(_02368_)
  );
  al_aoi21ftf _07614_ (
    .a(\DFF_710.Q ),
    .b(\DFF_760.Q ),
    .c(_02368_),
    .y(\DFF_761.D )
  );
  al_oa21ftt _07615_ (
    .a(\DFF_709.Q ),
    .b(\DFF_761.Q ),
    .c(RESET),
    .y(_02369_)
  );
  al_aoi21ftf _07616_ (
    .a(\DFF_709.Q ),
    .b(\DFF_761.Q ),
    .c(_02369_),
    .y(\DFF_762.D )
  );
  al_oa21ftt _07617_ (
    .a(\DFF_708.Q ),
    .b(\DFF_762.Q ),
    .c(RESET),
    .y(_02370_)
  );
  al_aoi21ftf _07618_ (
    .a(\DFF_708.Q ),
    .b(\DFF_762.Q ),
    .c(_02370_),
    .y(\DFF_763.D )
  );
  al_oa21ftt _07619_ (
    .a(\DFF_707.Q ),
    .b(\DFF_763.Q ),
    .c(RESET),
    .y(_02371_)
  );
  al_aoi21ftf _07620_ (
    .a(\DFF_707.Q ),
    .b(\DFF_763.Q ),
    .c(_02371_),
    .y(\DFF_764.D )
  );
  al_oa21ftt _07621_ (
    .a(\DFF_706.Q ),
    .b(\DFF_764.Q ),
    .c(RESET),
    .y(_02372_)
  );
  al_aoi21ftf _07622_ (
    .a(\DFF_706.Q ),
    .b(\DFF_764.Q ),
    .c(_02372_),
    .y(\DFF_765.D )
  );
  al_oa21ftt _07623_ (
    .a(\DFF_705.Q ),
    .b(\DFF_765.Q ),
    .c(RESET),
    .y(_02373_)
  );
  al_aoi21ftf _07624_ (
    .a(\DFF_705.Q ),
    .b(\DFF_765.Q ),
    .c(_02373_),
    .y(\DFF_766.D )
  );
  al_oa21ftt _07625_ (
    .a(\DFF_704.Q ),
    .b(\DFF_766.Q ),
    .c(RESET),
    .y(_02374_)
  );
  al_aoi21ftf _07626_ (
    .a(\DFF_704.Q ),
    .b(\DFF_766.Q ),
    .c(_02374_),
    .y(\DFF_767.D )
  );
  al_and2 _07627_ (
    .a(RESET),
    .b(\DFF_769.Q ),
    .y(\DFF_768.D )
  );
  al_and2 _07628_ (
    .a(RESET),
    .b(\DFF_770.Q ),
    .y(\DFF_769.D )
  );
  al_and2 _07629_ (
    .a(RESET),
    .b(\DFF_771.Q ),
    .y(\DFF_770.D )
  );
  al_and2 _07630_ (
    .a(RESET),
    .b(\DFF_772.Q ),
    .y(\DFF_771.D )
  );
  al_and2 _07631_ (
    .a(RESET),
    .b(\DFF_773.Q ),
    .y(\DFF_772.D )
  );
  al_and2 _07632_ (
    .a(RESET),
    .b(\DFF_774.Q ),
    .y(\DFF_773.D )
  );
  al_and2 _07633_ (
    .a(RESET),
    .b(\DFF_775.Q ),
    .y(\DFF_774.D )
  );
  al_and2 _07634_ (
    .a(RESET),
    .b(\DFF_776.Q ),
    .y(\DFF_775.D )
  );
  al_and2 _07635_ (
    .a(RESET),
    .b(\DFF_777.Q ),
    .y(\DFF_776.D )
  );
  al_and2 _07636_ (
    .a(RESET),
    .b(\DFF_778.Q ),
    .y(\DFF_777.D )
  );
  al_and2 _07637_ (
    .a(RESET),
    .b(\DFF_779.Q ),
    .y(\DFF_778.D )
  );
  al_and2 _07638_ (
    .a(RESET),
    .b(\DFF_780.Q ),
    .y(\DFF_779.D )
  );
  al_and2 _07639_ (
    .a(RESET),
    .b(\DFF_781.Q ),
    .y(\DFF_780.D )
  );
  al_and2 _07640_ (
    .a(RESET),
    .b(\DFF_782.Q ),
    .y(\DFF_781.D )
  );
  al_and2 _07641_ (
    .a(RESET),
    .b(\DFF_783.Q ),
    .y(\DFF_782.D )
  );
  al_and2 _07642_ (
    .a(RESET),
    .b(\DFF_784.Q ),
    .y(\DFF_783.D )
  );
  al_and2 _07643_ (
    .a(RESET),
    .b(\DFF_785.Q ),
    .y(\DFF_784.D )
  );
  al_and2 _07644_ (
    .a(RESET),
    .b(\DFF_786.Q ),
    .y(\DFF_785.D )
  );
  al_and2 _07645_ (
    .a(RESET),
    .b(\DFF_787.Q ),
    .y(\DFF_786.D )
  );
  al_and2 _07646_ (
    .a(RESET),
    .b(\DFF_788.Q ),
    .y(\DFF_787.D )
  );
  al_and2 _07647_ (
    .a(RESET),
    .b(\DFF_789.Q ),
    .y(\DFF_788.D )
  );
  al_and2 _07648_ (
    .a(RESET),
    .b(\DFF_790.Q ),
    .y(\DFF_789.D )
  );
  al_and2 _07649_ (
    .a(RESET),
    .b(\DFF_791.Q ),
    .y(\DFF_790.D )
  );
  al_and2 _07650_ (
    .a(RESET),
    .b(\DFF_792.Q ),
    .y(\DFF_791.D )
  );
  al_and2 _07651_ (
    .a(RESET),
    .b(\DFF_793.Q ),
    .y(\DFF_792.D )
  );
  al_and2 _07652_ (
    .a(RESET),
    .b(\DFF_794.Q ),
    .y(\DFF_793.D )
  );
  al_and2 _07653_ (
    .a(RESET),
    .b(\DFF_795.Q ),
    .y(\DFF_794.D )
  );
  al_and2 _07654_ (
    .a(RESET),
    .b(\DFF_796.Q ),
    .y(\DFF_795.D )
  );
  al_and2 _07655_ (
    .a(RESET),
    .b(\DFF_797.Q ),
    .y(\DFF_796.D )
  );
  al_and2 _07656_ (
    .a(RESET),
    .b(\DFF_798.Q ),
    .y(\DFF_797.D )
  );
  al_and2 _07657_ (
    .a(RESET),
    .b(\DFF_799.Q ),
    .y(\DFF_798.D )
  );
  al_and2ft _07658_ (
    .a(\DFF_768.Q ),
    .b(RESET),
    .y(\DFF_799.D )
  );
  al_or2 _07659_ (
    .a(TM1),
    .b(\DFF_1056.Q ),
    .y(_02375_)
  );
  al_nand2 _07660_ (
    .a(TM1),
    .b(\DFF_1056.Q ),
    .y(_02376_)
  );
  al_nand3 _07661_ (
    .a(\DFF_1088.Q ),
    .b(_02375_),
    .c(_02376_),
    .y(_02377_)
  );
  al_nand2ft _07662_ (
    .a(TM1),
    .b(\DFF_1056.Q ),
    .y(_02378_)
  );
  al_and2ft _07663_ (
    .a(\DFF_1056.Q ),
    .b(TM1),
    .y(_02379_)
  );
  al_and3fft _07664_ (
    .a(\DFF_1088.Q ),
    .b(_02379_),
    .c(_02378_),
    .y(_02380_)
  );
  al_and2ft _07665_ (
    .a(\DFF_1024.Q ),
    .b(\DFF_992.Q ),
    .y(_02381_)
  );
  al_nand2ft _07666_ (
    .a(\DFF_992.Q ),
    .b(\DFF_1024.Q ),
    .y(_02382_)
  );
  al_nand2ft _07667_ (
    .a(_02381_),
    .b(_02382_),
    .y(_02383_)
  );
  al_oai21ftf _07668_ (
    .a(_02377_),
    .b(_02380_),
    .c(_02383_),
    .y(_02384_)
  );
  al_nand3ftt _07669_ (
    .a(_02380_),
    .b(_02377_),
    .c(_02383_),
    .y(_02385_)
  );
  al_nand3 _07670_ (
    .a(_00448_),
    .b(_02384_),
    .c(_02385_),
    .y(_02386_)
  );
  al_aoi21 _07671_ (
    .a(TM0),
    .b(\DFF_959.Q ),
    .c(TM1),
    .y(_02387_)
  );
  al_nand2 _07672_ (
    .a(_02387_),
    .b(_02386_),
    .y(_02388_)
  );
  al_aoi21ttf _07673_ (
    .a(\DFF_768.Q ),
    .b(TM0),
    .c(TM1),
    .y(_02389_)
  );
  al_and2 _07674_ (
    .a(_02389_),
    .b(_01897_),
    .y(_02390_)
  );
  al_nor3fft _07675_ (
    .a(RESET),
    .b(_02388_),
    .c(_02390_),
    .y(\DFF_800.D )
  );
  al_or2 _07676_ (
    .a(TM1),
    .b(\DFF_1057.Q ),
    .y(_02391_)
  );
  al_nand2 _07677_ (
    .a(TM1),
    .b(\DFF_1057.Q ),
    .y(_02392_)
  );
  al_nand3 _07678_ (
    .a(\DFF_1089.Q ),
    .b(_02391_),
    .c(_02392_),
    .y(_02393_)
  );
  al_nand2ft _07679_ (
    .a(TM1),
    .b(\DFF_1057.Q ),
    .y(_02394_)
  );
  al_and2ft _07680_ (
    .a(\DFF_1057.Q ),
    .b(TM1),
    .y(_02395_)
  );
  al_and3fft _07681_ (
    .a(\DFF_1089.Q ),
    .b(_02395_),
    .c(_02394_),
    .y(_02396_)
  );
  al_and2ft _07682_ (
    .a(\DFF_1025.Q ),
    .b(\DFF_993.Q ),
    .y(_02397_)
  );
  al_nand2ft _07683_ (
    .a(\DFF_993.Q ),
    .b(\DFF_1025.Q ),
    .y(_02398_)
  );
  al_nand2ft _07684_ (
    .a(_02397_),
    .b(_02398_),
    .y(_02399_)
  );
  al_oai21ftf _07685_ (
    .a(_02393_),
    .b(_02396_),
    .c(_02399_),
    .y(_02400_)
  );
  al_nand3ftt _07686_ (
    .a(_02396_),
    .b(_02393_),
    .c(_02399_),
    .y(_02401_)
  );
  al_nand3 _07687_ (
    .a(_00448_),
    .b(_02400_),
    .c(_02401_),
    .y(_02402_)
  );
  al_aoi21 _07688_ (
    .a(TM0),
    .b(\DFF_958.Q ),
    .c(TM1),
    .y(_02403_)
  );
  al_nand2 _07689_ (
    .a(_02403_),
    .b(_02402_),
    .y(_02404_)
  );
  al_aoi21ttf _07690_ (
    .a(TM0),
    .b(\DFF_769.Q ),
    .c(TM1),
    .y(_02405_)
  );
  al_and2 _07691_ (
    .a(_02405_),
    .b(_01913_),
    .y(_02406_)
  );
  al_nor3fft _07692_ (
    .a(RESET),
    .b(_02404_),
    .c(_02406_),
    .y(\DFF_801.D )
  );
  al_or2 _07693_ (
    .a(TM1),
    .b(\DFF_1058.Q ),
    .y(_02407_)
  );
  al_nand2 _07694_ (
    .a(TM1),
    .b(\DFF_1058.Q ),
    .y(_02408_)
  );
  al_nand3 _07695_ (
    .a(\DFF_1090.Q ),
    .b(_02407_),
    .c(_02408_),
    .y(_02409_)
  );
  al_nand2ft _07696_ (
    .a(TM1),
    .b(\DFF_1058.Q ),
    .y(_02410_)
  );
  al_and2ft _07697_ (
    .a(\DFF_1058.Q ),
    .b(TM1),
    .y(_02411_)
  );
  al_and3fft _07698_ (
    .a(\DFF_1090.Q ),
    .b(_02411_),
    .c(_02410_),
    .y(_02412_)
  );
  al_and2ft _07699_ (
    .a(\DFF_1026.Q ),
    .b(\DFF_994.Q ),
    .y(_02413_)
  );
  al_nand2ft _07700_ (
    .a(\DFF_994.Q ),
    .b(\DFF_1026.Q ),
    .y(_02414_)
  );
  al_nand2ft _07701_ (
    .a(_02413_),
    .b(_02414_),
    .y(_02415_)
  );
  al_oai21ftf _07702_ (
    .a(_02409_),
    .b(_02412_),
    .c(_02415_),
    .y(_02416_)
  );
  al_nand3ftt _07703_ (
    .a(_02412_),
    .b(_02409_),
    .c(_02415_),
    .y(_02417_)
  );
  al_nand3 _07704_ (
    .a(_00448_),
    .b(_02416_),
    .c(_02417_),
    .y(_02418_)
  );
  al_aoi21 _07705_ (
    .a(TM0),
    .b(\DFF_957.Q ),
    .c(TM1),
    .y(_02419_)
  );
  al_nand2 _07706_ (
    .a(_02419_),
    .b(_02418_),
    .y(_02420_)
  );
  al_aoi21ttf _07707_ (
    .a(TM0),
    .b(\DFF_770.Q ),
    .c(TM1),
    .y(_02421_)
  );
  al_and2 _07708_ (
    .a(_02421_),
    .b(_01929_),
    .y(_02422_)
  );
  al_nor3fft _07709_ (
    .a(RESET),
    .b(_02420_),
    .c(_02422_),
    .y(\DFF_802.D )
  );
  al_or2 _07710_ (
    .a(TM1),
    .b(\DFF_1059.Q ),
    .y(_02423_)
  );
  al_nand2 _07711_ (
    .a(TM1),
    .b(\DFF_1059.Q ),
    .y(_02424_)
  );
  al_nand3 _07712_ (
    .a(\DFF_1091.Q ),
    .b(_02423_),
    .c(_02424_),
    .y(_02425_)
  );
  al_nand2ft _07713_ (
    .a(TM1),
    .b(\DFF_1059.Q ),
    .y(_02426_)
  );
  al_and2ft _07714_ (
    .a(\DFF_1059.Q ),
    .b(TM1),
    .y(_02427_)
  );
  al_and3fft _07715_ (
    .a(\DFF_1091.Q ),
    .b(_02427_),
    .c(_02426_),
    .y(_02428_)
  );
  al_and2ft _07716_ (
    .a(\DFF_1027.Q ),
    .b(\DFF_995.Q ),
    .y(_02429_)
  );
  al_nand2ft _07717_ (
    .a(\DFF_995.Q ),
    .b(\DFF_1027.Q ),
    .y(_02430_)
  );
  al_nand2ft _07718_ (
    .a(_02429_),
    .b(_02430_),
    .y(_02431_)
  );
  al_oai21ftf _07719_ (
    .a(_02425_),
    .b(_02428_),
    .c(_02431_),
    .y(_02432_)
  );
  al_nand3ftt _07720_ (
    .a(_02428_),
    .b(_02425_),
    .c(_02431_),
    .y(_02433_)
  );
  al_nand3 _07721_ (
    .a(_00448_),
    .b(_02432_),
    .c(_02433_),
    .y(_02434_)
  );
  al_aoi21 _07722_ (
    .a(TM0),
    .b(\DFF_956.Q ),
    .c(TM1),
    .y(_02435_)
  );
  al_nand2 _07723_ (
    .a(_02435_),
    .b(_02434_),
    .y(_02436_)
  );
  al_aoi21ttf _07724_ (
    .a(TM0),
    .b(\DFF_771.Q ),
    .c(TM1),
    .y(_02437_)
  );
  al_and2 _07725_ (
    .a(_02437_),
    .b(_01945_),
    .y(_02438_)
  );
  al_nor3fft _07726_ (
    .a(RESET),
    .b(_02436_),
    .c(_02438_),
    .y(\DFF_803.D )
  );
  al_or2 _07727_ (
    .a(TM1),
    .b(\DFF_1060.Q ),
    .y(_02439_)
  );
  al_nand2 _07728_ (
    .a(TM1),
    .b(\DFF_1060.Q ),
    .y(_02440_)
  );
  al_nand3 _07729_ (
    .a(\DFF_1092.Q ),
    .b(_02439_),
    .c(_02440_),
    .y(_02441_)
  );
  al_nand2ft _07730_ (
    .a(TM1),
    .b(\DFF_1060.Q ),
    .y(_02442_)
  );
  al_and2ft _07731_ (
    .a(\DFF_1060.Q ),
    .b(TM1),
    .y(_02443_)
  );
  al_and3fft _07732_ (
    .a(\DFF_1092.Q ),
    .b(_02443_),
    .c(_02442_),
    .y(_02444_)
  );
  al_and2ft _07733_ (
    .a(\DFF_1028.Q ),
    .b(\DFF_996.Q ),
    .y(_02445_)
  );
  al_nand2ft _07734_ (
    .a(\DFF_996.Q ),
    .b(\DFF_1028.Q ),
    .y(_02446_)
  );
  al_nand2ft _07735_ (
    .a(_02445_),
    .b(_02446_),
    .y(_02447_)
  );
  al_oai21ftf _07736_ (
    .a(_02441_),
    .b(_02444_),
    .c(_02447_),
    .y(_02448_)
  );
  al_nand3ftt _07737_ (
    .a(_02444_),
    .b(_02441_),
    .c(_02447_),
    .y(_02449_)
  );
  al_nand3 _07738_ (
    .a(_00448_),
    .b(_02448_),
    .c(_02449_),
    .y(_02450_)
  );
  al_aoi21 _07739_ (
    .a(TM0),
    .b(\DFF_955.Q ),
    .c(TM1),
    .y(_02451_)
  );
  al_nand2 _07740_ (
    .a(_02451_),
    .b(_02450_),
    .y(_02452_)
  );
  al_aoi21ttf _07741_ (
    .a(TM0),
    .b(\DFF_772.Q ),
    .c(TM1),
    .y(_02453_)
  );
  al_and2 _07742_ (
    .a(_02453_),
    .b(_01961_),
    .y(_02454_)
  );
  al_nor3fft _07743_ (
    .a(RESET),
    .b(_02452_),
    .c(_02454_),
    .y(\DFF_804.D )
  );
  al_or2 _07744_ (
    .a(TM1),
    .b(\DFF_1061.Q ),
    .y(_02455_)
  );
  al_nand2 _07745_ (
    .a(TM1),
    .b(\DFF_1061.Q ),
    .y(_02456_)
  );
  al_nand3 _07746_ (
    .a(\DFF_1093.Q ),
    .b(_02455_),
    .c(_02456_),
    .y(_02457_)
  );
  al_nand2ft _07747_ (
    .a(TM1),
    .b(\DFF_1061.Q ),
    .y(_02458_)
  );
  al_and2ft _07748_ (
    .a(\DFF_1061.Q ),
    .b(TM1),
    .y(_02459_)
  );
  al_and3fft _07749_ (
    .a(\DFF_1093.Q ),
    .b(_02459_),
    .c(_02458_),
    .y(_02460_)
  );
  al_and2ft _07750_ (
    .a(\DFF_1029.Q ),
    .b(\DFF_997.Q ),
    .y(_02461_)
  );
  al_nand2ft _07751_ (
    .a(\DFF_997.Q ),
    .b(\DFF_1029.Q ),
    .y(_02462_)
  );
  al_nand2ft _07752_ (
    .a(_02461_),
    .b(_02462_),
    .y(_02463_)
  );
  al_oai21ftf _07753_ (
    .a(_02457_),
    .b(_02460_),
    .c(_02463_),
    .y(_02464_)
  );
  al_nand3ftt _07754_ (
    .a(_02460_),
    .b(_02457_),
    .c(_02463_),
    .y(_02465_)
  );
  al_nand3 _07755_ (
    .a(_00448_),
    .b(_02464_),
    .c(_02465_),
    .y(_02466_)
  );
  al_aoi21 _07756_ (
    .a(TM0),
    .b(\DFF_954.Q ),
    .c(TM1),
    .y(_02467_)
  );
  al_nand2 _07757_ (
    .a(_02467_),
    .b(_02466_),
    .y(_02468_)
  );
  al_aoi21ttf _07758_ (
    .a(TM0),
    .b(\DFF_773.Q ),
    .c(TM1),
    .y(_02469_)
  );
  al_and2 _07759_ (
    .a(_02469_),
    .b(_01977_),
    .y(_02470_)
  );
  al_nor3fft _07760_ (
    .a(RESET),
    .b(_02468_),
    .c(_02470_),
    .y(\DFF_805.D )
  );
  al_or2 _07761_ (
    .a(TM1),
    .b(\DFF_1062.Q ),
    .y(_02471_)
  );
  al_nand2 _07762_ (
    .a(TM1),
    .b(\DFF_1062.Q ),
    .y(_02472_)
  );
  al_nand3 _07763_ (
    .a(\DFF_1094.Q ),
    .b(_02471_),
    .c(_02472_),
    .y(_02473_)
  );
  al_nand2ft _07764_ (
    .a(TM1),
    .b(\DFF_1062.Q ),
    .y(_02474_)
  );
  al_and2ft _07765_ (
    .a(\DFF_1062.Q ),
    .b(TM1),
    .y(_02475_)
  );
  al_and3fft _07766_ (
    .a(\DFF_1094.Q ),
    .b(_02475_),
    .c(_02474_),
    .y(_02476_)
  );
  al_and2ft _07767_ (
    .a(\DFF_1030.Q ),
    .b(\DFF_998.Q ),
    .y(_02477_)
  );
  al_nand2ft _07768_ (
    .a(\DFF_998.Q ),
    .b(\DFF_1030.Q ),
    .y(_02478_)
  );
  al_nand2ft _07769_ (
    .a(_02477_),
    .b(_02478_),
    .y(_02479_)
  );
  al_oai21ftf _07770_ (
    .a(_02473_),
    .b(_02476_),
    .c(_02479_),
    .y(_02480_)
  );
  al_nand3ftt _07771_ (
    .a(_02476_),
    .b(_02473_),
    .c(_02479_),
    .y(_02481_)
  );
  al_nand3 _07772_ (
    .a(_00448_),
    .b(_02480_),
    .c(_02481_),
    .y(_02482_)
  );
  al_aoi21 _07773_ (
    .a(TM0),
    .b(\DFF_953.Q ),
    .c(TM1),
    .y(_02483_)
  );
  al_nand2 _07774_ (
    .a(_02483_),
    .b(_02482_),
    .y(_02484_)
  );
  al_aoi21ttf _07775_ (
    .a(TM0),
    .b(\DFF_774.Q ),
    .c(TM1),
    .y(_02485_)
  );
  al_and2 _07776_ (
    .a(_02485_),
    .b(_01993_),
    .y(_02486_)
  );
  al_nor3fft _07777_ (
    .a(RESET),
    .b(_02484_),
    .c(_02486_),
    .y(\DFF_806.D )
  );
  al_or2 _07778_ (
    .a(TM1),
    .b(\DFF_1063.Q ),
    .y(_02487_)
  );
  al_nand2 _07779_ (
    .a(TM1),
    .b(\DFF_1063.Q ),
    .y(_02488_)
  );
  al_nand3 _07780_ (
    .a(\DFF_1095.Q ),
    .b(_02487_),
    .c(_02488_),
    .y(_02489_)
  );
  al_nand2ft _07781_ (
    .a(TM1),
    .b(\DFF_1063.Q ),
    .y(_02490_)
  );
  al_and2ft _07782_ (
    .a(\DFF_1063.Q ),
    .b(TM1),
    .y(_02491_)
  );
  al_and3fft _07783_ (
    .a(\DFF_1095.Q ),
    .b(_02491_),
    .c(_02490_),
    .y(_02492_)
  );
  al_and2ft _07784_ (
    .a(\DFF_1031.Q ),
    .b(\DFF_999.Q ),
    .y(_02493_)
  );
  al_nand2ft _07785_ (
    .a(\DFF_999.Q ),
    .b(\DFF_1031.Q ),
    .y(_02494_)
  );
  al_nand2ft _07786_ (
    .a(_02493_),
    .b(_02494_),
    .y(_02495_)
  );
  al_oai21ftf _07787_ (
    .a(_02489_),
    .b(_02492_),
    .c(_02495_),
    .y(_02496_)
  );
  al_nand3ftt _07788_ (
    .a(_02492_),
    .b(_02489_),
    .c(_02495_),
    .y(_02497_)
  );
  al_nand3 _07789_ (
    .a(_00448_),
    .b(_02496_),
    .c(_02497_),
    .y(_02498_)
  );
  al_aoi21 _07790_ (
    .a(TM0),
    .b(\DFF_952.Q ),
    .c(TM1),
    .y(_02499_)
  );
  al_nand2 _07791_ (
    .a(_02499_),
    .b(_02498_),
    .y(_02500_)
  );
  al_aoi21ttf _07792_ (
    .a(TM0),
    .b(\DFF_775.Q ),
    .c(TM1),
    .y(_02501_)
  );
  al_and2 _07793_ (
    .a(_02501_),
    .b(_02009_),
    .y(_02502_)
  );
  al_nor3fft _07794_ (
    .a(RESET),
    .b(_02500_),
    .c(_02502_),
    .y(\DFF_807.D )
  );
  al_or2 _07795_ (
    .a(TM1),
    .b(\DFF_1064.Q ),
    .y(_02503_)
  );
  al_nand2 _07796_ (
    .a(TM1),
    .b(\DFF_1064.Q ),
    .y(_02504_)
  );
  al_nand3 _07797_ (
    .a(\DFF_1096.Q ),
    .b(_02503_),
    .c(_02504_),
    .y(_02505_)
  );
  al_nand2ft _07798_ (
    .a(TM1),
    .b(\DFF_1064.Q ),
    .y(_02506_)
  );
  al_and2ft _07799_ (
    .a(\DFF_1064.Q ),
    .b(TM1),
    .y(_02507_)
  );
  al_and3fft _07800_ (
    .a(\DFF_1096.Q ),
    .b(_02507_),
    .c(_02506_),
    .y(_02508_)
  );
  al_and2ft _07801_ (
    .a(\DFF_1032.Q ),
    .b(\DFF_1000.Q ),
    .y(_02509_)
  );
  al_nand2ft _07802_ (
    .a(\DFF_1000.Q ),
    .b(\DFF_1032.Q ),
    .y(_02510_)
  );
  al_nand2ft _07803_ (
    .a(_02509_),
    .b(_02510_),
    .y(_02511_)
  );
  al_oai21ftf _07804_ (
    .a(_02505_),
    .b(_02508_),
    .c(_02511_),
    .y(_02512_)
  );
  al_nand3ftt _07805_ (
    .a(_02508_),
    .b(_02505_),
    .c(_02511_),
    .y(_02513_)
  );
  al_nand3 _07806_ (
    .a(_00448_),
    .b(_02512_),
    .c(_02513_),
    .y(_02514_)
  );
  al_aoi21 _07807_ (
    .a(TM0),
    .b(\DFF_951.Q ),
    .c(TM1),
    .y(_02515_)
  );
  al_nand2 _07808_ (
    .a(_02515_),
    .b(_02514_),
    .y(_02516_)
  );
  al_aoi21ttf _07809_ (
    .a(TM0),
    .b(\DFF_776.Q ),
    .c(TM1),
    .y(_02517_)
  );
  al_and2 _07810_ (
    .a(_02517_),
    .b(_02025_),
    .y(_02518_)
  );
  al_nor3fft _07811_ (
    .a(RESET),
    .b(_02516_),
    .c(_02518_),
    .y(\DFF_808.D )
  );
  al_or2 _07812_ (
    .a(TM1),
    .b(\DFF_1065.Q ),
    .y(_02519_)
  );
  al_nand2 _07813_ (
    .a(TM1),
    .b(\DFF_1065.Q ),
    .y(_02520_)
  );
  al_nand3 _07814_ (
    .a(\DFF_1097.Q ),
    .b(_02519_),
    .c(_02520_),
    .y(_02521_)
  );
  al_nand2ft _07815_ (
    .a(TM1),
    .b(\DFF_1065.Q ),
    .y(_02522_)
  );
  al_and2ft _07816_ (
    .a(\DFF_1065.Q ),
    .b(TM1),
    .y(_02523_)
  );
  al_and3fft _07817_ (
    .a(\DFF_1097.Q ),
    .b(_02523_),
    .c(_02522_),
    .y(_02524_)
  );
  al_and2ft _07818_ (
    .a(\DFF_1033.Q ),
    .b(\DFF_1001.Q ),
    .y(_02525_)
  );
  al_nand2ft _07819_ (
    .a(\DFF_1001.Q ),
    .b(\DFF_1033.Q ),
    .y(_02526_)
  );
  al_nand2ft _07820_ (
    .a(_02525_),
    .b(_02526_),
    .y(_02527_)
  );
  al_oai21ftf _07821_ (
    .a(_02521_),
    .b(_02524_),
    .c(_02527_),
    .y(_02528_)
  );
  al_nand3ftt _07822_ (
    .a(_02524_),
    .b(_02521_),
    .c(_02527_),
    .y(_02529_)
  );
  al_nand3 _07823_ (
    .a(_00448_),
    .b(_02528_),
    .c(_02529_),
    .y(_02530_)
  );
  al_aoi21 _07824_ (
    .a(TM0),
    .b(\DFF_950.Q ),
    .c(TM1),
    .y(_02531_)
  );
  al_nand2 _07825_ (
    .a(_02531_),
    .b(_02530_),
    .y(_02532_)
  );
  al_aoi21ttf _07826_ (
    .a(TM0),
    .b(\DFF_777.Q ),
    .c(TM1),
    .y(_02533_)
  );
  al_and2 _07827_ (
    .a(_02533_),
    .b(_02041_),
    .y(_02534_)
  );
  al_nor3fft _07828_ (
    .a(RESET),
    .b(_02532_),
    .c(_02534_),
    .y(\DFF_809.D )
  );
  al_or2 _07829_ (
    .a(TM1),
    .b(\DFF_1066.Q ),
    .y(_02535_)
  );
  al_nand2 _07830_ (
    .a(TM1),
    .b(\DFF_1066.Q ),
    .y(_02536_)
  );
  al_nand3 _07831_ (
    .a(\DFF_1098.Q ),
    .b(_02535_),
    .c(_02536_),
    .y(_02537_)
  );
  al_nand2ft _07832_ (
    .a(TM1),
    .b(\DFF_1066.Q ),
    .y(_02538_)
  );
  al_and2ft _07833_ (
    .a(\DFF_1066.Q ),
    .b(TM1),
    .y(_02539_)
  );
  al_and3fft _07834_ (
    .a(\DFF_1098.Q ),
    .b(_02539_),
    .c(_02538_),
    .y(_02540_)
  );
  al_and2ft _07835_ (
    .a(\DFF_1034.Q ),
    .b(\DFF_1002.Q ),
    .y(_02541_)
  );
  al_nand2ft _07836_ (
    .a(\DFF_1002.Q ),
    .b(\DFF_1034.Q ),
    .y(_02542_)
  );
  al_nand2ft _07837_ (
    .a(_02541_),
    .b(_02542_),
    .y(_02543_)
  );
  al_oai21ftf _07838_ (
    .a(_02537_),
    .b(_02540_),
    .c(_02543_),
    .y(_02544_)
  );
  al_nand3ftt _07839_ (
    .a(_02540_),
    .b(_02537_),
    .c(_02543_),
    .y(_02545_)
  );
  al_nand3 _07840_ (
    .a(_00448_),
    .b(_02544_),
    .c(_02545_),
    .y(_02546_)
  );
  al_aoi21 _07841_ (
    .a(TM0),
    .b(\DFF_949.Q ),
    .c(TM1),
    .y(_02547_)
  );
  al_nand2 _07842_ (
    .a(_02547_),
    .b(_02546_),
    .y(_02548_)
  );
  al_aoi21ttf _07843_ (
    .a(TM0),
    .b(\DFF_778.Q ),
    .c(TM1),
    .y(_02549_)
  );
  al_and2 _07844_ (
    .a(_02549_),
    .b(_02057_),
    .y(_02550_)
  );
  al_nor3fft _07845_ (
    .a(RESET),
    .b(_02548_),
    .c(_02550_),
    .y(\DFF_810.D )
  );
  al_or2 _07846_ (
    .a(TM1),
    .b(\DFF_1067.Q ),
    .y(_02551_)
  );
  al_nand2 _07847_ (
    .a(TM1),
    .b(\DFF_1067.Q ),
    .y(_02552_)
  );
  al_nand3 _07848_ (
    .a(\DFF_1099.Q ),
    .b(_02551_),
    .c(_02552_),
    .y(_02553_)
  );
  al_nand2ft _07849_ (
    .a(TM1),
    .b(\DFF_1067.Q ),
    .y(_02554_)
  );
  al_and2ft _07850_ (
    .a(\DFF_1067.Q ),
    .b(TM1),
    .y(_02555_)
  );
  al_and3fft _07851_ (
    .a(\DFF_1099.Q ),
    .b(_02555_),
    .c(_02554_),
    .y(_02556_)
  );
  al_and2ft _07852_ (
    .a(\DFF_1035.Q ),
    .b(\DFF_1003.Q ),
    .y(_02557_)
  );
  al_nand2ft _07853_ (
    .a(\DFF_1003.Q ),
    .b(\DFF_1035.Q ),
    .y(_02558_)
  );
  al_nand2ft _07854_ (
    .a(_02557_),
    .b(_02558_),
    .y(_02559_)
  );
  al_oai21ftf _07855_ (
    .a(_02553_),
    .b(_02556_),
    .c(_02559_),
    .y(_02560_)
  );
  al_nand3ftt _07856_ (
    .a(_02556_),
    .b(_02553_),
    .c(_02559_),
    .y(_02561_)
  );
  al_nand3 _07857_ (
    .a(_00448_),
    .b(_02560_),
    .c(_02561_),
    .y(_02562_)
  );
  al_aoi21 _07858_ (
    .a(TM0),
    .b(\DFF_948.Q ),
    .c(TM1),
    .y(_02563_)
  );
  al_nand2 _07859_ (
    .a(_02563_),
    .b(_02562_),
    .y(_02564_)
  );
  al_aoi21ttf _07860_ (
    .a(TM0),
    .b(\DFF_779.Q ),
    .c(TM1),
    .y(_02565_)
  );
  al_and2 _07861_ (
    .a(_02565_),
    .b(_02073_),
    .y(_02566_)
  );
  al_nor3fft _07862_ (
    .a(RESET),
    .b(_02564_),
    .c(_02566_),
    .y(\DFF_811.D )
  );
  al_or2 _07863_ (
    .a(TM1),
    .b(\DFF_1068.Q ),
    .y(_02567_)
  );
  al_nand2 _07864_ (
    .a(TM1),
    .b(\DFF_1068.Q ),
    .y(_02568_)
  );
  al_nand3 _07865_ (
    .a(\DFF_1100.Q ),
    .b(_02567_),
    .c(_02568_),
    .y(_02569_)
  );
  al_nand2ft _07866_ (
    .a(TM1),
    .b(\DFF_1068.Q ),
    .y(_02570_)
  );
  al_and2ft _07867_ (
    .a(\DFF_1068.Q ),
    .b(TM1),
    .y(_02571_)
  );
  al_and3fft _07868_ (
    .a(\DFF_1100.Q ),
    .b(_02571_),
    .c(_02570_),
    .y(_02572_)
  );
  al_and2ft _07869_ (
    .a(\DFF_1036.Q ),
    .b(\DFF_1004.Q ),
    .y(_02573_)
  );
  al_nand2ft _07870_ (
    .a(\DFF_1004.Q ),
    .b(\DFF_1036.Q ),
    .y(_02574_)
  );
  al_nand2ft _07871_ (
    .a(_02573_),
    .b(_02574_),
    .y(_02575_)
  );
  al_oai21ftf _07872_ (
    .a(_02569_),
    .b(_02572_),
    .c(_02575_),
    .y(_02576_)
  );
  al_nand3ftt _07873_ (
    .a(_02572_),
    .b(_02569_),
    .c(_02575_),
    .y(_02577_)
  );
  al_nand3 _07874_ (
    .a(_00448_),
    .b(_02576_),
    .c(_02577_),
    .y(_02578_)
  );
  al_aoi21 _07875_ (
    .a(TM0),
    .b(\DFF_947.Q ),
    .c(TM1),
    .y(_02579_)
  );
  al_nand2 _07876_ (
    .a(_02579_),
    .b(_02578_),
    .y(_02580_)
  );
  al_aoi21ttf _07877_ (
    .a(TM0),
    .b(\DFF_780.Q ),
    .c(TM1),
    .y(_02581_)
  );
  al_and2 _07878_ (
    .a(_02581_),
    .b(_02089_),
    .y(_02582_)
  );
  al_nor3fft _07879_ (
    .a(RESET),
    .b(_02580_),
    .c(_02582_),
    .y(\DFF_812.D )
  );
  al_or2 _07880_ (
    .a(TM1),
    .b(\DFF_1069.Q ),
    .y(_02583_)
  );
  al_nand2 _07881_ (
    .a(TM1),
    .b(\DFF_1069.Q ),
    .y(_02584_)
  );
  al_nand3 _07882_ (
    .a(\DFF_1101.Q ),
    .b(_02583_),
    .c(_02584_),
    .y(_02585_)
  );
  al_nand2ft _07883_ (
    .a(TM1),
    .b(\DFF_1069.Q ),
    .y(_02586_)
  );
  al_and2ft _07884_ (
    .a(\DFF_1069.Q ),
    .b(TM1),
    .y(_02587_)
  );
  al_and3fft _07885_ (
    .a(\DFF_1101.Q ),
    .b(_02587_),
    .c(_02586_),
    .y(_02588_)
  );
  al_and2ft _07886_ (
    .a(\DFF_1037.Q ),
    .b(\DFF_1005.Q ),
    .y(_02589_)
  );
  al_nand2ft _07887_ (
    .a(\DFF_1005.Q ),
    .b(\DFF_1037.Q ),
    .y(_02590_)
  );
  al_nand2ft _07888_ (
    .a(_02589_),
    .b(_02590_),
    .y(_02591_)
  );
  al_oai21ftf _07889_ (
    .a(_02585_),
    .b(_02588_),
    .c(_02591_),
    .y(_02592_)
  );
  al_nand3ftt _07890_ (
    .a(_02588_),
    .b(_02585_),
    .c(_02591_),
    .y(_02593_)
  );
  al_nand3 _07891_ (
    .a(_00448_),
    .b(_02592_),
    .c(_02593_),
    .y(_02594_)
  );
  al_aoi21 _07892_ (
    .a(TM0),
    .b(\DFF_946.Q ),
    .c(TM1),
    .y(_02595_)
  );
  al_nand2 _07893_ (
    .a(_02595_),
    .b(_02594_),
    .y(_02596_)
  );
  al_aoi21ttf _07894_ (
    .a(TM0),
    .b(\DFF_781.Q ),
    .c(TM1),
    .y(_02597_)
  );
  al_and2 _07895_ (
    .a(_02597_),
    .b(_02105_),
    .y(_02598_)
  );
  al_nor3fft _07896_ (
    .a(RESET),
    .b(_02596_),
    .c(_02598_),
    .y(\DFF_813.D )
  );
  al_or2 _07897_ (
    .a(TM1),
    .b(\DFF_1070.Q ),
    .y(_02599_)
  );
  al_nand2 _07898_ (
    .a(TM1),
    .b(\DFF_1070.Q ),
    .y(_02600_)
  );
  al_nand3 _07899_ (
    .a(\DFF_1102.Q ),
    .b(_02599_),
    .c(_02600_),
    .y(_02601_)
  );
  al_nand2ft _07900_ (
    .a(TM1),
    .b(\DFF_1070.Q ),
    .y(_02602_)
  );
  al_and2ft _07901_ (
    .a(\DFF_1070.Q ),
    .b(TM1),
    .y(_02603_)
  );
  al_and3fft _07902_ (
    .a(\DFF_1102.Q ),
    .b(_02603_),
    .c(_02602_),
    .y(_02604_)
  );
  al_and2ft _07903_ (
    .a(\DFF_1038.Q ),
    .b(\DFF_1006.Q ),
    .y(_02605_)
  );
  al_nand2ft _07904_ (
    .a(\DFF_1006.Q ),
    .b(\DFF_1038.Q ),
    .y(_02606_)
  );
  al_nand2ft _07905_ (
    .a(_02605_),
    .b(_02606_),
    .y(_02607_)
  );
  al_oai21ftf _07906_ (
    .a(_02601_),
    .b(_02604_),
    .c(_02607_),
    .y(_02608_)
  );
  al_nand3ftt _07907_ (
    .a(_02604_),
    .b(_02601_),
    .c(_02607_),
    .y(_02609_)
  );
  al_nand3 _07908_ (
    .a(_00448_),
    .b(_02608_),
    .c(_02609_),
    .y(_02610_)
  );
  al_aoi21 _07909_ (
    .a(TM0),
    .b(\DFF_945.Q ),
    .c(TM1),
    .y(_02611_)
  );
  al_nand2 _07910_ (
    .a(_02611_),
    .b(_02610_),
    .y(_02612_)
  );
  al_aoi21ttf _07911_ (
    .a(TM0),
    .b(\DFF_782.Q ),
    .c(TM1),
    .y(_02613_)
  );
  al_and2 _07912_ (
    .a(_02613_),
    .b(_02121_),
    .y(_02614_)
  );
  al_nor3fft _07913_ (
    .a(RESET),
    .b(_02612_),
    .c(_02614_),
    .y(\DFF_814.D )
  );
  al_or2 _07914_ (
    .a(TM1),
    .b(\DFF_1071.Q ),
    .y(_02615_)
  );
  al_nand2 _07915_ (
    .a(TM1),
    .b(\DFF_1071.Q ),
    .y(_02616_)
  );
  al_nand3 _07916_ (
    .a(\DFF_1103.Q ),
    .b(_02615_),
    .c(_02616_),
    .y(_02617_)
  );
  al_nand2ft _07917_ (
    .a(TM1),
    .b(\DFF_1071.Q ),
    .y(_02618_)
  );
  al_and2ft _07918_ (
    .a(\DFF_1071.Q ),
    .b(TM1),
    .y(_02619_)
  );
  al_and3fft _07919_ (
    .a(\DFF_1103.Q ),
    .b(_02619_),
    .c(_02618_),
    .y(_02620_)
  );
  al_and2ft _07920_ (
    .a(\DFF_1039.Q ),
    .b(\DFF_1007.Q ),
    .y(_02621_)
  );
  al_nand2ft _07921_ (
    .a(\DFF_1007.Q ),
    .b(\DFF_1039.Q ),
    .y(_02622_)
  );
  al_nand2ft _07922_ (
    .a(_02621_),
    .b(_02622_),
    .y(_02623_)
  );
  al_oai21ftf _07923_ (
    .a(_02617_),
    .b(_02620_),
    .c(_02623_),
    .y(_02624_)
  );
  al_nand3ftt _07924_ (
    .a(_02620_),
    .b(_02617_),
    .c(_02623_),
    .y(_02625_)
  );
  al_nand3 _07925_ (
    .a(_00448_),
    .b(_02624_),
    .c(_02625_),
    .y(_02626_)
  );
  al_aoi21 _07926_ (
    .a(TM0),
    .b(\DFF_944.Q ),
    .c(TM1),
    .y(_02627_)
  );
  al_nand2 _07927_ (
    .a(_02627_),
    .b(_02626_),
    .y(_02628_)
  );
  al_aoi21ttf _07928_ (
    .a(TM0),
    .b(\DFF_783.Q ),
    .c(TM1),
    .y(_02629_)
  );
  al_and2 _07929_ (
    .a(_02629_),
    .b(_02137_),
    .y(_02630_)
  );
  al_nor3fft _07930_ (
    .a(RESET),
    .b(_02628_),
    .c(_02630_),
    .y(\DFF_815.D )
  );
  al_nor2 _07931_ (
    .a(\DFF_1040.Q ),
    .b(\DFF_1072.Q ),
    .y(_02631_)
  );
  al_and2 _07932_ (
    .a(\DFF_1040.Q ),
    .b(\DFF_1072.Q ),
    .y(_02632_)
  );
  al_and2ft _07933_ (
    .a(\DFF_1008.Q ),
    .b(\DFF_1104.Q ),
    .y(_02633_)
  );
  al_nand2ft _07934_ (
    .a(\DFF_1104.Q ),
    .b(\DFF_1008.Q ),
    .y(_02634_)
  );
  al_nand2ft _07935_ (
    .a(_02633_),
    .b(_02634_),
    .y(_02635_)
  );
  al_oa21ttf _07936_ (
    .a(_02631_),
    .b(_02632_),
    .c(_02635_),
    .y(_02636_)
  );
  al_nand3fft _07937_ (
    .a(_02631_),
    .b(_02632_),
    .c(_02635_),
    .y(_02637_)
  );
  al_and3fft _07938_ (
    .a(TM0),
    .b(_02636_),
    .c(_02637_),
    .y(_02638_)
  );
  al_nand2 _07939_ (
    .a(TM0),
    .b(\DFF_943.Q ),
    .y(_02639_)
  );
  al_or3fft _07940_ (
    .a(_01652_),
    .b(_02639_),
    .c(_02638_),
    .y(_02640_)
  );
  al_and2 _07941_ (
    .a(TM0),
    .b(\DFF_784.Q ),
    .y(_02641_)
  );
  al_and3fft _07942_ (
    .a(_02641_),
    .b(_02149_),
    .c(TM1),
    .y(_02642_)
  );
  al_nor3fft _07943_ (
    .a(RESET),
    .b(_02640_),
    .c(_02642_),
    .y(\DFF_816.D )
  );
  al_nor2 _07944_ (
    .a(\DFF_1041.Q ),
    .b(\DFF_1073.Q ),
    .y(_02643_)
  );
  al_and2 _07945_ (
    .a(\DFF_1041.Q ),
    .b(\DFF_1073.Q ),
    .y(_02644_)
  );
  al_and2ft _07946_ (
    .a(\DFF_1009.Q ),
    .b(\DFF_1105.Q ),
    .y(_02645_)
  );
  al_nand2ft _07947_ (
    .a(\DFF_1105.Q ),
    .b(\DFF_1009.Q ),
    .y(_02646_)
  );
  al_nand2ft _07948_ (
    .a(_02645_),
    .b(_02646_),
    .y(_02647_)
  );
  al_oa21ttf _07949_ (
    .a(_02643_),
    .b(_02644_),
    .c(_02647_),
    .y(_02648_)
  );
  al_nand3fft _07950_ (
    .a(_02643_),
    .b(_02644_),
    .c(_02647_),
    .y(_02649_)
  );
  al_and3fft _07951_ (
    .a(TM0),
    .b(_02648_),
    .c(_02649_),
    .y(_02650_)
  );
  al_nand2 _07952_ (
    .a(TM0),
    .b(\DFF_942.Q ),
    .y(_02651_)
  );
  al_or3fft _07953_ (
    .a(_01652_),
    .b(_02651_),
    .c(_02650_),
    .y(_02652_)
  );
  al_and2 _07954_ (
    .a(TM0),
    .b(\DFF_785.Q ),
    .y(_02653_)
  );
  al_and3fft _07955_ (
    .a(_02653_),
    .b(_02161_),
    .c(TM1),
    .y(_02654_)
  );
  al_nor3fft _07956_ (
    .a(RESET),
    .b(_02652_),
    .c(_02654_),
    .y(\DFF_817.D )
  );
  al_nor2 _07957_ (
    .a(\DFF_1042.Q ),
    .b(\DFF_1074.Q ),
    .y(_02655_)
  );
  al_and2 _07958_ (
    .a(\DFF_1042.Q ),
    .b(\DFF_1074.Q ),
    .y(_02656_)
  );
  al_and2ft _07959_ (
    .a(\DFF_1010.Q ),
    .b(\DFF_1106.Q ),
    .y(_02657_)
  );
  al_nand2ft _07960_ (
    .a(\DFF_1106.Q ),
    .b(\DFF_1010.Q ),
    .y(_02658_)
  );
  al_nand2ft _07961_ (
    .a(_02657_),
    .b(_02658_),
    .y(_02659_)
  );
  al_oa21ttf _07962_ (
    .a(_02655_),
    .b(_02656_),
    .c(_02659_),
    .y(_02660_)
  );
  al_nand3fft _07963_ (
    .a(_02655_),
    .b(_02656_),
    .c(_02659_),
    .y(_02661_)
  );
  al_and3fft _07964_ (
    .a(TM0),
    .b(_02660_),
    .c(_02661_),
    .y(_02662_)
  );
  al_nand2 _07965_ (
    .a(TM0),
    .b(\DFF_941.Q ),
    .y(_02663_)
  );
  al_or3fft _07966_ (
    .a(_01652_),
    .b(_02663_),
    .c(_02662_),
    .y(_02664_)
  );
  al_and2 _07967_ (
    .a(TM0),
    .b(\DFF_786.Q ),
    .y(_02665_)
  );
  al_and3fft _07968_ (
    .a(_02665_),
    .b(_02173_),
    .c(TM1),
    .y(_02666_)
  );
  al_nor3fft _07969_ (
    .a(RESET),
    .b(_02664_),
    .c(_02666_),
    .y(\DFF_818.D )
  );
  al_nor2 _07970_ (
    .a(\DFF_1043.Q ),
    .b(\DFF_1075.Q ),
    .y(_02667_)
  );
  al_and2 _07971_ (
    .a(\DFF_1043.Q ),
    .b(\DFF_1075.Q ),
    .y(_02668_)
  );
  al_and2ft _07972_ (
    .a(\DFF_1011.Q ),
    .b(\DFF_1107.Q ),
    .y(_02669_)
  );
  al_nand2ft _07973_ (
    .a(\DFF_1107.Q ),
    .b(\DFF_1011.Q ),
    .y(_02670_)
  );
  al_nand2ft _07974_ (
    .a(_02669_),
    .b(_02670_),
    .y(_02671_)
  );
  al_oa21ttf _07975_ (
    .a(_02667_),
    .b(_02668_),
    .c(_02671_),
    .y(_02672_)
  );
  al_nand3fft _07976_ (
    .a(_02667_),
    .b(_02668_),
    .c(_02671_),
    .y(_02673_)
  );
  al_and3fft _07977_ (
    .a(TM0),
    .b(_02672_),
    .c(_02673_),
    .y(_02674_)
  );
  al_nand2 _07978_ (
    .a(TM0),
    .b(\DFF_940.Q ),
    .y(_02675_)
  );
  al_or3fft _07979_ (
    .a(_01652_),
    .b(_02675_),
    .c(_02674_),
    .y(_02676_)
  );
  al_and2 _07980_ (
    .a(TM0),
    .b(\DFF_787.Q ),
    .y(_02677_)
  );
  al_and3fft _07981_ (
    .a(_02677_),
    .b(_02185_),
    .c(TM1),
    .y(_02678_)
  );
  al_nor3fft _07982_ (
    .a(RESET),
    .b(_02676_),
    .c(_02678_),
    .y(\DFF_819.D )
  );
  al_nor2 _07983_ (
    .a(\DFF_1044.Q ),
    .b(\DFF_1076.Q ),
    .y(_02679_)
  );
  al_and2 _07984_ (
    .a(\DFF_1044.Q ),
    .b(\DFF_1076.Q ),
    .y(_02680_)
  );
  al_and2ft _07985_ (
    .a(\DFF_1012.Q ),
    .b(\DFF_1108.Q ),
    .y(_02681_)
  );
  al_nand2ft _07986_ (
    .a(\DFF_1108.Q ),
    .b(\DFF_1012.Q ),
    .y(_02682_)
  );
  al_nand2ft _07987_ (
    .a(_02681_),
    .b(_02682_),
    .y(_02683_)
  );
  al_oa21ttf _07988_ (
    .a(_02679_),
    .b(_02680_),
    .c(_02683_),
    .y(_02684_)
  );
  al_nand3fft _07989_ (
    .a(_02679_),
    .b(_02680_),
    .c(_02683_),
    .y(_02685_)
  );
  al_and3fft _07990_ (
    .a(TM0),
    .b(_02684_),
    .c(_02685_),
    .y(_02686_)
  );
  al_nand2 _07991_ (
    .a(TM0),
    .b(\DFF_939.Q ),
    .y(_02687_)
  );
  al_or3fft _07992_ (
    .a(_01652_),
    .b(_02687_),
    .c(_02686_),
    .y(_02688_)
  );
  al_and2 _07993_ (
    .a(TM0),
    .b(\DFF_788.Q ),
    .y(_02689_)
  );
  al_and3fft _07994_ (
    .a(_02689_),
    .b(_02197_),
    .c(TM1),
    .y(_02690_)
  );
  al_nor3fft _07995_ (
    .a(RESET),
    .b(_02688_),
    .c(_02690_),
    .y(\DFF_820.D )
  );
  al_nor2 _07996_ (
    .a(\DFF_1045.Q ),
    .b(\DFF_1077.Q ),
    .y(_02691_)
  );
  al_and2 _07997_ (
    .a(\DFF_1045.Q ),
    .b(\DFF_1077.Q ),
    .y(_02692_)
  );
  al_and2ft _07998_ (
    .a(\DFF_1013.Q ),
    .b(\DFF_1109.Q ),
    .y(_02693_)
  );
  al_nand2ft _07999_ (
    .a(\DFF_1109.Q ),
    .b(\DFF_1013.Q ),
    .y(_02694_)
  );
  al_nand2ft _08000_ (
    .a(_02693_),
    .b(_02694_),
    .y(_02695_)
  );
  al_oa21ttf _08001_ (
    .a(_02691_),
    .b(_02692_),
    .c(_02695_),
    .y(_02696_)
  );
  al_nand3fft _08002_ (
    .a(_02691_),
    .b(_02692_),
    .c(_02695_),
    .y(_02697_)
  );
  al_and3fft _08003_ (
    .a(TM0),
    .b(_02696_),
    .c(_02697_),
    .y(_02698_)
  );
  al_nand2 _08004_ (
    .a(TM0),
    .b(\DFF_938.Q ),
    .y(_02699_)
  );
  al_or3fft _08005_ (
    .a(_01652_),
    .b(_02699_),
    .c(_02698_),
    .y(_02700_)
  );
  al_and2 _08006_ (
    .a(TM0),
    .b(\DFF_789.Q ),
    .y(_02701_)
  );
  al_and3fft _08007_ (
    .a(_02701_),
    .b(_02209_),
    .c(TM1),
    .y(_02702_)
  );
  al_nor3fft _08008_ (
    .a(RESET),
    .b(_02700_),
    .c(_02702_),
    .y(\DFF_821.D )
  );
  al_nor2 _08009_ (
    .a(\DFF_1046.Q ),
    .b(\DFF_1078.Q ),
    .y(_02703_)
  );
  al_and2 _08010_ (
    .a(\DFF_1046.Q ),
    .b(\DFF_1078.Q ),
    .y(_02704_)
  );
  al_and2ft _08011_ (
    .a(\DFF_1014.Q ),
    .b(\DFF_1110.Q ),
    .y(_02705_)
  );
  al_nand2ft _08012_ (
    .a(\DFF_1110.Q ),
    .b(\DFF_1014.Q ),
    .y(_02706_)
  );
  al_nand2ft _08013_ (
    .a(_02705_),
    .b(_02706_),
    .y(_02707_)
  );
  al_oa21ttf _08014_ (
    .a(_02703_),
    .b(_02704_),
    .c(_02707_),
    .y(_02708_)
  );
  al_nand3fft _08015_ (
    .a(_02703_),
    .b(_02704_),
    .c(_02707_),
    .y(_02709_)
  );
  al_and3fft _08016_ (
    .a(TM0),
    .b(_02708_),
    .c(_02709_),
    .y(_02710_)
  );
  al_nand2 _08017_ (
    .a(TM0),
    .b(\DFF_937.Q ),
    .y(_02711_)
  );
  al_or3fft _08018_ (
    .a(_01652_),
    .b(_02711_),
    .c(_02710_),
    .y(_02712_)
  );
  al_and2 _08019_ (
    .a(TM0),
    .b(\DFF_790.Q ),
    .y(_02713_)
  );
  al_and3fft _08020_ (
    .a(_02713_),
    .b(_02221_),
    .c(TM1),
    .y(_02714_)
  );
  al_nor3fft _08021_ (
    .a(RESET),
    .b(_02712_),
    .c(_02714_),
    .y(\DFF_822.D )
  );
  al_nor2 _08022_ (
    .a(\DFF_1047.Q ),
    .b(\DFF_1079.Q ),
    .y(_02715_)
  );
  al_and2 _08023_ (
    .a(\DFF_1047.Q ),
    .b(\DFF_1079.Q ),
    .y(_02716_)
  );
  al_and2ft _08024_ (
    .a(\DFF_1015.Q ),
    .b(\DFF_1111.Q ),
    .y(_02717_)
  );
  al_nand2ft _08025_ (
    .a(\DFF_1111.Q ),
    .b(\DFF_1015.Q ),
    .y(_02718_)
  );
  al_nand2ft _08026_ (
    .a(_02717_),
    .b(_02718_),
    .y(_02719_)
  );
  al_oa21ttf _08027_ (
    .a(_02715_),
    .b(_02716_),
    .c(_02719_),
    .y(_02720_)
  );
  al_nand3fft _08028_ (
    .a(_02715_),
    .b(_02716_),
    .c(_02719_),
    .y(_02721_)
  );
  al_and3fft _08029_ (
    .a(TM0),
    .b(_02720_),
    .c(_02721_),
    .y(_02722_)
  );
  al_nand2 _08030_ (
    .a(TM0),
    .b(\DFF_936.Q ),
    .y(_02723_)
  );
  al_or3fft _08031_ (
    .a(_01652_),
    .b(_02723_),
    .c(_02722_),
    .y(_02724_)
  );
  al_and2 _08032_ (
    .a(TM0),
    .b(\DFF_791.Q ),
    .y(_02725_)
  );
  al_and3fft _08033_ (
    .a(_02725_),
    .b(_02233_),
    .c(TM1),
    .y(_02726_)
  );
  al_nor3fft _08034_ (
    .a(RESET),
    .b(_02724_),
    .c(_02726_),
    .y(\DFF_823.D )
  );
  al_nor2 _08035_ (
    .a(\DFF_1048.Q ),
    .b(\DFF_1080.Q ),
    .y(_02727_)
  );
  al_and2 _08036_ (
    .a(\DFF_1048.Q ),
    .b(\DFF_1080.Q ),
    .y(_02728_)
  );
  al_and2ft _08037_ (
    .a(\DFF_1016.Q ),
    .b(\DFF_1112.Q ),
    .y(_02729_)
  );
  al_nand2ft _08038_ (
    .a(\DFF_1112.Q ),
    .b(\DFF_1016.Q ),
    .y(_02730_)
  );
  al_nand2ft _08039_ (
    .a(_02729_),
    .b(_02730_),
    .y(_02731_)
  );
  al_oa21ttf _08040_ (
    .a(_02727_),
    .b(_02728_),
    .c(_02731_),
    .y(_02732_)
  );
  al_nand3fft _08041_ (
    .a(_02727_),
    .b(_02728_),
    .c(_02731_),
    .y(_02733_)
  );
  al_and3fft _08042_ (
    .a(TM0),
    .b(_02732_),
    .c(_02733_),
    .y(_02734_)
  );
  al_nand2 _08043_ (
    .a(TM0),
    .b(\DFF_935.Q ),
    .y(_02735_)
  );
  al_or3fft _08044_ (
    .a(_01652_),
    .b(_02735_),
    .c(_02734_),
    .y(_02736_)
  );
  al_and2 _08045_ (
    .a(TM0),
    .b(\DFF_792.Q ),
    .y(_02737_)
  );
  al_and3fft _08046_ (
    .a(_02737_),
    .b(_02245_),
    .c(TM1),
    .y(_02738_)
  );
  al_nor3fft _08047_ (
    .a(RESET),
    .b(_02736_),
    .c(_02738_),
    .y(\DFF_824.D )
  );
  al_nor2 _08048_ (
    .a(\DFF_1049.Q ),
    .b(\DFF_1081.Q ),
    .y(_02739_)
  );
  al_and2 _08049_ (
    .a(\DFF_1049.Q ),
    .b(\DFF_1081.Q ),
    .y(_02740_)
  );
  al_and2ft _08050_ (
    .a(\DFF_1017.Q ),
    .b(\DFF_1113.Q ),
    .y(_02741_)
  );
  al_nand2ft _08051_ (
    .a(\DFF_1113.Q ),
    .b(\DFF_1017.Q ),
    .y(_02742_)
  );
  al_nand2ft _08052_ (
    .a(_02741_),
    .b(_02742_),
    .y(_02743_)
  );
  al_oa21ttf _08053_ (
    .a(_02739_),
    .b(_02740_),
    .c(_02743_),
    .y(_02744_)
  );
  al_nand3fft _08054_ (
    .a(_02739_),
    .b(_02740_),
    .c(_02743_),
    .y(_02745_)
  );
  al_and3fft _08055_ (
    .a(TM0),
    .b(_02744_),
    .c(_02745_),
    .y(_02746_)
  );
  al_nand2 _08056_ (
    .a(TM0),
    .b(\DFF_934.Q ),
    .y(_02747_)
  );
  al_or3fft _08057_ (
    .a(_01652_),
    .b(_02747_),
    .c(_02746_),
    .y(_02748_)
  );
  al_and2 _08058_ (
    .a(TM0),
    .b(\DFF_793.Q ),
    .y(_02749_)
  );
  al_and3fft _08059_ (
    .a(_02749_),
    .b(_02257_),
    .c(TM1),
    .y(_02750_)
  );
  al_nor3fft _08060_ (
    .a(RESET),
    .b(_02748_),
    .c(_02750_),
    .y(\DFF_825.D )
  );
  al_nor2 _08061_ (
    .a(\DFF_1050.Q ),
    .b(\DFF_1082.Q ),
    .y(_02751_)
  );
  al_and2 _08062_ (
    .a(\DFF_1050.Q ),
    .b(\DFF_1082.Q ),
    .y(_02752_)
  );
  al_and2ft _08063_ (
    .a(\DFF_1018.Q ),
    .b(\DFF_1114.Q ),
    .y(_02753_)
  );
  al_nand2ft _08064_ (
    .a(\DFF_1114.Q ),
    .b(\DFF_1018.Q ),
    .y(_02754_)
  );
  al_nand2ft _08065_ (
    .a(_02753_),
    .b(_02754_),
    .y(_02755_)
  );
  al_oa21ttf _08066_ (
    .a(_02751_),
    .b(_02752_),
    .c(_02755_),
    .y(_02756_)
  );
  al_nand3fft _08067_ (
    .a(_02751_),
    .b(_02752_),
    .c(_02755_),
    .y(_02757_)
  );
  al_and3fft _08068_ (
    .a(TM0),
    .b(_02756_),
    .c(_02757_),
    .y(_02758_)
  );
  al_nand2 _08069_ (
    .a(TM0),
    .b(\DFF_933.Q ),
    .y(_02759_)
  );
  al_or3fft _08070_ (
    .a(_01652_),
    .b(_02759_),
    .c(_02758_),
    .y(_02760_)
  );
  al_and2 _08071_ (
    .a(TM0),
    .b(\DFF_794.Q ),
    .y(_02761_)
  );
  al_and3fft _08072_ (
    .a(_02761_),
    .b(_02269_),
    .c(TM1),
    .y(_02762_)
  );
  al_nor3fft _08073_ (
    .a(RESET),
    .b(_02760_),
    .c(_02762_),
    .y(\DFF_826.D )
  );
  al_nor2 _08074_ (
    .a(\DFF_1051.Q ),
    .b(\DFF_1083.Q ),
    .y(_02763_)
  );
  al_and2 _08075_ (
    .a(\DFF_1051.Q ),
    .b(\DFF_1083.Q ),
    .y(_02764_)
  );
  al_and2ft _08076_ (
    .a(\DFF_1019.Q ),
    .b(\DFF_1115.Q ),
    .y(_02765_)
  );
  al_nand2ft _08077_ (
    .a(\DFF_1115.Q ),
    .b(\DFF_1019.Q ),
    .y(_02766_)
  );
  al_nand2ft _08078_ (
    .a(_02765_),
    .b(_02766_),
    .y(_02767_)
  );
  al_oa21ttf _08079_ (
    .a(_02763_),
    .b(_02764_),
    .c(_02767_),
    .y(_02768_)
  );
  al_nand3fft _08080_ (
    .a(_02763_),
    .b(_02764_),
    .c(_02767_),
    .y(_02769_)
  );
  al_and3fft _08081_ (
    .a(TM0),
    .b(_02768_),
    .c(_02769_),
    .y(_02770_)
  );
  al_nand2 _08082_ (
    .a(TM0),
    .b(\DFF_932.Q ),
    .y(_02771_)
  );
  al_or3fft _08083_ (
    .a(_01652_),
    .b(_02771_),
    .c(_02770_),
    .y(_02772_)
  );
  al_and2 _08084_ (
    .a(TM0),
    .b(\DFF_795.Q ),
    .y(_02773_)
  );
  al_and3fft _08085_ (
    .a(_02773_),
    .b(_02281_),
    .c(TM1),
    .y(_02774_)
  );
  al_nor3fft _08086_ (
    .a(RESET),
    .b(_02772_),
    .c(_02774_),
    .y(\DFF_827.D )
  );
  al_nor2 _08087_ (
    .a(\DFF_1052.Q ),
    .b(\DFF_1084.Q ),
    .y(_02775_)
  );
  al_and2 _08088_ (
    .a(\DFF_1052.Q ),
    .b(\DFF_1084.Q ),
    .y(_02776_)
  );
  al_and2ft _08089_ (
    .a(\DFF_1020.Q ),
    .b(\DFF_1116.Q ),
    .y(_02777_)
  );
  al_nand2ft _08090_ (
    .a(\DFF_1116.Q ),
    .b(\DFF_1020.Q ),
    .y(_02778_)
  );
  al_nand2ft _08091_ (
    .a(_02777_),
    .b(_02778_),
    .y(_02779_)
  );
  al_oa21ttf _08092_ (
    .a(_02775_),
    .b(_02776_),
    .c(_02779_),
    .y(_02780_)
  );
  al_nand3fft _08093_ (
    .a(_02775_),
    .b(_02776_),
    .c(_02779_),
    .y(_02781_)
  );
  al_and3fft _08094_ (
    .a(TM0),
    .b(_02780_),
    .c(_02781_),
    .y(_02782_)
  );
  al_nand2 _08095_ (
    .a(TM0),
    .b(\DFF_931.Q ),
    .y(_02783_)
  );
  al_or3fft _08096_ (
    .a(_01652_),
    .b(_02783_),
    .c(_02782_),
    .y(_02784_)
  );
  al_and2 _08097_ (
    .a(TM0),
    .b(\DFF_796.Q ),
    .y(_02785_)
  );
  al_and3fft _08098_ (
    .a(_02785_),
    .b(_02293_),
    .c(TM1),
    .y(_02786_)
  );
  al_nor3fft _08099_ (
    .a(RESET),
    .b(_02784_),
    .c(_02786_),
    .y(\DFF_828.D )
  );
  al_nor2 _08100_ (
    .a(\DFF_1053.Q ),
    .b(\DFF_1085.Q ),
    .y(_02787_)
  );
  al_and2 _08101_ (
    .a(\DFF_1053.Q ),
    .b(\DFF_1085.Q ),
    .y(_02788_)
  );
  al_and2ft _08102_ (
    .a(\DFF_1021.Q ),
    .b(\DFF_1117.Q ),
    .y(_02789_)
  );
  al_nand2ft _08103_ (
    .a(\DFF_1117.Q ),
    .b(\DFF_1021.Q ),
    .y(_02790_)
  );
  al_nand2ft _08104_ (
    .a(_02789_),
    .b(_02790_),
    .y(_02791_)
  );
  al_oa21ttf _08105_ (
    .a(_02787_),
    .b(_02788_),
    .c(_02791_),
    .y(_02792_)
  );
  al_nand3fft _08106_ (
    .a(_02787_),
    .b(_02788_),
    .c(_02791_),
    .y(_02793_)
  );
  al_and3fft _08107_ (
    .a(TM0),
    .b(_02792_),
    .c(_02793_),
    .y(_02794_)
  );
  al_nand2 _08108_ (
    .a(TM0),
    .b(\DFF_930.Q ),
    .y(_02795_)
  );
  al_or3fft _08109_ (
    .a(_01652_),
    .b(_02795_),
    .c(_02794_),
    .y(_02796_)
  );
  al_and2 _08110_ (
    .a(TM0),
    .b(\DFF_797.Q ),
    .y(_02797_)
  );
  al_and3fft _08111_ (
    .a(_02797_),
    .b(_02305_),
    .c(TM1),
    .y(_02798_)
  );
  al_nor3fft _08112_ (
    .a(RESET),
    .b(_02796_),
    .c(_02798_),
    .y(\DFF_829.D )
  );
  al_nor2 _08113_ (
    .a(\DFF_1054.Q ),
    .b(\DFF_1086.Q ),
    .y(_02799_)
  );
  al_and2 _08114_ (
    .a(\DFF_1054.Q ),
    .b(\DFF_1086.Q ),
    .y(_02800_)
  );
  al_and2ft _08115_ (
    .a(\DFF_1022.Q ),
    .b(\DFF_1118.Q ),
    .y(_02801_)
  );
  al_nand2ft _08116_ (
    .a(\DFF_1118.Q ),
    .b(\DFF_1022.Q ),
    .y(_02802_)
  );
  al_nand2ft _08117_ (
    .a(_02801_),
    .b(_02802_),
    .y(_02803_)
  );
  al_oa21ttf _08118_ (
    .a(_02799_),
    .b(_02800_),
    .c(_02803_),
    .y(_02804_)
  );
  al_nand3fft _08119_ (
    .a(_02799_),
    .b(_02800_),
    .c(_02803_),
    .y(_02805_)
  );
  al_and3fft _08120_ (
    .a(TM0),
    .b(_02804_),
    .c(_02805_),
    .y(_02806_)
  );
  al_nand2 _08121_ (
    .a(TM0),
    .b(\DFF_929.Q ),
    .y(_02807_)
  );
  al_or3fft _08122_ (
    .a(_01652_),
    .b(_02807_),
    .c(_02806_),
    .y(_02808_)
  );
  al_and2 _08123_ (
    .a(TM0),
    .b(\DFF_798.Q ),
    .y(_02809_)
  );
  al_and3fft _08124_ (
    .a(_02809_),
    .b(_02317_),
    .c(TM1),
    .y(_02810_)
  );
  al_nor3fft _08125_ (
    .a(RESET),
    .b(_02808_),
    .c(_02810_),
    .y(\DFF_830.D )
  );
  al_nor2 _08126_ (
    .a(\DFF_1055.Q ),
    .b(\DFF_1087.Q ),
    .y(_02811_)
  );
  al_and2 _08127_ (
    .a(\DFF_1055.Q ),
    .b(\DFF_1087.Q ),
    .y(_02812_)
  );
  al_and2ft _08128_ (
    .a(\DFF_1023.Q ),
    .b(\DFF_1119.Q ),
    .y(_02813_)
  );
  al_nand2ft _08129_ (
    .a(\DFF_1119.Q ),
    .b(\DFF_1023.Q ),
    .y(_02814_)
  );
  al_nand2ft _08130_ (
    .a(_02813_),
    .b(_02814_),
    .y(_02815_)
  );
  al_oa21ttf _08131_ (
    .a(_02811_),
    .b(_02812_),
    .c(_02815_),
    .y(_02816_)
  );
  al_nand3fft _08132_ (
    .a(_02811_),
    .b(_02812_),
    .c(_02815_),
    .y(_02817_)
  );
  al_and3fft _08133_ (
    .a(TM0),
    .b(_02816_),
    .c(_02817_),
    .y(_02818_)
  );
  al_nand2 _08134_ (
    .a(TM0),
    .b(\DFF_928.Q ),
    .y(_02819_)
  );
  al_or3fft _08135_ (
    .a(_01652_),
    .b(_02819_),
    .c(_02818_),
    .y(_02820_)
  );
  al_and2 _08136_ (
    .a(TM0),
    .b(\DFF_799.Q ),
    .y(_02821_)
  );
  al_and3fft _08137_ (
    .a(_02821_),
    .b(_02329_),
    .c(TM1),
    .y(_02822_)
  );
  al_nor3fft _08138_ (
    .a(RESET),
    .b(_02820_),
    .c(_02822_),
    .y(\DFF_831.D )
  );
  al_and2 _08139_ (
    .a(RESET),
    .b(\DFF_800.Q ),
    .y(\DFF_832.D )
  );
  al_and2 _08140_ (
    .a(RESET),
    .b(\DFF_801.Q ),
    .y(\DFF_833.D )
  );
  al_and2 _08141_ (
    .a(RESET),
    .b(\DFF_802.Q ),
    .y(\DFF_834.D )
  );
  al_and2 _08142_ (
    .a(RESET),
    .b(\DFF_803.Q ),
    .y(\DFF_835.D )
  );
  al_and2 _08143_ (
    .a(RESET),
    .b(\DFF_804.Q ),
    .y(\DFF_836.D )
  );
  al_and2 _08144_ (
    .a(RESET),
    .b(\DFF_805.Q ),
    .y(\DFF_837.D )
  );
  al_and2 _08145_ (
    .a(RESET),
    .b(\DFF_806.Q ),
    .y(\DFF_838.D )
  );
  al_and2 _08146_ (
    .a(RESET),
    .b(\DFF_807.Q ),
    .y(\DFF_839.D )
  );
  al_and2 _08147_ (
    .a(RESET),
    .b(\DFF_808.Q ),
    .y(\DFF_840.D )
  );
  al_and2 _08148_ (
    .a(RESET),
    .b(\DFF_809.Q ),
    .y(\DFF_841.D )
  );
  al_and2 _08149_ (
    .a(RESET),
    .b(\DFF_810.Q ),
    .y(\DFF_842.D )
  );
  al_and2 _08150_ (
    .a(RESET),
    .b(\DFF_811.Q ),
    .y(\DFF_843.D )
  );
  al_and2 _08151_ (
    .a(RESET),
    .b(\DFF_812.Q ),
    .y(\DFF_844.D )
  );
  al_and2 _08152_ (
    .a(RESET),
    .b(\DFF_813.Q ),
    .y(\DFF_845.D )
  );
  al_and2 _08153_ (
    .a(RESET),
    .b(\DFF_814.Q ),
    .y(\DFF_846.D )
  );
  al_and2 _08154_ (
    .a(RESET),
    .b(\DFF_815.Q ),
    .y(\DFF_847.D )
  );
  al_and2 _08155_ (
    .a(RESET),
    .b(\DFF_816.Q ),
    .y(\DFF_848.D )
  );
  al_and2 _08156_ (
    .a(RESET),
    .b(\DFF_817.Q ),
    .y(\DFF_849.D )
  );
  al_and2 _08157_ (
    .a(RESET),
    .b(\DFF_818.Q ),
    .y(\DFF_850.D )
  );
  al_and2 _08158_ (
    .a(RESET),
    .b(\DFF_819.Q ),
    .y(\DFF_851.D )
  );
  al_and2 _08159_ (
    .a(RESET),
    .b(\DFF_820.Q ),
    .y(\DFF_852.D )
  );
  al_and2 _08160_ (
    .a(RESET),
    .b(\DFF_821.Q ),
    .y(\DFF_853.D )
  );
  al_and2 _08161_ (
    .a(RESET),
    .b(\DFF_822.Q ),
    .y(\DFF_854.D )
  );
  al_and2 _08162_ (
    .a(RESET),
    .b(\DFF_823.Q ),
    .y(\DFF_855.D )
  );
  al_and2 _08163_ (
    .a(RESET),
    .b(\DFF_824.Q ),
    .y(\DFF_856.D )
  );
  al_and2 _08164_ (
    .a(RESET),
    .b(\DFF_825.Q ),
    .y(\DFF_857.D )
  );
  al_and2 _08165_ (
    .a(RESET),
    .b(\DFF_826.Q ),
    .y(\DFF_858.D )
  );
  al_and2 _08166_ (
    .a(RESET),
    .b(\DFF_827.Q ),
    .y(\DFF_859.D )
  );
  al_and2 _08167_ (
    .a(RESET),
    .b(\DFF_828.Q ),
    .y(\DFF_860.D )
  );
  al_and2 _08168_ (
    .a(RESET),
    .b(\DFF_829.Q ),
    .y(\DFF_861.D )
  );
  al_and2 _08169_ (
    .a(RESET),
    .b(\DFF_830.Q ),
    .y(\DFF_862.D )
  );
  al_and2 _08170_ (
    .a(RESET),
    .b(\DFF_831.Q ),
    .y(\DFF_863.D )
  );
  al_and2 _08171_ (
    .a(RESET),
    .b(\DFF_832.Q ),
    .y(\DFF_864.D )
  );
  al_and2 _08172_ (
    .a(RESET),
    .b(\DFF_833.Q ),
    .y(\DFF_865.D )
  );
  al_and2 _08173_ (
    .a(RESET),
    .b(\DFF_834.Q ),
    .y(\DFF_866.D )
  );
  al_and2 _08174_ (
    .a(RESET),
    .b(\DFF_835.Q ),
    .y(\DFF_867.D )
  );
  al_and2 _08175_ (
    .a(RESET),
    .b(\DFF_836.Q ),
    .y(\DFF_868.D )
  );
  al_and2 _08176_ (
    .a(RESET),
    .b(\DFF_837.Q ),
    .y(\DFF_869.D )
  );
  al_and2 _08177_ (
    .a(RESET),
    .b(\DFF_838.Q ),
    .y(\DFF_870.D )
  );
  al_and2 _08178_ (
    .a(RESET),
    .b(\DFF_839.Q ),
    .y(\DFF_871.D )
  );
  al_and2 _08179_ (
    .a(RESET),
    .b(\DFF_840.Q ),
    .y(\DFF_872.D )
  );
  al_and2 _08180_ (
    .a(RESET),
    .b(\DFF_841.Q ),
    .y(\DFF_873.D )
  );
  al_and2 _08181_ (
    .a(RESET),
    .b(\DFF_842.Q ),
    .y(\DFF_874.D )
  );
  al_and2 _08182_ (
    .a(RESET),
    .b(\DFF_843.Q ),
    .y(\DFF_875.D )
  );
  al_and2 _08183_ (
    .a(RESET),
    .b(\DFF_844.Q ),
    .y(\DFF_876.D )
  );
  al_and2 _08184_ (
    .a(RESET),
    .b(\DFF_845.Q ),
    .y(\DFF_877.D )
  );
  al_and2 _08185_ (
    .a(RESET),
    .b(\DFF_846.Q ),
    .y(\DFF_878.D )
  );
  al_and2 _08186_ (
    .a(RESET),
    .b(\DFF_847.Q ),
    .y(\DFF_879.D )
  );
  al_and2 _08187_ (
    .a(RESET),
    .b(\DFF_848.Q ),
    .y(\DFF_880.D )
  );
  al_and2 _08188_ (
    .a(RESET),
    .b(\DFF_849.Q ),
    .y(\DFF_881.D )
  );
  al_and2 _08189_ (
    .a(RESET),
    .b(\DFF_850.Q ),
    .y(\DFF_882.D )
  );
  al_and2 _08190_ (
    .a(RESET),
    .b(\DFF_851.Q ),
    .y(\DFF_883.D )
  );
  al_and2 _08191_ (
    .a(RESET),
    .b(\DFF_852.Q ),
    .y(\DFF_884.D )
  );
  al_and2 _08192_ (
    .a(RESET),
    .b(\DFF_853.Q ),
    .y(\DFF_885.D )
  );
  al_and2 _08193_ (
    .a(RESET),
    .b(\DFF_854.Q ),
    .y(\DFF_886.D )
  );
  al_and2 _08194_ (
    .a(RESET),
    .b(\DFF_855.Q ),
    .y(\DFF_887.D )
  );
  al_and2 _08195_ (
    .a(RESET),
    .b(\DFF_856.Q ),
    .y(\DFF_888.D )
  );
  al_and2 _08196_ (
    .a(RESET),
    .b(\DFF_857.Q ),
    .y(\DFF_889.D )
  );
  al_and2 _08197_ (
    .a(RESET),
    .b(\DFF_858.Q ),
    .y(\DFF_890.D )
  );
  al_and2 _08198_ (
    .a(RESET),
    .b(\DFF_859.Q ),
    .y(\DFF_891.D )
  );
  al_and2 _08199_ (
    .a(RESET),
    .b(\DFF_860.Q ),
    .y(\DFF_892.D )
  );
  al_and2 _08200_ (
    .a(RESET),
    .b(\DFF_861.Q ),
    .y(\DFF_893.D )
  );
  al_and2 _08201_ (
    .a(RESET),
    .b(\DFF_862.Q ),
    .y(\DFF_894.D )
  );
  al_and2 _08202_ (
    .a(RESET),
    .b(\DFF_863.Q ),
    .y(\DFF_895.D )
  );
  al_and2 _08203_ (
    .a(RESET),
    .b(\DFF_864.Q ),
    .y(\DFF_896.D )
  );
  al_and2 _08204_ (
    .a(RESET),
    .b(\DFF_865.Q ),
    .y(\DFF_897.D )
  );
  al_and2 _08205_ (
    .a(RESET),
    .b(\DFF_866.Q ),
    .y(\DFF_898.D )
  );
  al_and2 _08206_ (
    .a(RESET),
    .b(\DFF_867.Q ),
    .y(\DFF_899.D )
  );
  al_and2 _08207_ (
    .a(RESET),
    .b(\DFF_868.Q ),
    .y(\DFF_900.D )
  );
  al_and2 _08208_ (
    .a(RESET),
    .b(\DFF_869.Q ),
    .y(\DFF_901.D )
  );
  al_and2 _08209_ (
    .a(RESET),
    .b(\DFF_870.Q ),
    .y(\DFF_902.D )
  );
  al_and2 _08210_ (
    .a(RESET),
    .b(\DFF_871.Q ),
    .y(\DFF_903.D )
  );
  al_and2 _08211_ (
    .a(RESET),
    .b(\DFF_872.Q ),
    .y(\DFF_904.D )
  );
  al_and2 _08212_ (
    .a(RESET),
    .b(\DFF_873.Q ),
    .y(\DFF_905.D )
  );
  al_and2 _08213_ (
    .a(RESET),
    .b(\DFF_874.Q ),
    .y(\DFF_906.D )
  );
  al_and2 _08214_ (
    .a(RESET),
    .b(\DFF_875.Q ),
    .y(\DFF_907.D )
  );
  al_and2 _08215_ (
    .a(RESET),
    .b(\DFF_876.Q ),
    .y(\DFF_908.D )
  );
  al_and2 _08216_ (
    .a(RESET),
    .b(\DFF_877.Q ),
    .y(\DFF_909.D )
  );
  al_and2 _08217_ (
    .a(RESET),
    .b(\DFF_878.Q ),
    .y(\DFF_910.D )
  );
  al_and2 _08218_ (
    .a(RESET),
    .b(\DFF_879.Q ),
    .y(\DFF_911.D )
  );
  al_and2 _08219_ (
    .a(RESET),
    .b(\DFF_880.Q ),
    .y(\DFF_912.D )
  );
  al_and2 _08220_ (
    .a(RESET),
    .b(\DFF_881.Q ),
    .y(\DFF_913.D )
  );
  al_and2 _08221_ (
    .a(RESET),
    .b(\DFF_882.Q ),
    .y(\DFF_914.D )
  );
  al_and2 _08222_ (
    .a(RESET),
    .b(\DFF_883.Q ),
    .y(\DFF_915.D )
  );
  al_and2 _08223_ (
    .a(RESET),
    .b(\DFF_884.Q ),
    .y(\DFF_916.D )
  );
  al_and2 _08224_ (
    .a(RESET),
    .b(\DFF_885.Q ),
    .y(\DFF_917.D )
  );
  al_and2 _08225_ (
    .a(RESET),
    .b(\DFF_886.Q ),
    .y(\DFF_918.D )
  );
  al_and2 _08226_ (
    .a(RESET),
    .b(\DFF_887.Q ),
    .y(\DFF_919.D )
  );
  al_and2 _08227_ (
    .a(RESET),
    .b(\DFF_888.Q ),
    .y(\DFF_920.D )
  );
  al_and2 _08228_ (
    .a(RESET),
    .b(\DFF_889.Q ),
    .y(\DFF_921.D )
  );
  al_and2 _08229_ (
    .a(RESET),
    .b(\DFF_890.Q ),
    .y(\DFF_922.D )
  );
  al_and2 _08230_ (
    .a(RESET),
    .b(\DFF_891.Q ),
    .y(\DFF_923.D )
  );
  al_and2 _08231_ (
    .a(RESET),
    .b(\DFF_892.Q ),
    .y(\DFF_924.D )
  );
  al_and2 _08232_ (
    .a(RESET),
    .b(\DFF_893.Q ),
    .y(\DFF_925.D )
  );
  al_and2 _08233_ (
    .a(RESET),
    .b(\DFF_894.Q ),
    .y(\DFF_926.D )
  );
  al_and2 _08234_ (
    .a(RESET),
    .b(\DFF_895.Q ),
    .y(\DFF_927.D )
  );
  al_oa21ftt _08235_ (
    .a(\DFF_927.Q ),
    .b(\DFF_959.Q ),
    .c(RESET),
    .y(_02823_)
  );
  al_aoi21ftf _08236_ (
    .a(\DFF_927.Q ),
    .b(\DFF_959.Q ),
    .c(_02823_),
    .y(\DFF_928.D )
  );
  al_oa21ftt _08237_ (
    .a(\DFF_926.Q ),
    .b(\DFF_928.Q ),
    .c(RESET),
    .y(_02824_)
  );
  al_aoi21ftf _08238_ (
    .a(\DFF_926.Q ),
    .b(\DFF_928.Q ),
    .c(_02824_),
    .y(\DFF_929.D )
  );
  al_oa21ftt _08239_ (
    .a(\DFF_925.Q ),
    .b(\DFF_929.Q ),
    .c(RESET),
    .y(_02825_)
  );
  al_aoi21ftf _08240_ (
    .a(\DFF_925.Q ),
    .b(\DFF_929.Q ),
    .c(_02825_),
    .y(\DFF_930.D )
  );
  al_oa21ftt _08241_ (
    .a(\DFF_924.Q ),
    .b(\DFF_930.Q ),
    .c(RESET),
    .y(_02826_)
  );
  al_aoi21ftf _08242_ (
    .a(\DFF_924.Q ),
    .b(\DFF_930.Q ),
    .c(_02826_),
    .y(\DFF_931.D )
  );
  al_nand2ft _08243_ (
    .a(\DFF_923.Q ),
    .b(\DFF_931.Q ),
    .y(_02827_)
  );
  al_nand2ft _08244_ (
    .a(\DFF_931.Q ),
    .b(\DFF_923.Q ),
    .y(_02828_)
  );
  al_ao21ttf _08245_ (
    .a(_02827_),
    .b(_02828_),
    .c(\DFF_959.Q ),
    .y(_02829_)
  );
  al_nand3ftt _08246_ (
    .a(\DFF_959.Q ),
    .b(_02827_),
    .c(_02828_),
    .y(_02830_)
  );
  al_aoi21 _08247_ (
    .a(_02830_),
    .b(_02829_),
    .c(_00451_),
    .y(\DFF_932.D )
  );
  al_oa21ftt _08248_ (
    .a(\DFF_922.Q ),
    .b(\DFF_932.Q ),
    .c(RESET),
    .y(_02831_)
  );
  al_aoi21ftf _08249_ (
    .a(\DFF_922.Q ),
    .b(\DFF_932.Q ),
    .c(_02831_),
    .y(\DFF_933.D )
  );
  al_oa21ftt _08250_ (
    .a(\DFF_921.Q ),
    .b(\DFF_933.Q ),
    .c(RESET),
    .y(_02832_)
  );
  al_aoi21ftf _08251_ (
    .a(\DFF_921.Q ),
    .b(\DFF_933.Q ),
    .c(_02832_),
    .y(\DFF_934.D )
  );
  al_oa21ftt _08252_ (
    .a(\DFF_920.Q ),
    .b(\DFF_934.Q ),
    .c(RESET),
    .y(_02833_)
  );
  al_aoi21ftf _08253_ (
    .a(\DFF_920.Q ),
    .b(\DFF_934.Q ),
    .c(_02833_),
    .y(\DFF_935.D )
  );
  al_oa21ftt _08254_ (
    .a(\DFF_919.Q ),
    .b(\DFF_935.Q ),
    .c(RESET),
    .y(_02834_)
  );
  al_aoi21ftf _08255_ (
    .a(\DFF_919.Q ),
    .b(\DFF_935.Q ),
    .c(_02834_),
    .y(\DFF_936.D )
  );
  al_oa21ftt _08256_ (
    .a(\DFF_918.Q ),
    .b(\DFF_936.Q ),
    .c(RESET),
    .y(_02835_)
  );
  al_aoi21ftf _08257_ (
    .a(\DFF_918.Q ),
    .b(\DFF_936.Q ),
    .c(_02835_),
    .y(\DFF_937.D )
  );
  al_oa21ftt _08258_ (
    .a(\DFF_917.Q ),
    .b(\DFF_937.Q ),
    .c(RESET),
    .y(_02836_)
  );
  al_aoi21ftf _08259_ (
    .a(\DFF_917.Q ),
    .b(\DFF_937.Q ),
    .c(_02836_),
    .y(\DFF_938.D )
  );
  al_nand2ft _08260_ (
    .a(\DFF_916.Q ),
    .b(\DFF_938.Q ),
    .y(_02837_)
  );
  al_nand2ft _08261_ (
    .a(\DFF_938.Q ),
    .b(\DFF_916.Q ),
    .y(_02838_)
  );
  al_ao21ttf _08262_ (
    .a(_02837_),
    .b(_02838_),
    .c(\DFF_959.Q ),
    .y(_02839_)
  );
  al_nand3ftt _08263_ (
    .a(\DFF_959.Q ),
    .b(_02837_),
    .c(_02838_),
    .y(_02840_)
  );
  al_aoi21 _08264_ (
    .a(_02840_),
    .b(_02839_),
    .c(_00451_),
    .y(\DFF_939.D )
  );
  al_oa21ftt _08265_ (
    .a(\DFF_915.Q ),
    .b(\DFF_939.Q ),
    .c(RESET),
    .y(_02841_)
  );
  al_aoi21ftf _08266_ (
    .a(\DFF_915.Q ),
    .b(\DFF_939.Q ),
    .c(_02841_),
    .y(\DFF_940.D )
  );
  al_oa21ftt _08267_ (
    .a(\DFF_914.Q ),
    .b(\DFF_940.Q ),
    .c(RESET),
    .y(_02842_)
  );
  al_aoi21ftf _08268_ (
    .a(\DFF_914.Q ),
    .b(\DFF_940.Q ),
    .c(_02842_),
    .y(\DFF_941.D )
  );
  al_oa21ftt _08269_ (
    .a(\DFF_913.Q ),
    .b(\DFF_941.Q ),
    .c(RESET),
    .y(_02843_)
  );
  al_aoi21ftf _08270_ (
    .a(\DFF_913.Q ),
    .b(\DFF_941.Q ),
    .c(_02843_),
    .y(\DFF_942.D )
  );
  al_oa21ftt _08271_ (
    .a(\DFF_912.Q ),
    .b(\DFF_942.Q ),
    .c(RESET),
    .y(_02844_)
  );
  al_aoi21ftf _08272_ (
    .a(\DFF_912.Q ),
    .b(\DFF_942.Q ),
    .c(_02844_),
    .y(\DFF_943.D )
  );
  al_nand2ft _08273_ (
    .a(\DFF_911.Q ),
    .b(\DFF_943.Q ),
    .y(_02845_)
  );
  al_nand2ft _08274_ (
    .a(\DFF_943.Q ),
    .b(\DFF_911.Q ),
    .y(_02846_)
  );
  al_ao21ttf _08275_ (
    .a(_02845_),
    .b(_02846_),
    .c(\DFF_959.Q ),
    .y(_02847_)
  );
  al_nand3ftt _08276_ (
    .a(\DFF_959.Q ),
    .b(_02845_),
    .c(_02846_),
    .y(_02848_)
  );
  al_aoi21 _08277_ (
    .a(_02848_),
    .b(_02847_),
    .c(_00451_),
    .y(\DFF_944.D )
  );
  al_oa21ftt _08278_ (
    .a(\DFF_910.Q ),
    .b(\DFF_944.Q ),
    .c(RESET),
    .y(_02849_)
  );
  al_aoi21ftf _08279_ (
    .a(\DFF_910.Q ),
    .b(\DFF_944.Q ),
    .c(_02849_),
    .y(\DFF_945.D )
  );
  al_oa21ftt _08280_ (
    .a(\DFF_909.Q ),
    .b(\DFF_945.Q ),
    .c(RESET),
    .y(_02850_)
  );
  al_aoi21ftf _08281_ (
    .a(\DFF_909.Q ),
    .b(\DFF_945.Q ),
    .c(_02850_),
    .y(\DFF_946.D )
  );
  al_oa21ftt _08282_ (
    .a(\DFF_908.Q ),
    .b(\DFF_946.Q ),
    .c(RESET),
    .y(_02851_)
  );
  al_aoi21ftf _08283_ (
    .a(\DFF_908.Q ),
    .b(\DFF_946.Q ),
    .c(_02851_),
    .y(\DFF_947.D )
  );
  al_oa21ftt _08284_ (
    .a(\DFF_907.Q ),
    .b(\DFF_947.Q ),
    .c(RESET),
    .y(_02852_)
  );
  al_aoi21ftf _08285_ (
    .a(\DFF_907.Q ),
    .b(\DFF_947.Q ),
    .c(_02852_),
    .y(\DFF_948.D )
  );
  al_oa21ftt _08286_ (
    .a(\DFF_906.Q ),
    .b(\DFF_948.Q ),
    .c(RESET),
    .y(_02853_)
  );
  al_aoi21ftf _08287_ (
    .a(\DFF_906.Q ),
    .b(\DFF_948.Q ),
    .c(_02853_),
    .y(\DFF_949.D )
  );
  al_oa21ftt _08288_ (
    .a(\DFF_905.Q ),
    .b(\DFF_949.Q ),
    .c(RESET),
    .y(_02854_)
  );
  al_aoi21ftf _08289_ (
    .a(\DFF_905.Q ),
    .b(\DFF_949.Q ),
    .c(_02854_),
    .y(\DFF_950.D )
  );
  al_oa21ftt _08290_ (
    .a(\DFF_904.Q ),
    .b(\DFF_950.Q ),
    .c(RESET),
    .y(_02855_)
  );
  al_aoi21ftf _08291_ (
    .a(\DFF_904.Q ),
    .b(\DFF_950.Q ),
    .c(_02855_),
    .y(\DFF_951.D )
  );
  al_oa21ftt _08292_ (
    .a(\DFF_903.Q ),
    .b(\DFF_951.Q ),
    .c(RESET),
    .y(_02856_)
  );
  al_aoi21ftf _08293_ (
    .a(\DFF_903.Q ),
    .b(\DFF_951.Q ),
    .c(_02856_),
    .y(\DFF_952.D )
  );
  al_oa21ftt _08294_ (
    .a(\DFF_902.Q ),
    .b(\DFF_952.Q ),
    .c(RESET),
    .y(_02857_)
  );
  al_aoi21ftf _08295_ (
    .a(\DFF_902.Q ),
    .b(\DFF_952.Q ),
    .c(_02857_),
    .y(\DFF_953.D )
  );
  al_oa21ftt _08296_ (
    .a(\DFF_901.Q ),
    .b(\DFF_953.Q ),
    .c(RESET),
    .y(_02858_)
  );
  al_aoi21ftf _08297_ (
    .a(\DFF_901.Q ),
    .b(\DFF_953.Q ),
    .c(_02858_),
    .y(\DFF_954.D )
  );
  al_oa21ftt _08298_ (
    .a(\DFF_900.Q ),
    .b(\DFF_954.Q ),
    .c(RESET),
    .y(_02859_)
  );
  al_aoi21ftf _08299_ (
    .a(\DFF_900.Q ),
    .b(\DFF_954.Q ),
    .c(_02859_),
    .y(\DFF_955.D )
  );
  al_oa21ftt _08300_ (
    .a(\DFF_899.Q ),
    .b(\DFF_955.Q ),
    .c(RESET),
    .y(_02860_)
  );
  al_aoi21ftf _08301_ (
    .a(\DFF_899.Q ),
    .b(\DFF_955.Q ),
    .c(_02860_),
    .y(\DFF_956.D )
  );
  al_oa21ftt _08302_ (
    .a(\DFF_898.Q ),
    .b(\DFF_956.Q ),
    .c(RESET),
    .y(_02861_)
  );
  al_aoi21ftf _08303_ (
    .a(\DFF_898.Q ),
    .b(\DFF_956.Q ),
    .c(_02861_),
    .y(\DFF_957.D )
  );
  al_oa21ftt _08304_ (
    .a(\DFF_897.Q ),
    .b(\DFF_957.Q ),
    .c(RESET),
    .y(_02862_)
  );
  al_aoi21ftf _08305_ (
    .a(\DFF_897.Q ),
    .b(\DFF_957.Q ),
    .c(_02862_),
    .y(\DFF_958.D )
  );
  al_oa21ftt _08306_ (
    .a(\DFF_896.Q ),
    .b(\DFF_958.Q ),
    .c(RESET),
    .y(_02863_)
  );
  al_aoi21ftf _08307_ (
    .a(\DFF_896.Q ),
    .b(\DFF_958.Q ),
    .c(_02863_),
    .y(\DFF_959.D )
  );
  al_and2 _08308_ (
    .a(RESET),
    .b(\DFF_961.Q ),
    .y(\DFF_960.D )
  );
  al_and2 _08309_ (
    .a(RESET),
    .b(\DFF_962.Q ),
    .y(\DFF_961.D )
  );
  al_and2 _08310_ (
    .a(RESET),
    .b(\DFF_963.Q ),
    .y(\DFF_962.D )
  );
  al_and2 _08311_ (
    .a(RESET),
    .b(\DFF_964.Q ),
    .y(\DFF_963.D )
  );
  al_and2 _08312_ (
    .a(RESET),
    .b(\DFF_965.Q ),
    .y(\DFF_964.D )
  );
  al_and2 _08313_ (
    .a(RESET),
    .b(\DFF_966.Q ),
    .y(\DFF_965.D )
  );
  al_and2 _08314_ (
    .a(RESET),
    .b(\DFF_967.Q ),
    .y(\DFF_966.D )
  );
  al_and2 _08315_ (
    .a(RESET),
    .b(\DFF_968.Q ),
    .y(\DFF_967.D )
  );
  al_and2 _08316_ (
    .a(RESET),
    .b(\DFF_969.Q ),
    .y(\DFF_968.D )
  );
  al_and2 _08317_ (
    .a(RESET),
    .b(\DFF_970.Q ),
    .y(\DFF_969.D )
  );
  al_and2 _08318_ (
    .a(RESET),
    .b(\DFF_971.Q ),
    .y(\DFF_970.D )
  );
  al_and2 _08319_ (
    .a(RESET),
    .b(\DFF_972.Q ),
    .y(\DFF_971.D )
  );
  al_and2 _08320_ (
    .a(RESET),
    .b(\DFF_973.Q ),
    .y(\DFF_972.D )
  );
  al_and2 _08321_ (
    .a(RESET),
    .b(\DFF_974.Q ),
    .y(\DFF_973.D )
  );
  al_and2 _08322_ (
    .a(RESET),
    .b(\DFF_975.Q ),
    .y(\DFF_974.D )
  );
  al_and2 _08323_ (
    .a(RESET),
    .b(\DFF_976.Q ),
    .y(\DFF_975.D )
  );
  al_and2 _08324_ (
    .a(RESET),
    .b(\DFF_977.Q ),
    .y(\DFF_976.D )
  );
  al_and2 _08325_ (
    .a(RESET),
    .b(\DFF_978.Q ),
    .y(\DFF_977.D )
  );
  al_and2 _08326_ (
    .a(RESET),
    .b(\DFF_979.Q ),
    .y(\DFF_978.D )
  );
  al_and2 _08327_ (
    .a(RESET),
    .b(\DFF_980.Q ),
    .y(\DFF_979.D )
  );
  al_and2 _08328_ (
    .a(RESET),
    .b(\DFF_981.Q ),
    .y(\DFF_980.D )
  );
  al_and2 _08329_ (
    .a(RESET),
    .b(\DFF_982.Q ),
    .y(\DFF_981.D )
  );
  al_and2 _08330_ (
    .a(RESET),
    .b(\DFF_983.Q ),
    .y(\DFF_982.D )
  );
  al_and2 _08331_ (
    .a(RESET),
    .b(\DFF_984.Q ),
    .y(\DFF_983.D )
  );
  al_and2 _08332_ (
    .a(RESET),
    .b(\DFF_985.Q ),
    .y(\DFF_984.D )
  );
  al_and2 _08333_ (
    .a(RESET),
    .b(\DFF_986.Q ),
    .y(\DFF_985.D )
  );
  al_and2 _08334_ (
    .a(RESET),
    .b(\DFF_987.Q ),
    .y(\DFF_986.D )
  );
  al_and2 _08335_ (
    .a(RESET),
    .b(\DFF_988.Q ),
    .y(\DFF_987.D )
  );
  al_and2 _08336_ (
    .a(RESET),
    .b(\DFF_989.Q ),
    .y(\DFF_988.D )
  );
  al_and2 _08337_ (
    .a(RESET),
    .b(\DFF_990.Q ),
    .y(\DFF_989.D )
  );
  al_and2 _08338_ (
    .a(RESET),
    .b(\DFF_991.Q ),
    .y(\DFF_990.D )
  );
  al_and2ft _08339_ (
    .a(\DFF_960.Q ),
    .b(RESET),
    .y(\DFF_991.D )
  );
  al_or2 _08340_ (
    .a(TM1),
    .b(\DFF_1248.Q ),
    .y(_02864_)
  );
  al_nand2 _08341_ (
    .a(TM1),
    .b(\DFF_1248.Q ),
    .y(_02865_)
  );
  al_nand3 _08342_ (
    .a(\DFF_1280.Q ),
    .b(_02864_),
    .c(_02865_),
    .y(_02866_)
  );
  al_nand2ft _08343_ (
    .a(TM1),
    .b(\DFF_1248.Q ),
    .y(_02867_)
  );
  al_and2ft _08344_ (
    .a(\DFF_1248.Q ),
    .b(TM1),
    .y(_02868_)
  );
  al_and3fft _08345_ (
    .a(\DFF_1280.Q ),
    .b(_02868_),
    .c(_02867_),
    .y(_02869_)
  );
  al_and2ft _08346_ (
    .a(\DFF_1216.Q ),
    .b(\DFF_1184.Q ),
    .y(_02870_)
  );
  al_nand2ft _08347_ (
    .a(\DFF_1184.Q ),
    .b(\DFF_1216.Q ),
    .y(_02871_)
  );
  al_nand2ft _08348_ (
    .a(_02870_),
    .b(_02871_),
    .y(_02872_)
  );
  al_oai21ftf _08349_ (
    .a(_02866_),
    .b(_02869_),
    .c(_02872_),
    .y(_02873_)
  );
  al_nand3ftt _08350_ (
    .a(_02869_),
    .b(_02866_),
    .c(_02872_),
    .y(_02874_)
  );
  al_nand3 _08351_ (
    .a(_00448_),
    .b(_02873_),
    .c(_02874_),
    .y(_02875_)
  );
  al_aoi21 _08352_ (
    .a(TM0),
    .b(\DFF_1151.Q ),
    .c(TM1),
    .y(_02876_)
  );
  al_nand2 _08353_ (
    .a(_02876_),
    .b(_02875_),
    .y(_02877_)
  );
  al_aoi21ttf _08354_ (
    .a(\DFF_960.Q ),
    .b(TM0),
    .c(TM1),
    .y(_02878_)
  );
  al_and2 _08355_ (
    .a(_02878_),
    .b(_02386_),
    .y(_02879_)
  );
  al_nor3fft _08356_ (
    .a(RESET),
    .b(_02877_),
    .c(_02879_),
    .y(\DFF_992.D )
  );
  al_or2 _08357_ (
    .a(TM1),
    .b(\DFF_1249.Q ),
    .y(_02880_)
  );
  al_nand2 _08358_ (
    .a(TM1),
    .b(\DFF_1249.Q ),
    .y(_02881_)
  );
  al_nand3 _08359_ (
    .a(\DFF_1281.Q ),
    .b(_02880_),
    .c(_02881_),
    .y(_02882_)
  );
  al_nand2ft _08360_ (
    .a(TM1),
    .b(\DFF_1249.Q ),
    .y(_02883_)
  );
  al_and2ft _08361_ (
    .a(\DFF_1249.Q ),
    .b(TM1),
    .y(_02884_)
  );
  al_and3fft _08362_ (
    .a(\DFF_1281.Q ),
    .b(_02884_),
    .c(_02883_),
    .y(_02885_)
  );
  al_and2ft _08363_ (
    .a(\DFF_1217.Q ),
    .b(\DFF_1185.Q ),
    .y(_02886_)
  );
  al_nand2ft _08364_ (
    .a(\DFF_1185.Q ),
    .b(\DFF_1217.Q ),
    .y(_02887_)
  );
  al_nand2ft _08365_ (
    .a(_02886_),
    .b(_02887_),
    .y(_02888_)
  );
  al_oai21ftf _08366_ (
    .a(_02882_),
    .b(_02885_),
    .c(_02888_),
    .y(_02889_)
  );
  al_nand3ftt _08367_ (
    .a(_02885_),
    .b(_02882_),
    .c(_02888_),
    .y(_02890_)
  );
  al_nand3 _08368_ (
    .a(_00448_),
    .b(_02889_),
    .c(_02890_),
    .y(_02891_)
  );
  al_aoi21 _08369_ (
    .a(TM0),
    .b(\DFF_1150.Q ),
    .c(TM1),
    .y(_02892_)
  );
  al_nand2 _08370_ (
    .a(_02892_),
    .b(_02891_),
    .y(_02893_)
  );
  al_aoi21ttf _08371_ (
    .a(TM0),
    .b(\DFF_961.Q ),
    .c(TM1),
    .y(_02894_)
  );
  al_and2 _08372_ (
    .a(_02894_),
    .b(_02402_),
    .y(_02895_)
  );
  al_nor3fft _08373_ (
    .a(RESET),
    .b(_02893_),
    .c(_02895_),
    .y(\DFF_993.D )
  );
  al_or2 _08374_ (
    .a(TM1),
    .b(\DFF_1250.Q ),
    .y(_02896_)
  );
  al_nand2 _08375_ (
    .a(TM1),
    .b(\DFF_1250.Q ),
    .y(_02897_)
  );
  al_nand3 _08376_ (
    .a(\DFF_1282.Q ),
    .b(_02896_),
    .c(_02897_),
    .y(_02898_)
  );
  al_nand2ft _08377_ (
    .a(TM1),
    .b(\DFF_1250.Q ),
    .y(_02899_)
  );
  al_and2ft _08378_ (
    .a(\DFF_1250.Q ),
    .b(TM1),
    .y(_02900_)
  );
  al_and3fft _08379_ (
    .a(\DFF_1282.Q ),
    .b(_02900_),
    .c(_02899_),
    .y(_02901_)
  );
  al_and2ft _08380_ (
    .a(\DFF_1218.Q ),
    .b(\DFF_1186.Q ),
    .y(_02902_)
  );
  al_nand2ft _08381_ (
    .a(\DFF_1186.Q ),
    .b(\DFF_1218.Q ),
    .y(_02903_)
  );
  al_nand2ft _08382_ (
    .a(_02902_),
    .b(_02903_),
    .y(_02904_)
  );
  al_oai21ftf _08383_ (
    .a(_02898_),
    .b(_02901_),
    .c(_02904_),
    .y(_02905_)
  );
  al_nand3ftt _08384_ (
    .a(_02901_),
    .b(_02898_),
    .c(_02904_),
    .y(_02906_)
  );
  al_nand3 _08385_ (
    .a(_00448_),
    .b(_02905_),
    .c(_02906_),
    .y(_02907_)
  );
  al_aoi21 _08386_ (
    .a(TM0),
    .b(\DFF_1149.Q ),
    .c(TM1),
    .y(_02908_)
  );
  al_nand2 _08387_ (
    .a(_02908_),
    .b(_02907_),
    .y(_02909_)
  );
  al_aoi21ttf _08388_ (
    .a(TM0),
    .b(\DFF_962.Q ),
    .c(TM1),
    .y(_02910_)
  );
  al_and2 _08389_ (
    .a(_02910_),
    .b(_02418_),
    .y(_02911_)
  );
  al_nor3fft _08390_ (
    .a(RESET),
    .b(_02909_),
    .c(_02911_),
    .y(\DFF_994.D )
  );
  al_or2 _08391_ (
    .a(TM1),
    .b(\DFF_1251.Q ),
    .y(_02912_)
  );
  al_nand2 _08392_ (
    .a(TM1),
    .b(\DFF_1251.Q ),
    .y(_02913_)
  );
  al_nand3 _08393_ (
    .a(\DFF_1283.Q ),
    .b(_02912_),
    .c(_02913_),
    .y(_02914_)
  );
  al_nand2ft _08394_ (
    .a(TM1),
    .b(\DFF_1251.Q ),
    .y(_02915_)
  );
  al_and2ft _08395_ (
    .a(\DFF_1251.Q ),
    .b(TM1),
    .y(_02916_)
  );
  al_and3fft _08396_ (
    .a(\DFF_1283.Q ),
    .b(_02916_),
    .c(_02915_),
    .y(_02917_)
  );
  al_and2ft _08397_ (
    .a(\DFF_1219.Q ),
    .b(\DFF_1187.Q ),
    .y(_02918_)
  );
  al_nand2ft _08398_ (
    .a(\DFF_1187.Q ),
    .b(\DFF_1219.Q ),
    .y(_02919_)
  );
  al_nand2ft _08399_ (
    .a(_02918_),
    .b(_02919_),
    .y(_02920_)
  );
  al_oai21ftf _08400_ (
    .a(_02914_),
    .b(_02917_),
    .c(_02920_),
    .y(_02921_)
  );
  al_nand3ftt _08401_ (
    .a(_02917_),
    .b(_02914_),
    .c(_02920_),
    .y(_02922_)
  );
  al_nand3 _08402_ (
    .a(_00448_),
    .b(_02921_),
    .c(_02922_),
    .y(_02923_)
  );
  al_aoi21 _08403_ (
    .a(TM0),
    .b(\DFF_1148.Q ),
    .c(TM1),
    .y(_02924_)
  );
  al_nand2 _08404_ (
    .a(_02924_),
    .b(_02923_),
    .y(_02925_)
  );
  al_aoi21ttf _08405_ (
    .a(TM0),
    .b(\DFF_963.Q ),
    .c(TM1),
    .y(_02926_)
  );
  al_and2 _08406_ (
    .a(_02926_),
    .b(_02434_),
    .y(_02927_)
  );
  al_nor3fft _08407_ (
    .a(RESET),
    .b(_02925_),
    .c(_02927_),
    .y(\DFF_995.D )
  );
  al_or2 _08408_ (
    .a(TM1),
    .b(\DFF_1252.Q ),
    .y(_02928_)
  );
  al_nand2 _08409_ (
    .a(TM1),
    .b(\DFF_1252.Q ),
    .y(_02929_)
  );
  al_nand3 _08410_ (
    .a(\DFF_1284.Q ),
    .b(_02928_),
    .c(_02929_),
    .y(_02930_)
  );
  al_nand2ft _08411_ (
    .a(TM1),
    .b(\DFF_1252.Q ),
    .y(_02931_)
  );
  al_and2ft _08412_ (
    .a(\DFF_1252.Q ),
    .b(TM1),
    .y(_02932_)
  );
  al_and3fft _08413_ (
    .a(\DFF_1284.Q ),
    .b(_02932_),
    .c(_02931_),
    .y(_02933_)
  );
  al_and2ft _08414_ (
    .a(\DFF_1220.Q ),
    .b(\DFF_1188.Q ),
    .y(_02934_)
  );
  al_nand2ft _08415_ (
    .a(\DFF_1188.Q ),
    .b(\DFF_1220.Q ),
    .y(_02935_)
  );
  al_nand2ft _08416_ (
    .a(_02934_),
    .b(_02935_),
    .y(_02936_)
  );
  al_oai21ftf _08417_ (
    .a(_02930_),
    .b(_02933_),
    .c(_02936_),
    .y(_02937_)
  );
  al_nand3ftt _08418_ (
    .a(_02933_),
    .b(_02930_),
    .c(_02936_),
    .y(_02938_)
  );
  al_nand3 _08419_ (
    .a(_00448_),
    .b(_02937_),
    .c(_02938_),
    .y(_02939_)
  );
  al_aoi21 _08420_ (
    .a(TM0),
    .b(\DFF_1147.Q ),
    .c(TM1),
    .y(_02940_)
  );
  al_nand2 _08421_ (
    .a(_02940_),
    .b(_02939_),
    .y(_02941_)
  );
  al_aoi21ttf _08422_ (
    .a(TM0),
    .b(\DFF_964.Q ),
    .c(TM1),
    .y(_02942_)
  );
  al_and2 _08423_ (
    .a(_02942_),
    .b(_02450_),
    .y(_02943_)
  );
  al_nor3fft _08424_ (
    .a(RESET),
    .b(_02941_),
    .c(_02943_),
    .y(\DFF_996.D )
  );
  al_or2 _08425_ (
    .a(TM1),
    .b(\DFF_1253.Q ),
    .y(_02944_)
  );
  al_nand2 _08426_ (
    .a(TM1),
    .b(\DFF_1253.Q ),
    .y(_02945_)
  );
  al_nand3 _08427_ (
    .a(\DFF_1285.Q ),
    .b(_02944_),
    .c(_02945_),
    .y(_02946_)
  );
  al_nand2ft _08428_ (
    .a(TM1),
    .b(\DFF_1253.Q ),
    .y(_02947_)
  );
  al_and2ft _08429_ (
    .a(\DFF_1253.Q ),
    .b(TM1),
    .y(_02948_)
  );
  al_and3fft _08430_ (
    .a(\DFF_1285.Q ),
    .b(_02948_),
    .c(_02947_),
    .y(_02949_)
  );
  al_and2ft _08431_ (
    .a(\DFF_1221.Q ),
    .b(\DFF_1189.Q ),
    .y(_02950_)
  );
  al_nand2ft _08432_ (
    .a(\DFF_1189.Q ),
    .b(\DFF_1221.Q ),
    .y(_02951_)
  );
  al_nand2ft _08433_ (
    .a(_02950_),
    .b(_02951_),
    .y(_02952_)
  );
  al_oai21ftf _08434_ (
    .a(_02946_),
    .b(_02949_),
    .c(_02952_),
    .y(_02953_)
  );
  al_nand3ftt _08435_ (
    .a(_02949_),
    .b(_02946_),
    .c(_02952_),
    .y(_02954_)
  );
  al_nand3 _08436_ (
    .a(_00448_),
    .b(_02953_),
    .c(_02954_),
    .y(_02955_)
  );
  al_aoi21 _08437_ (
    .a(TM0),
    .b(\DFF_1146.Q ),
    .c(TM1),
    .y(_02956_)
  );
  al_nand2 _08438_ (
    .a(_02956_),
    .b(_02955_),
    .y(_02957_)
  );
  al_aoi21ttf _08439_ (
    .a(TM0),
    .b(\DFF_965.Q ),
    .c(TM1),
    .y(_02958_)
  );
  al_and2 _08440_ (
    .a(_02958_),
    .b(_02466_),
    .y(_02959_)
  );
  al_nor3fft _08441_ (
    .a(RESET),
    .b(_02957_),
    .c(_02959_),
    .y(\DFF_997.D )
  );
  al_or2 _08442_ (
    .a(TM1),
    .b(\DFF_1254.Q ),
    .y(_02960_)
  );
  al_nand2 _08443_ (
    .a(TM1),
    .b(\DFF_1254.Q ),
    .y(_02961_)
  );
  al_nand3 _08444_ (
    .a(\DFF_1286.Q ),
    .b(_02960_),
    .c(_02961_),
    .y(_02962_)
  );
  al_nand2ft _08445_ (
    .a(TM1),
    .b(\DFF_1254.Q ),
    .y(_02963_)
  );
  al_and2ft _08446_ (
    .a(\DFF_1254.Q ),
    .b(TM1),
    .y(_02964_)
  );
  al_and3fft _08447_ (
    .a(\DFF_1286.Q ),
    .b(_02964_),
    .c(_02963_),
    .y(_02965_)
  );
  al_and2ft _08448_ (
    .a(\DFF_1222.Q ),
    .b(\DFF_1190.Q ),
    .y(_02966_)
  );
  al_nand2ft _08449_ (
    .a(\DFF_1190.Q ),
    .b(\DFF_1222.Q ),
    .y(_02967_)
  );
  al_nand2ft _08450_ (
    .a(_02966_),
    .b(_02967_),
    .y(_02968_)
  );
  al_oai21ftf _08451_ (
    .a(_02962_),
    .b(_02965_),
    .c(_02968_),
    .y(_02969_)
  );
  al_nand3ftt _08452_ (
    .a(_02965_),
    .b(_02962_),
    .c(_02968_),
    .y(_02970_)
  );
  al_nand3 _08453_ (
    .a(_00448_),
    .b(_02969_),
    .c(_02970_),
    .y(_02971_)
  );
  al_aoi21 _08454_ (
    .a(TM0),
    .b(\DFF_1145.Q ),
    .c(TM1),
    .y(_02972_)
  );
  al_nand2 _08455_ (
    .a(_02972_),
    .b(_02971_),
    .y(_02973_)
  );
  al_aoi21ttf _08456_ (
    .a(TM0),
    .b(\DFF_966.Q ),
    .c(TM1),
    .y(_02974_)
  );
  al_and2 _08457_ (
    .a(_02974_),
    .b(_02482_),
    .y(_02975_)
  );
  al_nor3fft _08458_ (
    .a(RESET),
    .b(_02973_),
    .c(_02975_),
    .y(\DFF_998.D )
  );
  al_or2 _08459_ (
    .a(TM1),
    .b(\DFF_1255.Q ),
    .y(_02976_)
  );
  al_nand2 _08460_ (
    .a(TM1),
    .b(\DFF_1255.Q ),
    .y(_02977_)
  );
  al_nand3 _08461_ (
    .a(\DFF_1287.Q ),
    .b(_02976_),
    .c(_02977_),
    .y(_02978_)
  );
  al_nand2ft _08462_ (
    .a(TM1),
    .b(\DFF_1255.Q ),
    .y(_02979_)
  );
  al_and2ft _08463_ (
    .a(\DFF_1255.Q ),
    .b(TM1),
    .y(_02980_)
  );
  al_and3fft _08464_ (
    .a(\DFF_1287.Q ),
    .b(_02980_),
    .c(_02979_),
    .y(_02981_)
  );
  al_and2ft _08465_ (
    .a(\DFF_1223.Q ),
    .b(\DFF_1191.Q ),
    .y(_02982_)
  );
  al_nand2ft _08466_ (
    .a(\DFF_1191.Q ),
    .b(\DFF_1223.Q ),
    .y(_02983_)
  );
  al_nand2ft _08467_ (
    .a(_02982_),
    .b(_02983_),
    .y(_02984_)
  );
  al_oai21ftf _08468_ (
    .a(_02978_),
    .b(_02981_),
    .c(_02984_),
    .y(_02985_)
  );
  al_nand3ftt _08469_ (
    .a(_02981_),
    .b(_02978_),
    .c(_02984_),
    .y(_02986_)
  );
  al_nand3 _08470_ (
    .a(_00448_),
    .b(_02985_),
    .c(_02986_),
    .y(_02987_)
  );
  al_aoi21 _08471_ (
    .a(TM0),
    .b(\DFF_1144.Q ),
    .c(TM1),
    .y(_02988_)
  );
  al_nand2 _08472_ (
    .a(_02988_),
    .b(_02987_),
    .y(_02989_)
  );
  al_aoi21ttf _08473_ (
    .a(TM0),
    .b(\DFF_967.Q ),
    .c(TM1),
    .y(_02990_)
  );
  al_and2 _08474_ (
    .a(_02990_),
    .b(_02498_),
    .y(_02991_)
  );
  al_nor3fft _08475_ (
    .a(RESET),
    .b(_02989_),
    .c(_02991_),
    .y(\DFF_999.D )
  );
  al_or2 _08476_ (
    .a(TM1),
    .b(\DFF_1256.Q ),
    .y(_02992_)
  );
  al_nand2 _08477_ (
    .a(TM1),
    .b(\DFF_1256.Q ),
    .y(_02993_)
  );
  al_nand3 _08478_ (
    .a(\DFF_1288.Q ),
    .b(_02992_),
    .c(_02993_),
    .y(_02994_)
  );
  al_nand2ft _08479_ (
    .a(TM1),
    .b(\DFF_1256.Q ),
    .y(_02995_)
  );
  al_and2ft _08480_ (
    .a(\DFF_1256.Q ),
    .b(TM1),
    .y(_02996_)
  );
  al_and3fft _08481_ (
    .a(\DFF_1288.Q ),
    .b(_02996_),
    .c(_02995_),
    .y(_02997_)
  );
  al_and2ft _08482_ (
    .a(\DFF_1224.Q ),
    .b(\DFF_1192.Q ),
    .y(_02998_)
  );
  al_nand2ft _08483_ (
    .a(\DFF_1192.Q ),
    .b(\DFF_1224.Q ),
    .y(_02999_)
  );
  al_nand2ft _08484_ (
    .a(_02998_),
    .b(_02999_),
    .y(_03000_)
  );
  al_oai21ftf _08485_ (
    .a(_02994_),
    .b(_02997_),
    .c(_03000_),
    .y(_03001_)
  );
  al_nand3ftt _08486_ (
    .a(_02997_),
    .b(_02994_),
    .c(_03000_),
    .y(_03002_)
  );
  al_nand3 _08487_ (
    .a(_00448_),
    .b(_03001_),
    .c(_03002_),
    .y(_03003_)
  );
  al_aoi21 _08488_ (
    .a(TM0),
    .b(\DFF_1143.Q ),
    .c(TM1),
    .y(_03004_)
  );
  al_nand2 _08489_ (
    .a(_03004_),
    .b(_03003_),
    .y(_03005_)
  );
  al_aoi21ttf _08490_ (
    .a(TM0),
    .b(\DFF_968.Q ),
    .c(TM1),
    .y(_03006_)
  );
  al_and2 _08491_ (
    .a(_03006_),
    .b(_02514_),
    .y(_03007_)
  );
  al_nor3fft _08492_ (
    .a(RESET),
    .b(_03005_),
    .c(_03007_),
    .y(\DFF_1000.D )
  );
  al_or2 _08493_ (
    .a(TM1),
    .b(\DFF_1257.Q ),
    .y(_03008_)
  );
  al_nand2 _08494_ (
    .a(TM1),
    .b(\DFF_1257.Q ),
    .y(_03009_)
  );
  al_nand3 _08495_ (
    .a(\DFF_1289.Q ),
    .b(_03008_),
    .c(_03009_),
    .y(_03010_)
  );
  al_nand2ft _08496_ (
    .a(TM1),
    .b(\DFF_1257.Q ),
    .y(_03011_)
  );
  al_and2ft _08497_ (
    .a(\DFF_1257.Q ),
    .b(TM1),
    .y(_03012_)
  );
  al_and3fft _08498_ (
    .a(\DFF_1289.Q ),
    .b(_03012_),
    .c(_03011_),
    .y(_03013_)
  );
  al_and2ft _08499_ (
    .a(\DFF_1225.Q ),
    .b(\DFF_1193.Q ),
    .y(_03014_)
  );
  al_nand2ft _08500_ (
    .a(\DFF_1193.Q ),
    .b(\DFF_1225.Q ),
    .y(_03015_)
  );
  al_nand2ft _08501_ (
    .a(_03014_),
    .b(_03015_),
    .y(_03016_)
  );
  al_oai21ftf _08502_ (
    .a(_03010_),
    .b(_03013_),
    .c(_03016_),
    .y(_03017_)
  );
  al_nand3ftt _08503_ (
    .a(_03013_),
    .b(_03010_),
    .c(_03016_),
    .y(_03018_)
  );
  al_nand3 _08504_ (
    .a(_00448_),
    .b(_03017_),
    .c(_03018_),
    .y(_03019_)
  );
  al_aoi21 _08505_ (
    .a(TM0),
    .b(\DFF_1142.Q ),
    .c(TM1),
    .y(_03020_)
  );
  al_nand2 _08506_ (
    .a(_03020_),
    .b(_03019_),
    .y(_03021_)
  );
  al_aoi21ttf _08507_ (
    .a(TM0),
    .b(\DFF_969.Q ),
    .c(TM1),
    .y(_03022_)
  );
  al_and2 _08508_ (
    .a(_03022_),
    .b(_02530_),
    .y(_03023_)
  );
  al_nor3fft _08509_ (
    .a(RESET),
    .b(_03021_),
    .c(_03023_),
    .y(\DFF_1001.D )
  );
  al_or2 _08510_ (
    .a(TM1),
    .b(\DFF_1258.Q ),
    .y(_03024_)
  );
  al_nand2 _08511_ (
    .a(TM1),
    .b(\DFF_1258.Q ),
    .y(_03025_)
  );
  al_nand3 _08512_ (
    .a(\DFF_1290.Q ),
    .b(_03024_),
    .c(_03025_),
    .y(_03026_)
  );
  al_nand2ft _08513_ (
    .a(TM1),
    .b(\DFF_1258.Q ),
    .y(_03027_)
  );
  al_and2ft _08514_ (
    .a(\DFF_1258.Q ),
    .b(TM1),
    .y(_03028_)
  );
  al_and3fft _08515_ (
    .a(\DFF_1290.Q ),
    .b(_03028_),
    .c(_03027_),
    .y(_03029_)
  );
  al_and2ft _08516_ (
    .a(\DFF_1226.Q ),
    .b(\DFF_1194.Q ),
    .y(_03030_)
  );
  al_nand2ft _08517_ (
    .a(\DFF_1194.Q ),
    .b(\DFF_1226.Q ),
    .y(_03031_)
  );
  al_nand2ft _08518_ (
    .a(_03030_),
    .b(_03031_),
    .y(_03032_)
  );
  al_oai21ftf _08519_ (
    .a(_03026_),
    .b(_03029_),
    .c(_03032_),
    .y(_03033_)
  );
  al_nand3ftt _08520_ (
    .a(_03029_),
    .b(_03026_),
    .c(_03032_),
    .y(_03034_)
  );
  al_nand3 _08521_ (
    .a(_00448_),
    .b(_03033_),
    .c(_03034_),
    .y(_03035_)
  );
  al_aoi21 _08522_ (
    .a(TM0),
    .b(\DFF_1141.Q ),
    .c(TM1),
    .y(_03036_)
  );
  al_nand2 _08523_ (
    .a(_03036_),
    .b(_03035_),
    .y(_03037_)
  );
  al_aoi21ttf _08524_ (
    .a(TM0),
    .b(\DFF_970.Q ),
    .c(TM1),
    .y(_03038_)
  );
  al_and2 _08525_ (
    .a(_03038_),
    .b(_02546_),
    .y(_03039_)
  );
  al_nor3fft _08526_ (
    .a(RESET),
    .b(_03037_),
    .c(_03039_),
    .y(\DFF_1002.D )
  );
  al_or2 _08527_ (
    .a(TM1),
    .b(\DFF_1259.Q ),
    .y(_03040_)
  );
  al_nand2 _08528_ (
    .a(TM1),
    .b(\DFF_1259.Q ),
    .y(_03041_)
  );
  al_nand3 _08529_ (
    .a(\DFF_1291.Q ),
    .b(_03040_),
    .c(_03041_),
    .y(_03042_)
  );
  al_nand2ft _08530_ (
    .a(TM1),
    .b(\DFF_1259.Q ),
    .y(_03043_)
  );
  al_and2ft _08531_ (
    .a(\DFF_1259.Q ),
    .b(TM1),
    .y(_03044_)
  );
  al_and3fft _08532_ (
    .a(\DFF_1291.Q ),
    .b(_03044_),
    .c(_03043_),
    .y(_03045_)
  );
  al_and2ft _08533_ (
    .a(\DFF_1227.Q ),
    .b(\DFF_1195.Q ),
    .y(_03046_)
  );
  al_nand2ft _08534_ (
    .a(\DFF_1195.Q ),
    .b(\DFF_1227.Q ),
    .y(_03047_)
  );
  al_nand2ft _08535_ (
    .a(_03046_),
    .b(_03047_),
    .y(_03048_)
  );
  al_oai21ftf _08536_ (
    .a(_03042_),
    .b(_03045_),
    .c(_03048_),
    .y(_03049_)
  );
  al_nand3ftt _08537_ (
    .a(_03045_),
    .b(_03042_),
    .c(_03048_),
    .y(_03050_)
  );
  al_nand3 _08538_ (
    .a(_00448_),
    .b(_03049_),
    .c(_03050_),
    .y(_03051_)
  );
  al_aoi21 _08539_ (
    .a(TM0),
    .b(\DFF_1140.Q ),
    .c(TM1),
    .y(_03052_)
  );
  al_nand2 _08540_ (
    .a(_03052_),
    .b(_03051_),
    .y(_03053_)
  );
  al_aoi21ttf _08541_ (
    .a(TM0),
    .b(\DFF_971.Q ),
    .c(TM1),
    .y(_03054_)
  );
  al_and2 _08542_ (
    .a(_03054_),
    .b(_02562_),
    .y(_03055_)
  );
  al_nor3fft _08543_ (
    .a(RESET),
    .b(_03053_),
    .c(_03055_),
    .y(\DFF_1003.D )
  );
  al_or2 _08544_ (
    .a(TM1),
    .b(\DFF_1260.Q ),
    .y(_03056_)
  );
  al_nand2 _08545_ (
    .a(TM1),
    .b(\DFF_1260.Q ),
    .y(_03057_)
  );
  al_nand3 _08546_ (
    .a(\DFF_1292.Q ),
    .b(_03056_),
    .c(_03057_),
    .y(_03058_)
  );
  al_nand2ft _08547_ (
    .a(TM1),
    .b(\DFF_1260.Q ),
    .y(_03059_)
  );
  al_and2ft _08548_ (
    .a(\DFF_1260.Q ),
    .b(TM1),
    .y(_03060_)
  );
  al_and3fft _08549_ (
    .a(\DFF_1292.Q ),
    .b(_03060_),
    .c(_03059_),
    .y(_03061_)
  );
  al_and2ft _08550_ (
    .a(\DFF_1228.Q ),
    .b(\DFF_1196.Q ),
    .y(_03062_)
  );
  al_nand2ft _08551_ (
    .a(\DFF_1196.Q ),
    .b(\DFF_1228.Q ),
    .y(_03063_)
  );
  al_nand2ft _08552_ (
    .a(_03062_),
    .b(_03063_),
    .y(_03064_)
  );
  al_oai21ftf _08553_ (
    .a(_03058_),
    .b(_03061_),
    .c(_03064_),
    .y(_03065_)
  );
  al_nand3ftt _08554_ (
    .a(_03061_),
    .b(_03058_),
    .c(_03064_),
    .y(_03066_)
  );
  al_nand3 _08555_ (
    .a(_00448_),
    .b(_03065_),
    .c(_03066_),
    .y(_03067_)
  );
  al_aoi21 _08556_ (
    .a(TM0),
    .b(\DFF_1139.Q ),
    .c(TM1),
    .y(_03068_)
  );
  al_nand2 _08557_ (
    .a(_03068_),
    .b(_03067_),
    .y(_03069_)
  );
  al_aoi21ttf _08558_ (
    .a(TM0),
    .b(\DFF_972.Q ),
    .c(TM1),
    .y(_03070_)
  );
  al_and2 _08559_ (
    .a(_03070_),
    .b(_02578_),
    .y(_03071_)
  );
  al_nor3fft _08560_ (
    .a(RESET),
    .b(_03069_),
    .c(_03071_),
    .y(\DFF_1004.D )
  );
  al_or2 _08561_ (
    .a(TM1),
    .b(\DFF_1261.Q ),
    .y(_03072_)
  );
  al_nand2 _08562_ (
    .a(TM1),
    .b(\DFF_1261.Q ),
    .y(_03073_)
  );
  al_nand3 _08563_ (
    .a(\DFF_1293.Q ),
    .b(_03072_),
    .c(_03073_),
    .y(_03074_)
  );
  al_nand2ft _08564_ (
    .a(TM1),
    .b(\DFF_1261.Q ),
    .y(_03075_)
  );
  al_and2ft _08565_ (
    .a(\DFF_1261.Q ),
    .b(TM1),
    .y(_03076_)
  );
  al_and3fft _08566_ (
    .a(\DFF_1293.Q ),
    .b(_03076_),
    .c(_03075_),
    .y(_03077_)
  );
  al_and2ft _08567_ (
    .a(\DFF_1229.Q ),
    .b(\DFF_1197.Q ),
    .y(_03078_)
  );
  al_nand2ft _08568_ (
    .a(\DFF_1197.Q ),
    .b(\DFF_1229.Q ),
    .y(_03079_)
  );
  al_nand2ft _08569_ (
    .a(_03078_),
    .b(_03079_),
    .y(_03080_)
  );
  al_oai21ftf _08570_ (
    .a(_03074_),
    .b(_03077_),
    .c(_03080_),
    .y(_03081_)
  );
  al_nand3ftt _08571_ (
    .a(_03077_),
    .b(_03074_),
    .c(_03080_),
    .y(_03082_)
  );
  al_nand3 _08572_ (
    .a(_00448_),
    .b(_03081_),
    .c(_03082_),
    .y(_03083_)
  );
  al_aoi21 _08573_ (
    .a(TM0),
    .b(\DFF_1138.Q ),
    .c(TM1),
    .y(_03084_)
  );
  al_nand2 _08574_ (
    .a(_03084_),
    .b(_03083_),
    .y(_03085_)
  );
  al_aoi21ttf _08575_ (
    .a(TM0),
    .b(\DFF_973.Q ),
    .c(TM1),
    .y(_03086_)
  );
  al_and2 _08576_ (
    .a(_03086_),
    .b(_02594_),
    .y(_03087_)
  );
  al_nor3fft _08577_ (
    .a(RESET),
    .b(_03085_),
    .c(_03087_),
    .y(\DFF_1005.D )
  );
  al_or2 _08578_ (
    .a(TM1),
    .b(\DFF_1262.Q ),
    .y(_03088_)
  );
  al_nand2 _08579_ (
    .a(TM1),
    .b(\DFF_1262.Q ),
    .y(_03089_)
  );
  al_nand3 _08580_ (
    .a(\DFF_1294.Q ),
    .b(_03088_),
    .c(_03089_),
    .y(_03090_)
  );
  al_nand2ft _08581_ (
    .a(TM1),
    .b(\DFF_1262.Q ),
    .y(_03091_)
  );
  al_and2ft _08582_ (
    .a(\DFF_1262.Q ),
    .b(TM1),
    .y(_03092_)
  );
  al_and3fft _08583_ (
    .a(\DFF_1294.Q ),
    .b(_03092_),
    .c(_03091_),
    .y(_03093_)
  );
  al_and2ft _08584_ (
    .a(\DFF_1230.Q ),
    .b(\DFF_1198.Q ),
    .y(_03094_)
  );
  al_nand2ft _08585_ (
    .a(\DFF_1198.Q ),
    .b(\DFF_1230.Q ),
    .y(_03095_)
  );
  al_nand2ft _08586_ (
    .a(_03094_),
    .b(_03095_),
    .y(_03096_)
  );
  al_oai21ftf _08587_ (
    .a(_03090_),
    .b(_03093_),
    .c(_03096_),
    .y(_03097_)
  );
  al_nand3ftt _08588_ (
    .a(_03093_),
    .b(_03090_),
    .c(_03096_),
    .y(_03098_)
  );
  al_nand3 _08589_ (
    .a(_00448_),
    .b(_03097_),
    .c(_03098_),
    .y(_03099_)
  );
  al_aoi21 _08590_ (
    .a(TM0),
    .b(\DFF_1137.Q ),
    .c(TM1),
    .y(_03100_)
  );
  al_nand2 _08591_ (
    .a(_03100_),
    .b(_03099_),
    .y(_03101_)
  );
  al_aoi21ttf _08592_ (
    .a(TM0),
    .b(\DFF_974.Q ),
    .c(TM1),
    .y(_03102_)
  );
  al_and2 _08593_ (
    .a(_03102_),
    .b(_02610_),
    .y(_03103_)
  );
  al_nor3fft _08594_ (
    .a(RESET),
    .b(_03101_),
    .c(_03103_),
    .y(\DFF_1006.D )
  );
  al_or2 _08595_ (
    .a(TM1),
    .b(\DFF_1263.Q ),
    .y(_03104_)
  );
  al_nand2 _08596_ (
    .a(TM1),
    .b(\DFF_1263.Q ),
    .y(_03105_)
  );
  al_nand3 _08597_ (
    .a(\DFF_1295.Q ),
    .b(_03104_),
    .c(_03105_),
    .y(_03106_)
  );
  al_nand2ft _08598_ (
    .a(TM1),
    .b(\DFF_1263.Q ),
    .y(_03107_)
  );
  al_and2ft _08599_ (
    .a(\DFF_1263.Q ),
    .b(TM1),
    .y(_03108_)
  );
  al_and3fft _08600_ (
    .a(\DFF_1295.Q ),
    .b(_03108_),
    .c(_03107_),
    .y(_03109_)
  );
  al_and2ft _08601_ (
    .a(\DFF_1231.Q ),
    .b(\DFF_1199.Q ),
    .y(_03110_)
  );
  al_nand2ft _08602_ (
    .a(\DFF_1199.Q ),
    .b(\DFF_1231.Q ),
    .y(_03111_)
  );
  al_nand2ft _08603_ (
    .a(_03110_),
    .b(_03111_),
    .y(_03112_)
  );
  al_oai21ftf _08604_ (
    .a(_03106_),
    .b(_03109_),
    .c(_03112_),
    .y(_03113_)
  );
  al_nand3ftt _08605_ (
    .a(_03109_),
    .b(_03106_),
    .c(_03112_),
    .y(_03114_)
  );
  al_nand3 _08606_ (
    .a(_00448_),
    .b(_03113_),
    .c(_03114_),
    .y(_03115_)
  );
  al_aoi21 _08607_ (
    .a(TM0),
    .b(\DFF_1136.Q ),
    .c(TM1),
    .y(_03116_)
  );
  al_nand2 _08608_ (
    .a(_03116_),
    .b(_03115_),
    .y(_03117_)
  );
  al_aoi21ttf _08609_ (
    .a(TM0),
    .b(\DFF_975.Q ),
    .c(TM1),
    .y(_03118_)
  );
  al_and2 _08610_ (
    .a(_03118_),
    .b(_02626_),
    .y(_03119_)
  );
  al_nor3fft _08611_ (
    .a(RESET),
    .b(_03117_),
    .c(_03119_),
    .y(\DFF_1007.D )
  );
  al_nor2 _08612_ (
    .a(\DFF_1232.Q ),
    .b(\DFF_1264.Q ),
    .y(_03120_)
  );
  al_and2 _08613_ (
    .a(\DFF_1232.Q ),
    .b(\DFF_1264.Q ),
    .y(_03121_)
  );
  al_and2ft _08614_ (
    .a(\DFF_1200.Q ),
    .b(\DFF_1296.Q ),
    .y(_03122_)
  );
  al_nand2ft _08615_ (
    .a(\DFF_1296.Q ),
    .b(\DFF_1200.Q ),
    .y(_03123_)
  );
  al_nand2ft _08616_ (
    .a(_03122_),
    .b(_03123_),
    .y(_03124_)
  );
  al_oa21ttf _08617_ (
    .a(_03120_),
    .b(_03121_),
    .c(_03124_),
    .y(_03125_)
  );
  al_nand3fft _08618_ (
    .a(_03120_),
    .b(_03121_),
    .c(_03124_),
    .y(_03126_)
  );
  al_and3fft _08619_ (
    .a(TM0),
    .b(_03125_),
    .c(_03126_),
    .y(_03127_)
  );
  al_nand2 _08620_ (
    .a(TM0),
    .b(\DFF_1135.Q ),
    .y(_03128_)
  );
  al_or3fft _08621_ (
    .a(_01652_),
    .b(_03128_),
    .c(_03127_),
    .y(_03129_)
  );
  al_and2 _08622_ (
    .a(TM0),
    .b(\DFF_976.Q ),
    .y(_03130_)
  );
  al_and3fft _08623_ (
    .a(_03130_),
    .b(_02638_),
    .c(TM1),
    .y(_03131_)
  );
  al_nor3fft _08624_ (
    .a(RESET),
    .b(_03129_),
    .c(_03131_),
    .y(\DFF_1008.D )
  );
  al_nor2 _08625_ (
    .a(\DFF_1233.Q ),
    .b(\DFF_1265.Q ),
    .y(_03132_)
  );
  al_and2 _08626_ (
    .a(\DFF_1233.Q ),
    .b(\DFF_1265.Q ),
    .y(_03133_)
  );
  al_and2ft _08627_ (
    .a(\DFF_1201.Q ),
    .b(\DFF_1297.Q ),
    .y(_03134_)
  );
  al_nand2ft _08628_ (
    .a(\DFF_1297.Q ),
    .b(\DFF_1201.Q ),
    .y(_03135_)
  );
  al_nand2ft _08629_ (
    .a(_03134_),
    .b(_03135_),
    .y(_03136_)
  );
  al_oa21ttf _08630_ (
    .a(_03132_),
    .b(_03133_),
    .c(_03136_),
    .y(_03137_)
  );
  al_nand3fft _08631_ (
    .a(_03132_),
    .b(_03133_),
    .c(_03136_),
    .y(_03138_)
  );
  al_and3fft _08632_ (
    .a(TM0),
    .b(_03137_),
    .c(_03138_),
    .y(_03139_)
  );
  al_nand2 _08633_ (
    .a(TM0),
    .b(\DFF_1134.Q ),
    .y(_03140_)
  );
  al_or3fft _08634_ (
    .a(_01652_),
    .b(_03140_),
    .c(_03139_),
    .y(_03141_)
  );
  al_and2 _08635_ (
    .a(TM0),
    .b(\DFF_977.Q ),
    .y(_03142_)
  );
  al_and3fft _08636_ (
    .a(_03142_),
    .b(_02650_),
    .c(TM1),
    .y(_03143_)
  );
  al_nor3fft _08637_ (
    .a(RESET),
    .b(_03141_),
    .c(_03143_),
    .y(\DFF_1009.D )
  );
  al_nor2 _08638_ (
    .a(\DFF_1234.Q ),
    .b(\DFF_1266.Q ),
    .y(_03144_)
  );
  al_and2 _08639_ (
    .a(\DFF_1234.Q ),
    .b(\DFF_1266.Q ),
    .y(_03145_)
  );
  al_and2ft _08640_ (
    .a(\DFF_1202.Q ),
    .b(\DFF_1298.Q ),
    .y(_03146_)
  );
  al_nand2ft _08641_ (
    .a(\DFF_1298.Q ),
    .b(\DFF_1202.Q ),
    .y(_03147_)
  );
  al_nand2ft _08642_ (
    .a(_03146_),
    .b(_03147_),
    .y(_03148_)
  );
  al_oa21ttf _08643_ (
    .a(_03144_),
    .b(_03145_),
    .c(_03148_),
    .y(_03149_)
  );
  al_nand3fft _08644_ (
    .a(_03144_),
    .b(_03145_),
    .c(_03148_),
    .y(_03150_)
  );
  al_and3fft _08645_ (
    .a(TM0),
    .b(_03149_),
    .c(_03150_),
    .y(_03151_)
  );
  al_nand2 _08646_ (
    .a(TM0),
    .b(\DFF_1133.Q ),
    .y(_03152_)
  );
  al_or3fft _08647_ (
    .a(_01652_),
    .b(_03152_),
    .c(_03151_),
    .y(_03153_)
  );
  al_and2 _08648_ (
    .a(TM0),
    .b(\DFF_978.Q ),
    .y(_03154_)
  );
  al_and3fft _08649_ (
    .a(_03154_),
    .b(_02662_),
    .c(TM1),
    .y(_03155_)
  );
  al_nor3fft _08650_ (
    .a(RESET),
    .b(_03153_),
    .c(_03155_),
    .y(\DFF_1010.D )
  );
  al_nor2 _08651_ (
    .a(\DFF_1235.Q ),
    .b(\DFF_1267.Q ),
    .y(_03156_)
  );
  al_and2 _08652_ (
    .a(\DFF_1235.Q ),
    .b(\DFF_1267.Q ),
    .y(_03157_)
  );
  al_and2ft _08653_ (
    .a(\DFF_1203.Q ),
    .b(\DFF_1299.Q ),
    .y(_03158_)
  );
  al_nand2ft _08654_ (
    .a(\DFF_1299.Q ),
    .b(\DFF_1203.Q ),
    .y(_03159_)
  );
  al_nand2ft _08655_ (
    .a(_03158_),
    .b(_03159_),
    .y(_03160_)
  );
  al_oa21ttf _08656_ (
    .a(_03156_),
    .b(_03157_),
    .c(_03160_),
    .y(_03161_)
  );
  al_nand3fft _08657_ (
    .a(_03156_),
    .b(_03157_),
    .c(_03160_),
    .y(_03162_)
  );
  al_and3fft _08658_ (
    .a(TM0),
    .b(_03161_),
    .c(_03162_),
    .y(_03163_)
  );
  al_nand2 _08659_ (
    .a(TM0),
    .b(\DFF_1132.Q ),
    .y(_03164_)
  );
  al_or3fft _08660_ (
    .a(_01652_),
    .b(_03164_),
    .c(_03163_),
    .y(_03165_)
  );
  al_and2 _08661_ (
    .a(TM0),
    .b(\DFF_979.Q ),
    .y(_03166_)
  );
  al_and3fft _08662_ (
    .a(_03166_),
    .b(_02674_),
    .c(TM1),
    .y(_03167_)
  );
  al_nor3fft _08663_ (
    .a(RESET),
    .b(_03165_),
    .c(_03167_),
    .y(\DFF_1011.D )
  );
  al_nor2 _08664_ (
    .a(\DFF_1236.Q ),
    .b(\DFF_1268.Q ),
    .y(_03168_)
  );
  al_and2 _08665_ (
    .a(\DFF_1236.Q ),
    .b(\DFF_1268.Q ),
    .y(_03169_)
  );
  al_and2ft _08666_ (
    .a(\DFF_1204.Q ),
    .b(\DFF_1300.Q ),
    .y(_03170_)
  );
  al_nand2ft _08667_ (
    .a(\DFF_1300.Q ),
    .b(\DFF_1204.Q ),
    .y(_03171_)
  );
  al_nand2ft _08668_ (
    .a(_03170_),
    .b(_03171_),
    .y(_03172_)
  );
  al_oa21ttf _08669_ (
    .a(_03168_),
    .b(_03169_),
    .c(_03172_),
    .y(_03173_)
  );
  al_nand3fft _08670_ (
    .a(_03168_),
    .b(_03169_),
    .c(_03172_),
    .y(_03174_)
  );
  al_and3fft _08671_ (
    .a(TM0),
    .b(_03173_),
    .c(_03174_),
    .y(_03175_)
  );
  al_nand2 _08672_ (
    .a(TM0),
    .b(\DFF_1131.Q ),
    .y(_03176_)
  );
  al_or3fft _08673_ (
    .a(_01652_),
    .b(_03176_),
    .c(_03175_),
    .y(_03177_)
  );
  al_and2 _08674_ (
    .a(TM0),
    .b(\DFF_980.Q ),
    .y(_03178_)
  );
  al_and3fft _08675_ (
    .a(_03178_),
    .b(_02686_),
    .c(TM1),
    .y(_03179_)
  );
  al_nor3fft _08676_ (
    .a(RESET),
    .b(_03177_),
    .c(_03179_),
    .y(\DFF_1012.D )
  );
  al_nor2 _08677_ (
    .a(\DFF_1237.Q ),
    .b(\DFF_1269.Q ),
    .y(_03180_)
  );
  al_and2 _08678_ (
    .a(\DFF_1237.Q ),
    .b(\DFF_1269.Q ),
    .y(_03181_)
  );
  al_and2ft _08679_ (
    .a(\DFF_1205.Q ),
    .b(\DFF_1301.Q ),
    .y(_03182_)
  );
  al_nand2ft _08680_ (
    .a(\DFF_1301.Q ),
    .b(\DFF_1205.Q ),
    .y(_03183_)
  );
  al_nand2ft _08681_ (
    .a(_03182_),
    .b(_03183_),
    .y(_03184_)
  );
  al_oa21ttf _08682_ (
    .a(_03180_),
    .b(_03181_),
    .c(_03184_),
    .y(_03185_)
  );
  al_nand3fft _08683_ (
    .a(_03180_),
    .b(_03181_),
    .c(_03184_),
    .y(_03186_)
  );
  al_and3fft _08684_ (
    .a(TM0),
    .b(_03185_),
    .c(_03186_),
    .y(_03187_)
  );
  al_nand2 _08685_ (
    .a(TM0),
    .b(\DFF_1130.Q ),
    .y(_03188_)
  );
  al_or3fft _08686_ (
    .a(_01652_),
    .b(_03188_),
    .c(_03187_),
    .y(_03189_)
  );
  al_and2 _08687_ (
    .a(TM0),
    .b(\DFF_981.Q ),
    .y(_03190_)
  );
  al_and3fft _08688_ (
    .a(_03190_),
    .b(_02698_),
    .c(TM1),
    .y(_03191_)
  );
  al_nor3fft _08689_ (
    .a(RESET),
    .b(_03189_),
    .c(_03191_),
    .y(\DFF_1013.D )
  );
  al_nor2 _08690_ (
    .a(\DFF_1238.Q ),
    .b(\DFF_1270.Q ),
    .y(_03192_)
  );
  al_and2 _08691_ (
    .a(\DFF_1238.Q ),
    .b(\DFF_1270.Q ),
    .y(_03193_)
  );
  al_and2ft _08692_ (
    .a(\DFF_1206.Q ),
    .b(\DFF_1302.Q ),
    .y(_03194_)
  );
  al_nand2ft _08693_ (
    .a(\DFF_1302.Q ),
    .b(\DFF_1206.Q ),
    .y(_03195_)
  );
  al_nand2ft _08694_ (
    .a(_03194_),
    .b(_03195_),
    .y(_03196_)
  );
  al_oa21ttf _08695_ (
    .a(_03192_),
    .b(_03193_),
    .c(_03196_),
    .y(_03197_)
  );
  al_nand3fft _08696_ (
    .a(_03192_),
    .b(_03193_),
    .c(_03196_),
    .y(_03198_)
  );
  al_and3fft _08697_ (
    .a(TM0),
    .b(_03197_),
    .c(_03198_),
    .y(_03199_)
  );
  al_nand2 _08698_ (
    .a(TM0),
    .b(\DFF_1129.Q ),
    .y(_03200_)
  );
  al_or3fft _08699_ (
    .a(_01652_),
    .b(_03200_),
    .c(_03199_),
    .y(_03201_)
  );
  al_and2 _08700_ (
    .a(TM0),
    .b(\DFF_982.Q ),
    .y(_03202_)
  );
  al_and3fft _08701_ (
    .a(_03202_),
    .b(_02710_),
    .c(TM1),
    .y(_03203_)
  );
  al_nor3fft _08702_ (
    .a(RESET),
    .b(_03201_),
    .c(_03203_),
    .y(\DFF_1014.D )
  );
  al_nor2 _08703_ (
    .a(\DFF_1239.Q ),
    .b(\DFF_1271.Q ),
    .y(_03204_)
  );
  al_and2 _08704_ (
    .a(\DFF_1239.Q ),
    .b(\DFF_1271.Q ),
    .y(_03205_)
  );
  al_and2ft _08705_ (
    .a(\DFF_1207.Q ),
    .b(\DFF_1303.Q ),
    .y(_03206_)
  );
  al_nand2ft _08706_ (
    .a(\DFF_1303.Q ),
    .b(\DFF_1207.Q ),
    .y(_03207_)
  );
  al_nand2ft _08707_ (
    .a(_03206_),
    .b(_03207_),
    .y(_03208_)
  );
  al_oa21ttf _08708_ (
    .a(_03204_),
    .b(_03205_),
    .c(_03208_),
    .y(_03209_)
  );
  al_nand3fft _08709_ (
    .a(_03204_),
    .b(_03205_),
    .c(_03208_),
    .y(_03210_)
  );
  al_and3fft _08710_ (
    .a(TM0),
    .b(_03209_),
    .c(_03210_),
    .y(_03211_)
  );
  al_nand2 _08711_ (
    .a(TM0),
    .b(\DFF_1128.Q ),
    .y(_03212_)
  );
  al_or3fft _08712_ (
    .a(_01652_),
    .b(_03212_),
    .c(_03211_),
    .y(_03213_)
  );
  al_and2 _08713_ (
    .a(TM0),
    .b(\DFF_983.Q ),
    .y(_03214_)
  );
  al_and3fft _08714_ (
    .a(_03214_),
    .b(_02722_),
    .c(TM1),
    .y(_03215_)
  );
  al_nor3fft _08715_ (
    .a(RESET),
    .b(_03213_),
    .c(_03215_),
    .y(\DFF_1015.D )
  );
  al_nor2 _08716_ (
    .a(\DFF_1240.Q ),
    .b(\DFF_1272.Q ),
    .y(_03216_)
  );
  al_and2 _08717_ (
    .a(\DFF_1240.Q ),
    .b(\DFF_1272.Q ),
    .y(_03217_)
  );
  al_and2ft _08718_ (
    .a(\DFF_1208.Q ),
    .b(\DFF_1304.Q ),
    .y(_03218_)
  );
  al_nand2ft _08719_ (
    .a(\DFF_1304.Q ),
    .b(\DFF_1208.Q ),
    .y(_03219_)
  );
  al_nand2ft _08720_ (
    .a(_03218_),
    .b(_03219_),
    .y(_03220_)
  );
  al_oa21ttf _08721_ (
    .a(_03216_),
    .b(_03217_),
    .c(_03220_),
    .y(_03221_)
  );
  al_nand3fft _08722_ (
    .a(_03216_),
    .b(_03217_),
    .c(_03220_),
    .y(_03222_)
  );
  al_and3fft _08723_ (
    .a(TM0),
    .b(_03221_),
    .c(_03222_),
    .y(_03223_)
  );
  al_nand2 _08724_ (
    .a(TM0),
    .b(\DFF_1127.Q ),
    .y(_03224_)
  );
  al_or3fft _08725_ (
    .a(_01652_),
    .b(_03224_),
    .c(_03223_),
    .y(_03225_)
  );
  al_and2 _08726_ (
    .a(TM0),
    .b(\DFF_984.Q ),
    .y(_03226_)
  );
  al_and3fft _08727_ (
    .a(_03226_),
    .b(_02734_),
    .c(TM1),
    .y(_03227_)
  );
  al_nor3fft _08728_ (
    .a(RESET),
    .b(_03225_),
    .c(_03227_),
    .y(\DFF_1016.D )
  );
  al_nor2 _08729_ (
    .a(\DFF_1241.Q ),
    .b(\DFF_1273.Q ),
    .y(_03228_)
  );
  al_and2 _08730_ (
    .a(\DFF_1241.Q ),
    .b(\DFF_1273.Q ),
    .y(_03229_)
  );
  al_and2ft _08731_ (
    .a(\DFF_1209.Q ),
    .b(\DFF_1305.Q ),
    .y(_03230_)
  );
  al_nand2ft _08732_ (
    .a(\DFF_1305.Q ),
    .b(\DFF_1209.Q ),
    .y(_03231_)
  );
  al_nand2ft _08733_ (
    .a(_03230_),
    .b(_03231_),
    .y(_03232_)
  );
  al_oa21ttf _08734_ (
    .a(_03228_),
    .b(_03229_),
    .c(_03232_),
    .y(_03233_)
  );
  al_nand3fft _08735_ (
    .a(_03228_),
    .b(_03229_),
    .c(_03232_),
    .y(_03234_)
  );
  al_and3fft _08736_ (
    .a(TM0),
    .b(_03233_),
    .c(_03234_),
    .y(_03235_)
  );
  al_nand2 _08737_ (
    .a(TM0),
    .b(\DFF_1126.Q ),
    .y(_03236_)
  );
  al_or3fft _08738_ (
    .a(_01652_),
    .b(_03236_),
    .c(_03235_),
    .y(_03237_)
  );
  al_and2 _08739_ (
    .a(TM0),
    .b(\DFF_985.Q ),
    .y(_03238_)
  );
  al_and3fft _08740_ (
    .a(_03238_),
    .b(_02746_),
    .c(TM1),
    .y(_03239_)
  );
  al_nor3fft _08741_ (
    .a(RESET),
    .b(_03237_),
    .c(_03239_),
    .y(\DFF_1017.D )
  );
  al_nor2 _08742_ (
    .a(\DFF_1242.Q ),
    .b(\DFF_1274.Q ),
    .y(_03240_)
  );
  al_and2 _08743_ (
    .a(\DFF_1242.Q ),
    .b(\DFF_1274.Q ),
    .y(_03241_)
  );
  al_and2ft _08744_ (
    .a(\DFF_1210.Q ),
    .b(\DFF_1306.Q ),
    .y(_03242_)
  );
  al_nand2ft _08745_ (
    .a(\DFF_1306.Q ),
    .b(\DFF_1210.Q ),
    .y(_03243_)
  );
  al_nand2ft _08746_ (
    .a(_03242_),
    .b(_03243_),
    .y(_03244_)
  );
  al_oa21ttf _08747_ (
    .a(_03240_),
    .b(_03241_),
    .c(_03244_),
    .y(_03245_)
  );
  al_nand3fft _08748_ (
    .a(_03240_),
    .b(_03241_),
    .c(_03244_),
    .y(_03246_)
  );
  al_and3fft _08749_ (
    .a(TM0),
    .b(_03245_),
    .c(_03246_),
    .y(_03247_)
  );
  al_nand2 _08750_ (
    .a(TM0),
    .b(\DFF_1125.Q ),
    .y(_03248_)
  );
  al_or3fft _08751_ (
    .a(_01652_),
    .b(_03248_),
    .c(_03247_),
    .y(_03249_)
  );
  al_and2 _08752_ (
    .a(TM0),
    .b(\DFF_986.Q ),
    .y(_03250_)
  );
  al_and3fft _08753_ (
    .a(_03250_),
    .b(_02758_),
    .c(TM1),
    .y(_03251_)
  );
  al_nor3fft _08754_ (
    .a(RESET),
    .b(_03249_),
    .c(_03251_),
    .y(\DFF_1018.D )
  );
  al_nor2 _08755_ (
    .a(\DFF_1243.Q ),
    .b(\DFF_1275.Q ),
    .y(_03252_)
  );
  al_and2 _08756_ (
    .a(\DFF_1243.Q ),
    .b(\DFF_1275.Q ),
    .y(_03253_)
  );
  al_and2ft _08757_ (
    .a(\DFF_1211.Q ),
    .b(\DFF_1307.Q ),
    .y(_03254_)
  );
  al_nand2ft _08758_ (
    .a(\DFF_1307.Q ),
    .b(\DFF_1211.Q ),
    .y(_03255_)
  );
  al_nand2ft _08759_ (
    .a(_03254_),
    .b(_03255_),
    .y(_03256_)
  );
  al_oa21ttf _08760_ (
    .a(_03252_),
    .b(_03253_),
    .c(_03256_),
    .y(_03257_)
  );
  al_nand3fft _08761_ (
    .a(_03252_),
    .b(_03253_),
    .c(_03256_),
    .y(_03258_)
  );
  al_and3fft _08762_ (
    .a(TM0),
    .b(_03257_),
    .c(_03258_),
    .y(_03259_)
  );
  al_nand2 _08763_ (
    .a(TM0),
    .b(\DFF_1124.Q ),
    .y(_03260_)
  );
  al_or3fft _08764_ (
    .a(_01652_),
    .b(_03260_),
    .c(_03259_),
    .y(_03261_)
  );
  al_and2 _08765_ (
    .a(TM0),
    .b(\DFF_987.Q ),
    .y(_03262_)
  );
  al_and3fft _08766_ (
    .a(_03262_),
    .b(_02770_),
    .c(TM1),
    .y(_03263_)
  );
  al_nor3fft _08767_ (
    .a(RESET),
    .b(_03261_),
    .c(_03263_),
    .y(\DFF_1019.D )
  );
  al_nor2 _08768_ (
    .a(\DFF_1244.Q ),
    .b(\DFF_1276.Q ),
    .y(_03264_)
  );
  al_and2 _08769_ (
    .a(\DFF_1244.Q ),
    .b(\DFF_1276.Q ),
    .y(_03265_)
  );
  al_and2ft _08770_ (
    .a(\DFF_1212.Q ),
    .b(\DFF_1308.Q ),
    .y(_03266_)
  );
  al_nand2ft _08771_ (
    .a(\DFF_1308.Q ),
    .b(\DFF_1212.Q ),
    .y(_03267_)
  );
  al_nand2ft _08772_ (
    .a(_03266_),
    .b(_03267_),
    .y(_03268_)
  );
  al_oa21ttf _08773_ (
    .a(_03264_),
    .b(_03265_),
    .c(_03268_),
    .y(_03269_)
  );
  al_nand3fft _08774_ (
    .a(_03264_),
    .b(_03265_),
    .c(_03268_),
    .y(_03270_)
  );
  al_and3fft _08775_ (
    .a(TM0),
    .b(_03269_),
    .c(_03270_),
    .y(_03271_)
  );
  al_nand2 _08776_ (
    .a(TM0),
    .b(\DFF_1123.Q ),
    .y(_03272_)
  );
  al_or3fft _08777_ (
    .a(_01652_),
    .b(_03272_),
    .c(_03271_),
    .y(_03273_)
  );
  al_and2 _08778_ (
    .a(TM0),
    .b(\DFF_988.Q ),
    .y(_03274_)
  );
  al_and3fft _08779_ (
    .a(_03274_),
    .b(_02782_),
    .c(TM1),
    .y(_03275_)
  );
  al_nor3fft _08780_ (
    .a(RESET),
    .b(_03273_),
    .c(_03275_),
    .y(\DFF_1020.D )
  );
  al_nor2 _08781_ (
    .a(\DFF_1245.Q ),
    .b(\DFF_1277.Q ),
    .y(_03276_)
  );
  al_and2 _08782_ (
    .a(\DFF_1245.Q ),
    .b(\DFF_1277.Q ),
    .y(_03277_)
  );
  al_and2ft _08783_ (
    .a(\DFF_1213.Q ),
    .b(\DFF_1309.Q ),
    .y(_03278_)
  );
  al_nand2ft _08784_ (
    .a(\DFF_1309.Q ),
    .b(\DFF_1213.Q ),
    .y(_03279_)
  );
  al_nand2ft _08785_ (
    .a(_03278_),
    .b(_03279_),
    .y(_03280_)
  );
  al_oa21ttf _08786_ (
    .a(_03276_),
    .b(_03277_),
    .c(_03280_),
    .y(_03281_)
  );
  al_nand3fft _08787_ (
    .a(_03276_),
    .b(_03277_),
    .c(_03280_),
    .y(_03282_)
  );
  al_and3fft _08788_ (
    .a(TM0),
    .b(_03281_),
    .c(_03282_),
    .y(_03283_)
  );
  al_nand2 _08789_ (
    .a(TM0),
    .b(\DFF_1122.Q ),
    .y(_03284_)
  );
  al_or3fft _08790_ (
    .a(_01652_),
    .b(_03284_),
    .c(_03283_),
    .y(_03285_)
  );
  al_and2 _08791_ (
    .a(TM0),
    .b(\DFF_989.Q ),
    .y(_03286_)
  );
  al_and3fft _08792_ (
    .a(_03286_),
    .b(_02794_),
    .c(TM1),
    .y(_03287_)
  );
  al_nor3fft _08793_ (
    .a(RESET),
    .b(_03285_),
    .c(_03287_),
    .y(\DFF_1021.D )
  );
  al_nor2 _08794_ (
    .a(\DFF_1246.Q ),
    .b(\DFF_1278.Q ),
    .y(_03288_)
  );
  al_and2 _08795_ (
    .a(\DFF_1246.Q ),
    .b(\DFF_1278.Q ),
    .y(_03289_)
  );
  al_and2ft _08796_ (
    .a(\DFF_1214.Q ),
    .b(\DFF_1310.Q ),
    .y(_03290_)
  );
  al_nand2ft _08797_ (
    .a(\DFF_1310.Q ),
    .b(\DFF_1214.Q ),
    .y(_03291_)
  );
  al_nand2ft _08798_ (
    .a(_03290_),
    .b(_03291_),
    .y(_03292_)
  );
  al_oa21ttf _08799_ (
    .a(_03288_),
    .b(_03289_),
    .c(_03292_),
    .y(_03293_)
  );
  al_nand3fft _08800_ (
    .a(_03288_),
    .b(_03289_),
    .c(_03292_),
    .y(_03294_)
  );
  al_and3fft _08801_ (
    .a(TM0),
    .b(_03293_),
    .c(_03294_),
    .y(_03295_)
  );
  al_nand2 _08802_ (
    .a(TM0),
    .b(\DFF_1121.Q ),
    .y(_03296_)
  );
  al_or3fft _08803_ (
    .a(_01652_),
    .b(_03296_),
    .c(_03295_),
    .y(_03297_)
  );
  al_and2 _08804_ (
    .a(TM0),
    .b(\DFF_990.Q ),
    .y(_03298_)
  );
  al_and3fft _08805_ (
    .a(_03298_),
    .b(_02806_),
    .c(TM1),
    .y(_03299_)
  );
  al_nor3fft _08806_ (
    .a(RESET),
    .b(_03297_),
    .c(_03299_),
    .y(\DFF_1022.D )
  );
  al_nor2 _08807_ (
    .a(\DFF_1247.Q ),
    .b(\DFF_1279.Q ),
    .y(_03300_)
  );
  al_and2 _08808_ (
    .a(\DFF_1247.Q ),
    .b(\DFF_1279.Q ),
    .y(_03301_)
  );
  al_and2ft _08809_ (
    .a(\DFF_1215.Q ),
    .b(\DFF_1311.Q ),
    .y(_03302_)
  );
  al_nand2ft _08810_ (
    .a(\DFF_1311.Q ),
    .b(\DFF_1215.Q ),
    .y(_03303_)
  );
  al_nand2ft _08811_ (
    .a(_03302_),
    .b(_03303_),
    .y(_03304_)
  );
  al_oa21ttf _08812_ (
    .a(_03300_),
    .b(_03301_),
    .c(_03304_),
    .y(_03305_)
  );
  al_nand3fft _08813_ (
    .a(_03300_),
    .b(_03301_),
    .c(_03304_),
    .y(_03306_)
  );
  al_and3fft _08814_ (
    .a(TM0),
    .b(_03305_),
    .c(_03306_),
    .y(_03307_)
  );
  al_nand2 _08815_ (
    .a(TM0),
    .b(\DFF_1120.Q ),
    .y(_03308_)
  );
  al_or3fft _08816_ (
    .a(_01652_),
    .b(_03308_),
    .c(_03307_),
    .y(_03309_)
  );
  al_and2 _08817_ (
    .a(TM0),
    .b(\DFF_991.Q ),
    .y(_03310_)
  );
  al_and3fft _08818_ (
    .a(_03310_),
    .b(_02818_),
    .c(TM1),
    .y(_03311_)
  );
  al_nor3fft _08819_ (
    .a(RESET),
    .b(_03309_),
    .c(_03311_),
    .y(\DFF_1023.D )
  );
  al_and2 _08820_ (
    .a(RESET),
    .b(\DFF_992.Q ),
    .y(\DFF_1024.D )
  );
  al_and2 _08821_ (
    .a(RESET),
    .b(\DFF_993.Q ),
    .y(\DFF_1025.D )
  );
  al_and2 _08822_ (
    .a(RESET),
    .b(\DFF_994.Q ),
    .y(\DFF_1026.D )
  );
  al_and2 _08823_ (
    .a(RESET),
    .b(\DFF_995.Q ),
    .y(\DFF_1027.D )
  );
  al_and2 _08824_ (
    .a(RESET),
    .b(\DFF_996.Q ),
    .y(\DFF_1028.D )
  );
  al_and2 _08825_ (
    .a(RESET),
    .b(\DFF_997.Q ),
    .y(\DFF_1029.D )
  );
  al_and2 _08826_ (
    .a(RESET),
    .b(\DFF_998.Q ),
    .y(\DFF_1030.D )
  );
  al_and2 _08827_ (
    .a(RESET),
    .b(\DFF_999.Q ),
    .y(\DFF_1031.D )
  );
  al_and2 _08828_ (
    .a(RESET),
    .b(\DFF_1000.Q ),
    .y(\DFF_1032.D )
  );
  al_and2 _08829_ (
    .a(RESET),
    .b(\DFF_1001.Q ),
    .y(\DFF_1033.D )
  );
  al_and2 _08830_ (
    .a(RESET),
    .b(\DFF_1002.Q ),
    .y(\DFF_1034.D )
  );
  al_and2 _08831_ (
    .a(RESET),
    .b(\DFF_1003.Q ),
    .y(\DFF_1035.D )
  );
  al_and2 _08832_ (
    .a(RESET),
    .b(\DFF_1004.Q ),
    .y(\DFF_1036.D )
  );
  al_and2 _08833_ (
    .a(RESET),
    .b(\DFF_1005.Q ),
    .y(\DFF_1037.D )
  );
  al_and2 _08834_ (
    .a(RESET),
    .b(\DFF_1006.Q ),
    .y(\DFF_1038.D )
  );
  al_and2 _08835_ (
    .a(RESET),
    .b(\DFF_1007.Q ),
    .y(\DFF_1039.D )
  );
  al_and2 _08836_ (
    .a(RESET),
    .b(\DFF_1008.Q ),
    .y(\DFF_1040.D )
  );
  al_and2 _08837_ (
    .a(RESET),
    .b(\DFF_1009.Q ),
    .y(\DFF_1041.D )
  );
  al_and2 _08838_ (
    .a(RESET),
    .b(\DFF_1010.Q ),
    .y(\DFF_1042.D )
  );
  al_and2 _08839_ (
    .a(RESET),
    .b(\DFF_1011.Q ),
    .y(\DFF_1043.D )
  );
  al_and2 _08840_ (
    .a(RESET),
    .b(\DFF_1012.Q ),
    .y(\DFF_1044.D )
  );
  al_and2 _08841_ (
    .a(RESET),
    .b(\DFF_1013.Q ),
    .y(\DFF_1045.D )
  );
  al_and2 _08842_ (
    .a(RESET),
    .b(\DFF_1014.Q ),
    .y(\DFF_1046.D )
  );
  al_and2 _08843_ (
    .a(RESET),
    .b(\DFF_1015.Q ),
    .y(\DFF_1047.D )
  );
  al_and2 _08844_ (
    .a(RESET),
    .b(\DFF_1016.Q ),
    .y(\DFF_1048.D )
  );
  al_and2 _08845_ (
    .a(RESET),
    .b(\DFF_1017.Q ),
    .y(\DFF_1049.D )
  );
  al_and2 _08846_ (
    .a(RESET),
    .b(\DFF_1018.Q ),
    .y(\DFF_1050.D )
  );
  al_and2 _08847_ (
    .a(RESET),
    .b(\DFF_1019.Q ),
    .y(\DFF_1051.D )
  );
  al_and2 _08848_ (
    .a(RESET),
    .b(\DFF_1020.Q ),
    .y(\DFF_1052.D )
  );
  al_and2 _08849_ (
    .a(RESET),
    .b(\DFF_1021.Q ),
    .y(\DFF_1053.D )
  );
  al_and2 _08850_ (
    .a(RESET),
    .b(\DFF_1022.Q ),
    .y(\DFF_1054.D )
  );
  al_and2 _08851_ (
    .a(RESET),
    .b(\DFF_1023.Q ),
    .y(\DFF_1055.D )
  );
  al_and2 _08852_ (
    .a(RESET),
    .b(\DFF_1024.Q ),
    .y(\DFF_1056.D )
  );
  al_and2 _08853_ (
    .a(RESET),
    .b(\DFF_1025.Q ),
    .y(\DFF_1057.D )
  );
  al_and2 _08854_ (
    .a(RESET),
    .b(\DFF_1026.Q ),
    .y(\DFF_1058.D )
  );
  al_and2 _08855_ (
    .a(RESET),
    .b(\DFF_1027.Q ),
    .y(\DFF_1059.D )
  );
  al_and2 _08856_ (
    .a(RESET),
    .b(\DFF_1028.Q ),
    .y(\DFF_1060.D )
  );
  al_and2 _08857_ (
    .a(RESET),
    .b(\DFF_1029.Q ),
    .y(\DFF_1061.D )
  );
  al_and2 _08858_ (
    .a(RESET),
    .b(\DFF_1030.Q ),
    .y(\DFF_1062.D )
  );
  al_and2 _08859_ (
    .a(RESET),
    .b(\DFF_1031.Q ),
    .y(\DFF_1063.D )
  );
  al_and2 _08860_ (
    .a(RESET),
    .b(\DFF_1032.Q ),
    .y(\DFF_1064.D )
  );
  al_and2 _08861_ (
    .a(RESET),
    .b(\DFF_1033.Q ),
    .y(\DFF_1065.D )
  );
  al_and2 _08862_ (
    .a(RESET),
    .b(\DFF_1034.Q ),
    .y(\DFF_1066.D )
  );
  al_and2 _08863_ (
    .a(RESET),
    .b(\DFF_1035.Q ),
    .y(\DFF_1067.D )
  );
  al_and2 _08864_ (
    .a(RESET),
    .b(\DFF_1036.Q ),
    .y(\DFF_1068.D )
  );
  al_and2 _08865_ (
    .a(RESET),
    .b(\DFF_1037.Q ),
    .y(\DFF_1069.D )
  );
  al_and2 _08866_ (
    .a(RESET),
    .b(\DFF_1038.Q ),
    .y(\DFF_1070.D )
  );
  al_and2 _08867_ (
    .a(RESET),
    .b(\DFF_1039.Q ),
    .y(\DFF_1071.D )
  );
  al_and2 _08868_ (
    .a(RESET),
    .b(\DFF_1040.Q ),
    .y(\DFF_1072.D )
  );
  al_and2 _08869_ (
    .a(RESET),
    .b(\DFF_1041.Q ),
    .y(\DFF_1073.D )
  );
  al_and2 _08870_ (
    .a(RESET),
    .b(\DFF_1042.Q ),
    .y(\DFF_1074.D )
  );
  al_and2 _08871_ (
    .a(RESET),
    .b(\DFF_1043.Q ),
    .y(\DFF_1075.D )
  );
  al_and2 _08872_ (
    .a(RESET),
    .b(\DFF_1044.Q ),
    .y(\DFF_1076.D )
  );
  al_and2 _08873_ (
    .a(RESET),
    .b(\DFF_1045.Q ),
    .y(\DFF_1077.D )
  );
  al_and2 _08874_ (
    .a(RESET),
    .b(\DFF_1046.Q ),
    .y(\DFF_1078.D )
  );
  al_and2 _08875_ (
    .a(RESET),
    .b(\DFF_1047.Q ),
    .y(\DFF_1079.D )
  );
  al_and2 _08876_ (
    .a(RESET),
    .b(\DFF_1048.Q ),
    .y(\DFF_1080.D )
  );
  al_and2 _08877_ (
    .a(RESET),
    .b(\DFF_1049.Q ),
    .y(\DFF_1081.D )
  );
  al_and2 _08878_ (
    .a(RESET),
    .b(\DFF_1050.Q ),
    .y(\DFF_1082.D )
  );
  al_and2 _08879_ (
    .a(RESET),
    .b(\DFF_1051.Q ),
    .y(\DFF_1083.D )
  );
  al_and2 _08880_ (
    .a(RESET),
    .b(\DFF_1052.Q ),
    .y(\DFF_1084.D )
  );
  al_and2 _08881_ (
    .a(RESET),
    .b(\DFF_1053.Q ),
    .y(\DFF_1085.D )
  );
  al_and2 _08882_ (
    .a(RESET),
    .b(\DFF_1054.Q ),
    .y(\DFF_1086.D )
  );
  al_and2 _08883_ (
    .a(RESET),
    .b(\DFF_1055.Q ),
    .y(\DFF_1087.D )
  );
  al_and2 _08884_ (
    .a(RESET),
    .b(\DFF_1056.Q ),
    .y(\DFF_1088.D )
  );
  al_and2 _08885_ (
    .a(RESET),
    .b(\DFF_1057.Q ),
    .y(\DFF_1089.D )
  );
  al_and2 _08886_ (
    .a(RESET),
    .b(\DFF_1058.Q ),
    .y(\DFF_1090.D )
  );
  al_and2 _08887_ (
    .a(RESET),
    .b(\DFF_1059.Q ),
    .y(\DFF_1091.D )
  );
  al_and2 _08888_ (
    .a(RESET),
    .b(\DFF_1060.Q ),
    .y(\DFF_1092.D )
  );
  al_and2 _08889_ (
    .a(RESET),
    .b(\DFF_1061.Q ),
    .y(\DFF_1093.D )
  );
  al_and2 _08890_ (
    .a(RESET),
    .b(\DFF_1062.Q ),
    .y(\DFF_1094.D )
  );
  al_and2 _08891_ (
    .a(RESET),
    .b(\DFF_1063.Q ),
    .y(\DFF_1095.D )
  );
  al_and2 _08892_ (
    .a(RESET),
    .b(\DFF_1064.Q ),
    .y(\DFF_1096.D )
  );
  al_and2 _08893_ (
    .a(RESET),
    .b(\DFF_1065.Q ),
    .y(\DFF_1097.D )
  );
  al_and2 _08894_ (
    .a(RESET),
    .b(\DFF_1066.Q ),
    .y(\DFF_1098.D )
  );
  al_and2 _08895_ (
    .a(RESET),
    .b(\DFF_1067.Q ),
    .y(\DFF_1099.D )
  );
  al_and2 _08896_ (
    .a(RESET),
    .b(\DFF_1068.Q ),
    .y(\DFF_1100.D )
  );
  al_and2 _08897_ (
    .a(RESET),
    .b(\DFF_1069.Q ),
    .y(\DFF_1101.D )
  );
  al_and2 _08898_ (
    .a(RESET),
    .b(\DFF_1070.Q ),
    .y(\DFF_1102.D )
  );
  al_and2 _08899_ (
    .a(RESET),
    .b(\DFF_1071.Q ),
    .y(\DFF_1103.D )
  );
  al_and2 _08900_ (
    .a(RESET),
    .b(\DFF_1072.Q ),
    .y(\DFF_1104.D )
  );
  al_and2 _08901_ (
    .a(RESET),
    .b(\DFF_1073.Q ),
    .y(\DFF_1105.D )
  );
  al_and2 _08902_ (
    .a(RESET),
    .b(\DFF_1074.Q ),
    .y(\DFF_1106.D )
  );
  al_and2 _08903_ (
    .a(RESET),
    .b(\DFF_1075.Q ),
    .y(\DFF_1107.D )
  );
  al_and2 _08904_ (
    .a(RESET),
    .b(\DFF_1076.Q ),
    .y(\DFF_1108.D )
  );
  al_and2 _08905_ (
    .a(RESET),
    .b(\DFF_1077.Q ),
    .y(\DFF_1109.D )
  );
  al_and2 _08906_ (
    .a(RESET),
    .b(\DFF_1078.Q ),
    .y(\DFF_1110.D )
  );
  al_and2 _08907_ (
    .a(RESET),
    .b(\DFF_1079.Q ),
    .y(\DFF_1111.D )
  );
  al_and2 _08908_ (
    .a(RESET),
    .b(\DFF_1080.Q ),
    .y(\DFF_1112.D )
  );
  al_and2 _08909_ (
    .a(RESET),
    .b(\DFF_1081.Q ),
    .y(\DFF_1113.D )
  );
  al_and2 _08910_ (
    .a(RESET),
    .b(\DFF_1082.Q ),
    .y(\DFF_1114.D )
  );
  al_and2 _08911_ (
    .a(RESET),
    .b(\DFF_1083.Q ),
    .y(\DFF_1115.D )
  );
  al_and2 _08912_ (
    .a(RESET),
    .b(\DFF_1084.Q ),
    .y(\DFF_1116.D )
  );
  al_and2 _08913_ (
    .a(RESET),
    .b(\DFF_1085.Q ),
    .y(\DFF_1117.D )
  );
  al_and2 _08914_ (
    .a(RESET),
    .b(\DFF_1086.Q ),
    .y(\DFF_1118.D )
  );
  al_and2 _08915_ (
    .a(RESET),
    .b(\DFF_1087.Q ),
    .y(\DFF_1119.D )
  );
  al_oa21ftt _08916_ (
    .a(\DFF_1119.Q ),
    .b(\DFF_1151.Q ),
    .c(RESET),
    .y(_03312_)
  );
  al_aoi21ftf _08917_ (
    .a(\DFF_1119.Q ),
    .b(\DFF_1151.Q ),
    .c(_03312_),
    .y(\DFF_1120.D )
  );
  al_oa21ftt _08918_ (
    .a(\DFF_1118.Q ),
    .b(\DFF_1120.Q ),
    .c(RESET),
    .y(_03313_)
  );
  al_aoi21ftf _08919_ (
    .a(\DFF_1118.Q ),
    .b(\DFF_1120.Q ),
    .c(_03313_),
    .y(\DFF_1121.D )
  );
  al_oa21ftt _08920_ (
    .a(\DFF_1117.Q ),
    .b(\DFF_1121.Q ),
    .c(RESET),
    .y(_03314_)
  );
  al_aoi21ftf _08921_ (
    .a(\DFF_1117.Q ),
    .b(\DFF_1121.Q ),
    .c(_03314_),
    .y(\DFF_1122.D )
  );
  al_oa21ftt _08922_ (
    .a(\DFF_1116.Q ),
    .b(\DFF_1122.Q ),
    .c(RESET),
    .y(_03315_)
  );
  al_aoi21ftf _08923_ (
    .a(\DFF_1116.Q ),
    .b(\DFF_1122.Q ),
    .c(_03315_),
    .y(\DFF_1123.D )
  );
  al_nand2ft _08924_ (
    .a(\DFF_1115.Q ),
    .b(\DFF_1123.Q ),
    .y(_03316_)
  );
  al_nand2ft _08925_ (
    .a(\DFF_1123.Q ),
    .b(\DFF_1115.Q ),
    .y(_03317_)
  );
  al_ao21ttf _08926_ (
    .a(_03316_),
    .b(_03317_),
    .c(\DFF_1151.Q ),
    .y(_03318_)
  );
  al_nand3ftt _08927_ (
    .a(\DFF_1151.Q ),
    .b(_03316_),
    .c(_03317_),
    .y(_03319_)
  );
  al_aoi21 _08928_ (
    .a(_03319_),
    .b(_03318_),
    .c(_00451_),
    .y(\DFF_1124.D )
  );
  al_oa21ftt _08929_ (
    .a(\DFF_1114.Q ),
    .b(\DFF_1124.Q ),
    .c(RESET),
    .y(_03320_)
  );
  al_aoi21ftf _08930_ (
    .a(\DFF_1114.Q ),
    .b(\DFF_1124.Q ),
    .c(_03320_),
    .y(\DFF_1125.D )
  );
  al_oa21ftt _08931_ (
    .a(\DFF_1113.Q ),
    .b(\DFF_1125.Q ),
    .c(RESET),
    .y(_03321_)
  );
  al_aoi21ftf _08932_ (
    .a(\DFF_1113.Q ),
    .b(\DFF_1125.Q ),
    .c(_03321_),
    .y(\DFF_1126.D )
  );
  al_oa21ftt _08933_ (
    .a(\DFF_1112.Q ),
    .b(\DFF_1126.Q ),
    .c(RESET),
    .y(_03322_)
  );
  al_aoi21ftf _08934_ (
    .a(\DFF_1112.Q ),
    .b(\DFF_1126.Q ),
    .c(_03322_),
    .y(\DFF_1127.D )
  );
  al_oa21ftt _08935_ (
    .a(\DFF_1111.Q ),
    .b(\DFF_1127.Q ),
    .c(RESET),
    .y(_03323_)
  );
  al_aoi21ftf _08936_ (
    .a(\DFF_1111.Q ),
    .b(\DFF_1127.Q ),
    .c(_03323_),
    .y(\DFF_1128.D )
  );
  al_oa21ftt _08937_ (
    .a(\DFF_1110.Q ),
    .b(\DFF_1128.Q ),
    .c(RESET),
    .y(_03324_)
  );
  al_aoi21ftf _08938_ (
    .a(\DFF_1110.Q ),
    .b(\DFF_1128.Q ),
    .c(_03324_),
    .y(\DFF_1129.D )
  );
  al_oa21ftt _08939_ (
    .a(\DFF_1109.Q ),
    .b(\DFF_1129.Q ),
    .c(RESET),
    .y(_03325_)
  );
  al_aoi21ftf _08940_ (
    .a(\DFF_1109.Q ),
    .b(\DFF_1129.Q ),
    .c(_03325_),
    .y(\DFF_1130.D )
  );
  al_nand2ft _08941_ (
    .a(\DFF_1108.Q ),
    .b(\DFF_1130.Q ),
    .y(_03326_)
  );
  al_nand2ft _08942_ (
    .a(\DFF_1130.Q ),
    .b(\DFF_1108.Q ),
    .y(_03327_)
  );
  al_ao21ttf _08943_ (
    .a(_03326_),
    .b(_03327_),
    .c(\DFF_1151.Q ),
    .y(_03328_)
  );
  al_nand3ftt _08944_ (
    .a(\DFF_1151.Q ),
    .b(_03326_),
    .c(_03327_),
    .y(_03329_)
  );
  al_aoi21 _08945_ (
    .a(_03329_),
    .b(_03328_),
    .c(_00451_),
    .y(\DFF_1131.D )
  );
  al_oa21ftt _08946_ (
    .a(\DFF_1107.Q ),
    .b(\DFF_1131.Q ),
    .c(RESET),
    .y(_03330_)
  );
  al_aoi21ftf _08947_ (
    .a(\DFF_1107.Q ),
    .b(\DFF_1131.Q ),
    .c(_03330_),
    .y(\DFF_1132.D )
  );
  al_oa21ftt _08948_ (
    .a(\DFF_1106.Q ),
    .b(\DFF_1132.Q ),
    .c(RESET),
    .y(_03331_)
  );
  al_aoi21ftf _08949_ (
    .a(\DFF_1106.Q ),
    .b(\DFF_1132.Q ),
    .c(_03331_),
    .y(\DFF_1133.D )
  );
  al_oa21ftt _08950_ (
    .a(\DFF_1105.Q ),
    .b(\DFF_1133.Q ),
    .c(RESET),
    .y(_03332_)
  );
  al_aoi21ftf _08951_ (
    .a(\DFF_1105.Q ),
    .b(\DFF_1133.Q ),
    .c(_03332_),
    .y(\DFF_1134.D )
  );
  al_oa21ftt _08952_ (
    .a(\DFF_1104.Q ),
    .b(\DFF_1134.Q ),
    .c(RESET),
    .y(_03333_)
  );
  al_aoi21ftf _08953_ (
    .a(\DFF_1104.Q ),
    .b(\DFF_1134.Q ),
    .c(_03333_),
    .y(\DFF_1135.D )
  );
  al_nand2ft _08954_ (
    .a(\DFF_1103.Q ),
    .b(\DFF_1135.Q ),
    .y(_03334_)
  );
  al_nand2ft _08955_ (
    .a(\DFF_1135.Q ),
    .b(\DFF_1103.Q ),
    .y(_03335_)
  );
  al_ao21ttf _08956_ (
    .a(_03334_),
    .b(_03335_),
    .c(\DFF_1151.Q ),
    .y(_03336_)
  );
  al_nand3ftt _08957_ (
    .a(\DFF_1151.Q ),
    .b(_03334_),
    .c(_03335_),
    .y(_03337_)
  );
  al_aoi21 _08958_ (
    .a(_03337_),
    .b(_03336_),
    .c(_00451_),
    .y(\DFF_1136.D )
  );
  al_oa21ftt _08959_ (
    .a(\DFF_1102.Q ),
    .b(\DFF_1136.Q ),
    .c(RESET),
    .y(_03338_)
  );
  al_aoi21ftf _08960_ (
    .a(\DFF_1102.Q ),
    .b(\DFF_1136.Q ),
    .c(_03338_),
    .y(\DFF_1137.D )
  );
  al_oa21ftt _08961_ (
    .a(\DFF_1101.Q ),
    .b(\DFF_1137.Q ),
    .c(RESET),
    .y(_03339_)
  );
  al_aoi21ftf _08962_ (
    .a(\DFF_1101.Q ),
    .b(\DFF_1137.Q ),
    .c(_03339_),
    .y(\DFF_1138.D )
  );
  al_oa21ftt _08963_ (
    .a(\DFF_1100.Q ),
    .b(\DFF_1138.Q ),
    .c(RESET),
    .y(_03340_)
  );
  al_aoi21ftf _08964_ (
    .a(\DFF_1100.Q ),
    .b(\DFF_1138.Q ),
    .c(_03340_),
    .y(\DFF_1139.D )
  );
  al_oa21ftt _08965_ (
    .a(\DFF_1099.Q ),
    .b(\DFF_1139.Q ),
    .c(RESET),
    .y(_03341_)
  );
  al_aoi21ftf _08966_ (
    .a(\DFF_1099.Q ),
    .b(\DFF_1139.Q ),
    .c(_03341_),
    .y(\DFF_1140.D )
  );
  al_oa21ftt _08967_ (
    .a(\DFF_1098.Q ),
    .b(\DFF_1140.Q ),
    .c(RESET),
    .y(_03342_)
  );
  al_aoi21ftf _08968_ (
    .a(\DFF_1098.Q ),
    .b(\DFF_1140.Q ),
    .c(_03342_),
    .y(\DFF_1141.D )
  );
  al_oa21ftt _08969_ (
    .a(\DFF_1097.Q ),
    .b(\DFF_1141.Q ),
    .c(RESET),
    .y(_03343_)
  );
  al_aoi21ftf _08970_ (
    .a(\DFF_1097.Q ),
    .b(\DFF_1141.Q ),
    .c(_03343_),
    .y(\DFF_1142.D )
  );
  al_oa21ftt _08971_ (
    .a(\DFF_1096.Q ),
    .b(\DFF_1142.Q ),
    .c(RESET),
    .y(_03344_)
  );
  al_aoi21ftf _08972_ (
    .a(\DFF_1096.Q ),
    .b(\DFF_1142.Q ),
    .c(_03344_),
    .y(\DFF_1143.D )
  );
  al_oa21ftt _08973_ (
    .a(\DFF_1095.Q ),
    .b(\DFF_1143.Q ),
    .c(RESET),
    .y(_03345_)
  );
  al_aoi21ftf _08974_ (
    .a(\DFF_1095.Q ),
    .b(\DFF_1143.Q ),
    .c(_03345_),
    .y(\DFF_1144.D )
  );
  al_oa21ftt _08975_ (
    .a(\DFF_1094.Q ),
    .b(\DFF_1144.Q ),
    .c(RESET),
    .y(_03346_)
  );
  al_aoi21ftf _08976_ (
    .a(\DFF_1094.Q ),
    .b(\DFF_1144.Q ),
    .c(_03346_),
    .y(\DFF_1145.D )
  );
  al_oa21ftt _08977_ (
    .a(\DFF_1093.Q ),
    .b(\DFF_1145.Q ),
    .c(RESET),
    .y(_03347_)
  );
  al_aoi21ftf _08978_ (
    .a(\DFF_1093.Q ),
    .b(\DFF_1145.Q ),
    .c(_03347_),
    .y(\DFF_1146.D )
  );
  al_oa21ftt _08979_ (
    .a(\DFF_1092.Q ),
    .b(\DFF_1146.Q ),
    .c(RESET),
    .y(_03348_)
  );
  al_aoi21ftf _08980_ (
    .a(\DFF_1092.Q ),
    .b(\DFF_1146.Q ),
    .c(_03348_),
    .y(\DFF_1147.D )
  );
  al_oa21ftt _08981_ (
    .a(\DFF_1091.Q ),
    .b(\DFF_1147.Q ),
    .c(RESET),
    .y(_03349_)
  );
  al_aoi21ftf _08982_ (
    .a(\DFF_1091.Q ),
    .b(\DFF_1147.Q ),
    .c(_03349_),
    .y(\DFF_1148.D )
  );
  al_oa21ftt _08983_ (
    .a(\DFF_1090.Q ),
    .b(\DFF_1148.Q ),
    .c(RESET),
    .y(_03350_)
  );
  al_aoi21ftf _08984_ (
    .a(\DFF_1090.Q ),
    .b(\DFF_1148.Q ),
    .c(_03350_),
    .y(\DFF_1149.D )
  );
  al_oa21ftt _08985_ (
    .a(\DFF_1089.Q ),
    .b(\DFF_1149.Q ),
    .c(RESET),
    .y(_03351_)
  );
  al_aoi21ftf _08986_ (
    .a(\DFF_1089.Q ),
    .b(\DFF_1149.Q ),
    .c(_03351_),
    .y(\DFF_1150.D )
  );
  al_oa21ftt _08987_ (
    .a(\DFF_1088.Q ),
    .b(\DFF_1150.Q ),
    .c(RESET),
    .y(_03352_)
  );
  al_aoi21ftf _08988_ (
    .a(\DFF_1088.Q ),
    .b(\DFF_1150.Q ),
    .c(_03352_),
    .y(\DFF_1151.D )
  );
  al_and2 _08989_ (
    .a(RESET),
    .b(\DFF_1153.Q ),
    .y(\DFF_1152.D )
  );
  al_and2 _08990_ (
    .a(RESET),
    .b(\DFF_1154.Q ),
    .y(\DFF_1153.D )
  );
  al_and2 _08991_ (
    .a(RESET),
    .b(\DFF_1155.Q ),
    .y(\DFF_1154.D )
  );
  al_and2 _08992_ (
    .a(RESET),
    .b(\DFF_1156.Q ),
    .y(\DFF_1155.D )
  );
  al_and2 _08993_ (
    .a(RESET),
    .b(\DFF_1157.Q ),
    .y(\DFF_1156.D )
  );
  al_and2 _08994_ (
    .a(RESET),
    .b(\DFF_1158.Q ),
    .y(\DFF_1157.D )
  );
  al_and2 _08995_ (
    .a(RESET),
    .b(\DFF_1159.Q ),
    .y(\DFF_1158.D )
  );
  al_and2 _08996_ (
    .a(RESET),
    .b(\DFF_1160.Q ),
    .y(\DFF_1159.D )
  );
  al_and2 _08997_ (
    .a(RESET),
    .b(\DFF_1161.Q ),
    .y(\DFF_1160.D )
  );
  al_and2 _08998_ (
    .a(RESET),
    .b(\DFF_1162.Q ),
    .y(\DFF_1161.D )
  );
  al_and2 _08999_ (
    .a(RESET),
    .b(\DFF_1163.Q ),
    .y(\DFF_1162.D )
  );
  al_and2 _09000_ (
    .a(RESET),
    .b(\DFF_1164.Q ),
    .y(\DFF_1163.D )
  );
  al_and2 _09001_ (
    .a(RESET),
    .b(\DFF_1165.Q ),
    .y(\DFF_1164.D )
  );
  al_and2 _09002_ (
    .a(RESET),
    .b(\DFF_1166.Q ),
    .y(\DFF_1165.D )
  );
  al_and2 _09003_ (
    .a(RESET),
    .b(\DFF_1167.Q ),
    .y(\DFF_1166.D )
  );
  al_and2 _09004_ (
    .a(RESET),
    .b(\DFF_1168.Q ),
    .y(\DFF_1167.D )
  );
  al_and2 _09005_ (
    .a(RESET),
    .b(\DFF_1169.Q ),
    .y(\DFF_1168.D )
  );
  al_and2 _09006_ (
    .a(RESET),
    .b(\DFF_1170.Q ),
    .y(\DFF_1169.D )
  );
  al_and2 _09007_ (
    .a(RESET),
    .b(\DFF_1171.Q ),
    .y(\DFF_1170.D )
  );
  al_and2 _09008_ (
    .a(RESET),
    .b(\DFF_1172.Q ),
    .y(\DFF_1171.D )
  );
  al_and2 _09009_ (
    .a(RESET),
    .b(\DFF_1173.Q ),
    .y(\DFF_1172.D )
  );
  al_and2 _09010_ (
    .a(RESET),
    .b(\DFF_1174.Q ),
    .y(\DFF_1173.D )
  );
  al_and2 _09011_ (
    .a(RESET),
    .b(\DFF_1175.Q ),
    .y(\DFF_1174.D )
  );
  al_and2 _09012_ (
    .a(RESET),
    .b(\DFF_1176.Q ),
    .y(\DFF_1175.D )
  );
  al_and2 _09013_ (
    .a(RESET),
    .b(\DFF_1177.Q ),
    .y(\DFF_1176.D )
  );
  al_and2 _09014_ (
    .a(RESET),
    .b(\DFF_1178.Q ),
    .y(\DFF_1177.D )
  );
  al_and2 _09015_ (
    .a(RESET),
    .b(\DFF_1179.Q ),
    .y(\DFF_1178.D )
  );
  al_and2 _09016_ (
    .a(RESET),
    .b(\DFF_1180.Q ),
    .y(\DFF_1179.D )
  );
  al_and2 _09017_ (
    .a(RESET),
    .b(\DFF_1181.Q ),
    .y(\DFF_1180.D )
  );
  al_and2 _09018_ (
    .a(RESET),
    .b(\DFF_1182.Q ),
    .y(\DFF_1181.D )
  );
  al_and2 _09019_ (
    .a(RESET),
    .b(\DFF_1183.Q ),
    .y(\DFF_1182.D )
  );
  al_and2ft _09020_ (
    .a(\DFF_1152.Q ),
    .b(RESET),
    .y(\DFF_1183.D )
  );
  al_or2 _09021_ (
    .a(TM1),
    .b(\DFF_1440.Q ),
    .y(_03353_)
  );
  al_nand2 _09022_ (
    .a(TM1),
    .b(\DFF_1440.Q ),
    .y(_03354_)
  );
  al_nand3 _09023_ (
    .a(\DFF_1472.Q ),
    .b(_03353_),
    .c(_03354_),
    .y(_03355_)
  );
  al_nand2ft _09024_ (
    .a(TM1),
    .b(\DFF_1440.Q ),
    .y(_03356_)
  );
  al_and2ft _09025_ (
    .a(\DFF_1440.Q ),
    .b(TM1),
    .y(_03357_)
  );
  al_and3fft _09026_ (
    .a(\DFF_1472.Q ),
    .b(_03357_),
    .c(_03356_),
    .y(_03358_)
  );
  al_and2ft _09027_ (
    .a(\DFF_1408.Q ),
    .b(\DFF_1376.Q ),
    .y(_03359_)
  );
  al_nand2ft _09028_ (
    .a(\DFF_1376.Q ),
    .b(\DFF_1408.Q ),
    .y(_03360_)
  );
  al_nand2ft _09029_ (
    .a(_03359_),
    .b(_03360_),
    .y(_03361_)
  );
  al_oai21ftf _09030_ (
    .a(_03355_),
    .b(_03358_),
    .c(_03361_),
    .y(_03362_)
  );
  al_nand3ftt _09031_ (
    .a(_03358_),
    .b(_03355_),
    .c(_03361_),
    .y(_03363_)
  );
  al_nand3 _09032_ (
    .a(_00448_),
    .b(_03362_),
    .c(_03363_),
    .y(_03364_)
  );
  al_aoi21 _09033_ (
    .a(TM0),
    .b(\DFF_1343.Q ),
    .c(TM1),
    .y(_03365_)
  );
  al_nand2 _09034_ (
    .a(_03365_),
    .b(_03364_),
    .y(_03366_)
  );
  al_aoi21ttf _09035_ (
    .a(\DFF_1152.Q ),
    .b(TM0),
    .c(TM1),
    .y(_03367_)
  );
  al_and2 _09036_ (
    .a(_03367_),
    .b(_02875_),
    .y(_03368_)
  );
  al_nor3fft _09037_ (
    .a(RESET),
    .b(_03366_),
    .c(_03368_),
    .y(\DFF_1184.D )
  );
  al_or2 _09038_ (
    .a(TM1),
    .b(\DFF_1441.Q ),
    .y(_03369_)
  );
  al_nand2 _09039_ (
    .a(TM1),
    .b(\DFF_1441.Q ),
    .y(_03370_)
  );
  al_nand3 _09040_ (
    .a(\DFF_1473.Q ),
    .b(_03369_),
    .c(_03370_),
    .y(_03371_)
  );
  al_nand2ft _09041_ (
    .a(TM1),
    .b(\DFF_1441.Q ),
    .y(_03372_)
  );
  al_and2ft _09042_ (
    .a(\DFF_1441.Q ),
    .b(TM1),
    .y(_03373_)
  );
  al_and3fft _09043_ (
    .a(\DFF_1473.Q ),
    .b(_03373_),
    .c(_03372_),
    .y(_03374_)
  );
  al_and2ft _09044_ (
    .a(\DFF_1409.Q ),
    .b(\DFF_1377.Q ),
    .y(_03375_)
  );
  al_nand2ft _09045_ (
    .a(\DFF_1377.Q ),
    .b(\DFF_1409.Q ),
    .y(_03376_)
  );
  al_nand2ft _09046_ (
    .a(_03375_),
    .b(_03376_),
    .y(_03377_)
  );
  al_oai21ftf _09047_ (
    .a(_03371_),
    .b(_03374_),
    .c(_03377_),
    .y(_03378_)
  );
  al_nand3ftt _09048_ (
    .a(_03374_),
    .b(_03371_),
    .c(_03377_),
    .y(_03379_)
  );
  al_nand3 _09049_ (
    .a(_00448_),
    .b(_03378_),
    .c(_03379_),
    .y(_03380_)
  );
  al_aoi21 _09050_ (
    .a(TM0),
    .b(\DFF_1342.Q ),
    .c(TM1),
    .y(_03381_)
  );
  al_nand2 _09051_ (
    .a(_03381_),
    .b(_03380_),
    .y(_03382_)
  );
  al_aoi21ttf _09052_ (
    .a(TM0),
    .b(\DFF_1153.Q ),
    .c(TM1),
    .y(_03383_)
  );
  al_and2 _09053_ (
    .a(_03383_),
    .b(_02891_),
    .y(_03384_)
  );
  al_nor3fft _09054_ (
    .a(RESET),
    .b(_03382_),
    .c(_03384_),
    .y(\DFF_1185.D )
  );
  al_or2 _09055_ (
    .a(TM1),
    .b(\DFF_1442.Q ),
    .y(_03385_)
  );
  al_nand2 _09056_ (
    .a(TM1),
    .b(\DFF_1442.Q ),
    .y(_03386_)
  );
  al_nand3 _09057_ (
    .a(\DFF_1474.Q ),
    .b(_03385_),
    .c(_03386_),
    .y(_03387_)
  );
  al_nand2ft _09058_ (
    .a(TM1),
    .b(\DFF_1442.Q ),
    .y(_03388_)
  );
  al_and2ft _09059_ (
    .a(\DFF_1442.Q ),
    .b(TM1),
    .y(_03389_)
  );
  al_and3fft _09060_ (
    .a(\DFF_1474.Q ),
    .b(_03389_),
    .c(_03388_),
    .y(_03390_)
  );
  al_and2ft _09061_ (
    .a(\DFF_1410.Q ),
    .b(\DFF_1378.Q ),
    .y(_03391_)
  );
  al_nand2ft _09062_ (
    .a(\DFF_1378.Q ),
    .b(\DFF_1410.Q ),
    .y(_03392_)
  );
  al_nand2ft _09063_ (
    .a(_03391_),
    .b(_03392_),
    .y(_03393_)
  );
  al_oai21ftf _09064_ (
    .a(_03387_),
    .b(_03390_),
    .c(_03393_),
    .y(_03394_)
  );
  al_nand3ftt _09065_ (
    .a(_03390_),
    .b(_03387_),
    .c(_03393_),
    .y(_03395_)
  );
  al_nand3 _09066_ (
    .a(_00448_),
    .b(_03394_),
    .c(_03395_),
    .y(_03396_)
  );
  al_aoi21 _09067_ (
    .a(TM0),
    .b(\DFF_1341.Q ),
    .c(TM1),
    .y(_03397_)
  );
  al_nand2 _09068_ (
    .a(_03397_),
    .b(_03396_),
    .y(_03398_)
  );
  al_aoi21ttf _09069_ (
    .a(TM0),
    .b(\DFF_1154.Q ),
    .c(TM1),
    .y(_03399_)
  );
  al_and2 _09070_ (
    .a(_03399_),
    .b(_02907_),
    .y(_03400_)
  );
  al_nor3fft _09071_ (
    .a(RESET),
    .b(_03398_),
    .c(_03400_),
    .y(\DFF_1186.D )
  );
  al_or2 _09072_ (
    .a(TM1),
    .b(\DFF_1443.Q ),
    .y(_03401_)
  );
  al_nand2 _09073_ (
    .a(TM1),
    .b(\DFF_1443.Q ),
    .y(_03402_)
  );
  al_nand3 _09074_ (
    .a(\DFF_1475.Q ),
    .b(_03401_),
    .c(_03402_),
    .y(_03403_)
  );
  al_nand2ft _09075_ (
    .a(TM1),
    .b(\DFF_1443.Q ),
    .y(_03404_)
  );
  al_and2ft _09076_ (
    .a(\DFF_1443.Q ),
    .b(TM1),
    .y(_03405_)
  );
  al_and3fft _09077_ (
    .a(\DFF_1475.Q ),
    .b(_03405_),
    .c(_03404_),
    .y(_03406_)
  );
  al_and2ft _09078_ (
    .a(\DFF_1411.Q ),
    .b(\DFF_1379.Q ),
    .y(_03407_)
  );
  al_nand2ft _09079_ (
    .a(\DFF_1379.Q ),
    .b(\DFF_1411.Q ),
    .y(_03408_)
  );
  al_nand2ft _09080_ (
    .a(_03407_),
    .b(_03408_),
    .y(_03409_)
  );
  al_oai21ftf _09081_ (
    .a(_03403_),
    .b(_03406_),
    .c(_03409_),
    .y(_03410_)
  );
  al_nand3ftt _09082_ (
    .a(_03406_),
    .b(_03403_),
    .c(_03409_),
    .y(_03411_)
  );
  al_nand3 _09083_ (
    .a(_00448_),
    .b(_03410_),
    .c(_03411_),
    .y(_03412_)
  );
  al_aoi21 _09084_ (
    .a(TM0),
    .b(\DFF_1340.Q ),
    .c(TM1),
    .y(_03413_)
  );
  al_nand2 _09085_ (
    .a(_03413_),
    .b(_03412_),
    .y(_03414_)
  );
  al_aoi21ttf _09086_ (
    .a(TM0),
    .b(\DFF_1155.Q ),
    .c(TM1),
    .y(_03415_)
  );
  al_and2 _09087_ (
    .a(_03415_),
    .b(_02923_),
    .y(_03416_)
  );
  al_nor3fft _09088_ (
    .a(RESET),
    .b(_03414_),
    .c(_03416_),
    .y(\DFF_1187.D )
  );
  al_or2 _09089_ (
    .a(TM1),
    .b(\DFF_1444.Q ),
    .y(_03417_)
  );
  al_nand2 _09090_ (
    .a(TM1),
    .b(\DFF_1444.Q ),
    .y(_03418_)
  );
  al_nand3 _09091_ (
    .a(\DFF_1476.Q ),
    .b(_03417_),
    .c(_03418_),
    .y(_03419_)
  );
  al_nand2ft _09092_ (
    .a(TM1),
    .b(\DFF_1444.Q ),
    .y(_03420_)
  );
  al_and2ft _09093_ (
    .a(\DFF_1444.Q ),
    .b(TM1),
    .y(_03421_)
  );
  al_and3fft _09094_ (
    .a(\DFF_1476.Q ),
    .b(_03421_),
    .c(_03420_),
    .y(_03422_)
  );
  al_and2ft _09095_ (
    .a(\DFF_1412.Q ),
    .b(\DFF_1380.Q ),
    .y(_03423_)
  );
  al_nand2ft _09096_ (
    .a(\DFF_1380.Q ),
    .b(\DFF_1412.Q ),
    .y(_03424_)
  );
  al_nand2ft _09097_ (
    .a(_03423_),
    .b(_03424_),
    .y(_03425_)
  );
  al_oai21ftf _09098_ (
    .a(_03419_),
    .b(_03422_),
    .c(_03425_),
    .y(_03426_)
  );
  al_nand3ftt _09099_ (
    .a(_03422_),
    .b(_03419_),
    .c(_03425_),
    .y(_03427_)
  );
  al_nand3 _09100_ (
    .a(_00448_),
    .b(_03426_),
    .c(_03427_),
    .y(_03428_)
  );
  al_aoi21 _09101_ (
    .a(TM0),
    .b(\DFF_1339.Q ),
    .c(TM1),
    .y(_03429_)
  );
  al_nand2 _09102_ (
    .a(_03429_),
    .b(_03428_),
    .y(_03430_)
  );
  al_aoi21ttf _09103_ (
    .a(TM0),
    .b(\DFF_1156.Q ),
    .c(TM1),
    .y(_03431_)
  );
  al_and2 _09104_ (
    .a(_03431_),
    .b(_02939_),
    .y(_03432_)
  );
  al_nor3fft _09105_ (
    .a(RESET),
    .b(_03430_),
    .c(_03432_),
    .y(\DFF_1188.D )
  );
  al_or2 _09106_ (
    .a(TM1),
    .b(\DFF_1445.Q ),
    .y(_03433_)
  );
  al_nand2 _09107_ (
    .a(TM1),
    .b(\DFF_1445.Q ),
    .y(_03434_)
  );
  al_nand3 _09108_ (
    .a(\DFF_1477.Q ),
    .b(_03433_),
    .c(_03434_),
    .y(_03435_)
  );
  al_nand2ft _09109_ (
    .a(TM1),
    .b(\DFF_1445.Q ),
    .y(_03436_)
  );
  al_and2ft _09110_ (
    .a(\DFF_1445.Q ),
    .b(TM1),
    .y(_03437_)
  );
  al_and3fft _09111_ (
    .a(\DFF_1477.Q ),
    .b(_03437_),
    .c(_03436_),
    .y(_03438_)
  );
  al_and2ft _09112_ (
    .a(\DFF_1413.Q ),
    .b(\DFF_1381.Q ),
    .y(_03439_)
  );
  al_nand2ft _09113_ (
    .a(\DFF_1381.Q ),
    .b(\DFF_1413.Q ),
    .y(_03440_)
  );
  al_nand2ft _09114_ (
    .a(_03439_),
    .b(_03440_),
    .y(_03441_)
  );
  al_oai21ftf _09115_ (
    .a(_03435_),
    .b(_03438_),
    .c(_03441_),
    .y(_03442_)
  );
  al_nand3ftt _09116_ (
    .a(_03438_),
    .b(_03435_),
    .c(_03441_),
    .y(_03443_)
  );
  al_nand3 _09117_ (
    .a(_00448_),
    .b(_03442_),
    .c(_03443_),
    .y(_03444_)
  );
  al_aoi21 _09118_ (
    .a(TM0),
    .b(\DFF_1338.Q ),
    .c(TM1),
    .y(_03445_)
  );
  al_nand2 _09119_ (
    .a(_03445_),
    .b(_03444_),
    .y(_03446_)
  );
  al_aoi21ttf _09120_ (
    .a(TM0),
    .b(\DFF_1157.Q ),
    .c(TM1),
    .y(_03447_)
  );
  al_and2 _09121_ (
    .a(_03447_),
    .b(_02955_),
    .y(_03448_)
  );
  al_nor3fft _09122_ (
    .a(RESET),
    .b(_03446_),
    .c(_03448_),
    .y(\DFF_1189.D )
  );
  al_or2 _09123_ (
    .a(TM1),
    .b(\DFF_1446.Q ),
    .y(_03449_)
  );
  al_nand2 _09124_ (
    .a(TM1),
    .b(\DFF_1446.Q ),
    .y(_03450_)
  );
  al_nand3 _09125_ (
    .a(\DFF_1478.Q ),
    .b(_03449_),
    .c(_03450_),
    .y(_03451_)
  );
  al_nand2ft _09126_ (
    .a(TM1),
    .b(\DFF_1446.Q ),
    .y(_03452_)
  );
  al_and2ft _09127_ (
    .a(\DFF_1446.Q ),
    .b(TM1),
    .y(_03453_)
  );
  al_and3fft _09128_ (
    .a(\DFF_1478.Q ),
    .b(_03453_),
    .c(_03452_),
    .y(_03454_)
  );
  al_and2ft _09129_ (
    .a(\DFF_1414.Q ),
    .b(\DFF_1382.Q ),
    .y(_03455_)
  );
  al_nand2ft _09130_ (
    .a(\DFF_1382.Q ),
    .b(\DFF_1414.Q ),
    .y(_03456_)
  );
  al_nand2ft _09131_ (
    .a(_03455_),
    .b(_03456_),
    .y(_03457_)
  );
  al_oai21ftf _09132_ (
    .a(_03451_),
    .b(_03454_),
    .c(_03457_),
    .y(_03458_)
  );
  al_nand3ftt _09133_ (
    .a(_03454_),
    .b(_03451_),
    .c(_03457_),
    .y(_03459_)
  );
  al_nand3 _09134_ (
    .a(_00448_),
    .b(_03458_),
    .c(_03459_),
    .y(_03460_)
  );
  al_aoi21 _09135_ (
    .a(TM0),
    .b(\DFF_1337.Q ),
    .c(TM1),
    .y(_03461_)
  );
  al_nand2 _09136_ (
    .a(_03461_),
    .b(_03460_),
    .y(_03462_)
  );
  al_aoi21ttf _09137_ (
    .a(TM0),
    .b(\DFF_1158.Q ),
    .c(TM1),
    .y(_03463_)
  );
  al_and2 _09138_ (
    .a(_03463_),
    .b(_02971_),
    .y(_03464_)
  );
  al_nor3fft _09139_ (
    .a(RESET),
    .b(_03462_),
    .c(_03464_),
    .y(\DFF_1190.D )
  );
  al_or2 _09140_ (
    .a(TM1),
    .b(\DFF_1447.Q ),
    .y(_03465_)
  );
  al_nand2 _09141_ (
    .a(TM1),
    .b(\DFF_1447.Q ),
    .y(_03466_)
  );
  al_nand3 _09142_ (
    .a(\DFF_1479.Q ),
    .b(_03465_),
    .c(_03466_),
    .y(_03467_)
  );
  al_nand2ft _09143_ (
    .a(TM1),
    .b(\DFF_1447.Q ),
    .y(_03468_)
  );
  al_and2ft _09144_ (
    .a(\DFF_1447.Q ),
    .b(TM1),
    .y(_03469_)
  );
  al_and3fft _09145_ (
    .a(\DFF_1479.Q ),
    .b(_03469_),
    .c(_03468_),
    .y(_03470_)
  );
  al_and2ft _09146_ (
    .a(\DFF_1415.Q ),
    .b(\DFF_1383.Q ),
    .y(_03471_)
  );
  al_nand2ft _09147_ (
    .a(\DFF_1383.Q ),
    .b(\DFF_1415.Q ),
    .y(_03472_)
  );
  al_nand2ft _09148_ (
    .a(_03471_),
    .b(_03472_),
    .y(_03473_)
  );
  al_oai21ftf _09149_ (
    .a(_03467_),
    .b(_03470_),
    .c(_03473_),
    .y(_03474_)
  );
  al_nand3ftt _09150_ (
    .a(_03470_),
    .b(_03467_),
    .c(_03473_),
    .y(_03475_)
  );
  al_nand3 _09151_ (
    .a(_00448_),
    .b(_03474_),
    .c(_03475_),
    .y(_03476_)
  );
  al_aoi21 _09152_ (
    .a(TM0),
    .b(\DFF_1336.Q ),
    .c(TM1),
    .y(_03477_)
  );
  al_nand2 _09153_ (
    .a(_03477_),
    .b(_03476_),
    .y(_03478_)
  );
  al_aoi21ttf _09154_ (
    .a(TM0),
    .b(\DFF_1159.Q ),
    .c(TM1),
    .y(_03479_)
  );
  al_and2 _09155_ (
    .a(_03479_),
    .b(_02987_),
    .y(_03480_)
  );
  al_nor3fft _09156_ (
    .a(RESET),
    .b(_03478_),
    .c(_03480_),
    .y(\DFF_1191.D )
  );
  al_or2 _09157_ (
    .a(TM1),
    .b(\DFF_1448.Q ),
    .y(_03481_)
  );
  al_nand2 _09158_ (
    .a(TM1),
    .b(\DFF_1448.Q ),
    .y(_03482_)
  );
  al_nand3 _09159_ (
    .a(\DFF_1480.Q ),
    .b(_03481_),
    .c(_03482_),
    .y(_03483_)
  );
  al_nand2ft _09160_ (
    .a(TM1),
    .b(\DFF_1448.Q ),
    .y(_03484_)
  );
  al_and2ft _09161_ (
    .a(\DFF_1448.Q ),
    .b(TM1),
    .y(_03485_)
  );
  al_and3fft _09162_ (
    .a(\DFF_1480.Q ),
    .b(_03485_),
    .c(_03484_),
    .y(_03486_)
  );
  al_and2ft _09163_ (
    .a(\DFF_1416.Q ),
    .b(\DFF_1384.Q ),
    .y(_03487_)
  );
  al_nand2ft _09164_ (
    .a(\DFF_1384.Q ),
    .b(\DFF_1416.Q ),
    .y(_03488_)
  );
  al_nand2ft _09165_ (
    .a(_03487_),
    .b(_03488_),
    .y(_03489_)
  );
  al_oai21ftf _09166_ (
    .a(_03483_),
    .b(_03486_),
    .c(_03489_),
    .y(_03490_)
  );
  al_nand3ftt _09167_ (
    .a(_03486_),
    .b(_03483_),
    .c(_03489_),
    .y(_03491_)
  );
  al_nand3 _09168_ (
    .a(_00448_),
    .b(_03490_),
    .c(_03491_),
    .y(_03492_)
  );
  al_aoi21 _09169_ (
    .a(TM0),
    .b(\DFF_1335.Q ),
    .c(TM1),
    .y(_03493_)
  );
  al_nand2 _09170_ (
    .a(_03493_),
    .b(_03492_),
    .y(_03494_)
  );
  al_aoi21ttf _09171_ (
    .a(TM0),
    .b(\DFF_1160.Q ),
    .c(TM1),
    .y(_03495_)
  );
  al_and2 _09172_ (
    .a(_03495_),
    .b(_03003_),
    .y(_03496_)
  );
  al_nor3fft _09173_ (
    .a(RESET),
    .b(_03494_),
    .c(_03496_),
    .y(\DFF_1192.D )
  );
  al_or2 _09174_ (
    .a(TM1),
    .b(\DFF_1449.Q ),
    .y(_03497_)
  );
  al_nand2 _09175_ (
    .a(TM1),
    .b(\DFF_1449.Q ),
    .y(_03498_)
  );
  al_nand3 _09176_ (
    .a(\DFF_1481.Q ),
    .b(_03497_),
    .c(_03498_),
    .y(_03499_)
  );
  al_nand2ft _09177_ (
    .a(TM1),
    .b(\DFF_1449.Q ),
    .y(_03500_)
  );
  al_and2ft _09178_ (
    .a(\DFF_1449.Q ),
    .b(TM1),
    .y(_03501_)
  );
  al_and3fft _09179_ (
    .a(\DFF_1481.Q ),
    .b(_03501_),
    .c(_03500_),
    .y(_03502_)
  );
  al_and2ft _09180_ (
    .a(\DFF_1417.Q ),
    .b(\DFF_1385.Q ),
    .y(_03503_)
  );
  al_nand2ft _09181_ (
    .a(\DFF_1385.Q ),
    .b(\DFF_1417.Q ),
    .y(_03504_)
  );
  al_nand2ft _09182_ (
    .a(_03503_),
    .b(_03504_),
    .y(_03505_)
  );
  al_oai21ftf _09183_ (
    .a(_03499_),
    .b(_03502_),
    .c(_03505_),
    .y(_03506_)
  );
  al_nand3ftt _09184_ (
    .a(_03502_),
    .b(_03499_),
    .c(_03505_),
    .y(_03507_)
  );
  al_nand3 _09185_ (
    .a(_00448_),
    .b(_03506_),
    .c(_03507_),
    .y(_03508_)
  );
  al_aoi21 _09186_ (
    .a(TM0),
    .b(\DFF_1334.Q ),
    .c(TM1),
    .y(_03509_)
  );
  al_nand2 _09187_ (
    .a(_03509_),
    .b(_03508_),
    .y(_03510_)
  );
  al_aoi21ttf _09188_ (
    .a(TM0),
    .b(\DFF_1161.Q ),
    .c(TM1),
    .y(_03511_)
  );
  al_and2 _09189_ (
    .a(_03511_),
    .b(_03019_),
    .y(_03512_)
  );
  al_nor3fft _09190_ (
    .a(RESET),
    .b(_03510_),
    .c(_03512_),
    .y(\DFF_1193.D )
  );
  al_or2 _09191_ (
    .a(TM1),
    .b(\DFF_1450.Q ),
    .y(_03513_)
  );
  al_nand2 _09192_ (
    .a(TM1),
    .b(\DFF_1450.Q ),
    .y(_03514_)
  );
  al_nand3 _09193_ (
    .a(\DFF_1482.Q ),
    .b(_03513_),
    .c(_03514_),
    .y(_03515_)
  );
  al_nand2ft _09194_ (
    .a(TM1),
    .b(\DFF_1450.Q ),
    .y(_03516_)
  );
  al_and2ft _09195_ (
    .a(\DFF_1450.Q ),
    .b(TM1),
    .y(_03517_)
  );
  al_and3fft _09196_ (
    .a(\DFF_1482.Q ),
    .b(_03517_),
    .c(_03516_),
    .y(_03518_)
  );
  al_and2ft _09197_ (
    .a(\DFF_1418.Q ),
    .b(\DFF_1386.Q ),
    .y(_03519_)
  );
  al_nand2ft _09198_ (
    .a(\DFF_1386.Q ),
    .b(\DFF_1418.Q ),
    .y(_03520_)
  );
  al_nand2ft _09199_ (
    .a(_03519_),
    .b(_03520_),
    .y(_03521_)
  );
  al_oai21ftf _09200_ (
    .a(_03515_),
    .b(_03518_),
    .c(_03521_),
    .y(_03522_)
  );
  al_nand3ftt _09201_ (
    .a(_03518_),
    .b(_03515_),
    .c(_03521_),
    .y(_03523_)
  );
  al_nand3 _09202_ (
    .a(_00448_),
    .b(_03522_),
    .c(_03523_),
    .y(_03524_)
  );
  al_aoi21 _09203_ (
    .a(TM0),
    .b(\DFF_1333.Q ),
    .c(TM1),
    .y(_03525_)
  );
  al_nand2 _09204_ (
    .a(_03525_),
    .b(_03524_),
    .y(_03526_)
  );
  al_aoi21ttf _09205_ (
    .a(TM0),
    .b(\DFF_1162.Q ),
    .c(TM1),
    .y(_03527_)
  );
  al_and2 _09206_ (
    .a(_03527_),
    .b(_03035_),
    .y(_03528_)
  );
  al_nor3fft _09207_ (
    .a(RESET),
    .b(_03526_),
    .c(_03528_),
    .y(\DFF_1194.D )
  );
  al_or2 _09208_ (
    .a(TM1),
    .b(\DFF_1451.Q ),
    .y(_03529_)
  );
  al_nand2 _09209_ (
    .a(TM1),
    .b(\DFF_1451.Q ),
    .y(_03530_)
  );
  al_nand3 _09210_ (
    .a(\DFF_1483.Q ),
    .b(_03529_),
    .c(_03530_),
    .y(_03531_)
  );
  al_nand2ft _09211_ (
    .a(TM1),
    .b(\DFF_1451.Q ),
    .y(_03532_)
  );
  al_and2ft _09212_ (
    .a(\DFF_1451.Q ),
    .b(TM1),
    .y(_03533_)
  );
  al_and3fft _09213_ (
    .a(\DFF_1483.Q ),
    .b(_03533_),
    .c(_03532_),
    .y(_03534_)
  );
  al_and2ft _09214_ (
    .a(\DFF_1419.Q ),
    .b(\DFF_1387.Q ),
    .y(_03535_)
  );
  al_nand2ft _09215_ (
    .a(\DFF_1387.Q ),
    .b(\DFF_1419.Q ),
    .y(_03536_)
  );
  al_nand2ft _09216_ (
    .a(_03535_),
    .b(_03536_),
    .y(_03537_)
  );
  al_oai21ftf _09217_ (
    .a(_03531_),
    .b(_03534_),
    .c(_03537_),
    .y(_03538_)
  );
  al_nand3ftt _09218_ (
    .a(_03534_),
    .b(_03531_),
    .c(_03537_),
    .y(_03539_)
  );
  al_nand3 _09219_ (
    .a(_00448_),
    .b(_03538_),
    .c(_03539_),
    .y(_03540_)
  );
  al_aoi21 _09220_ (
    .a(TM0),
    .b(\DFF_1332.Q ),
    .c(TM1),
    .y(_03541_)
  );
  al_nand2 _09221_ (
    .a(_03541_),
    .b(_03540_),
    .y(_03542_)
  );
  al_aoi21ttf _09222_ (
    .a(TM0),
    .b(\DFF_1163.Q ),
    .c(TM1),
    .y(_03543_)
  );
  al_and2 _09223_ (
    .a(_03543_),
    .b(_03051_),
    .y(_03544_)
  );
  al_nor3fft _09224_ (
    .a(RESET),
    .b(_03542_),
    .c(_03544_),
    .y(\DFF_1195.D )
  );
  al_or2 _09225_ (
    .a(TM1),
    .b(\DFF_1452.Q ),
    .y(_03545_)
  );
  al_nand2 _09226_ (
    .a(TM1),
    .b(\DFF_1452.Q ),
    .y(_03546_)
  );
  al_nand3 _09227_ (
    .a(\DFF_1484.Q ),
    .b(_03545_),
    .c(_03546_),
    .y(_03547_)
  );
  al_nand2ft _09228_ (
    .a(TM1),
    .b(\DFF_1452.Q ),
    .y(_03548_)
  );
  al_and2ft _09229_ (
    .a(\DFF_1452.Q ),
    .b(TM1),
    .y(_03549_)
  );
  al_and3fft _09230_ (
    .a(\DFF_1484.Q ),
    .b(_03549_),
    .c(_03548_),
    .y(_03550_)
  );
  al_and2ft _09231_ (
    .a(\DFF_1420.Q ),
    .b(\DFF_1388.Q ),
    .y(_03551_)
  );
  al_nand2ft _09232_ (
    .a(\DFF_1388.Q ),
    .b(\DFF_1420.Q ),
    .y(_03552_)
  );
  al_nand2ft _09233_ (
    .a(_03551_),
    .b(_03552_),
    .y(_03553_)
  );
  al_oai21ftf _09234_ (
    .a(_03547_),
    .b(_03550_),
    .c(_03553_),
    .y(_03554_)
  );
  al_nand3ftt _09235_ (
    .a(_03550_),
    .b(_03547_),
    .c(_03553_),
    .y(_03555_)
  );
  al_nand3 _09236_ (
    .a(_00448_),
    .b(_03554_),
    .c(_03555_),
    .y(_03556_)
  );
  al_aoi21 _09237_ (
    .a(TM0),
    .b(\DFF_1331.Q ),
    .c(TM1),
    .y(_03557_)
  );
  al_nand2 _09238_ (
    .a(_03557_),
    .b(_03556_),
    .y(_03558_)
  );
  al_aoi21ttf _09239_ (
    .a(TM0),
    .b(\DFF_1164.Q ),
    .c(TM1),
    .y(_03559_)
  );
  al_and2 _09240_ (
    .a(_03559_),
    .b(_03067_),
    .y(_03560_)
  );
  al_nor3fft _09241_ (
    .a(RESET),
    .b(_03558_),
    .c(_03560_),
    .y(\DFF_1196.D )
  );
  al_or2 _09242_ (
    .a(TM1),
    .b(\DFF_1453.Q ),
    .y(_03561_)
  );
  al_nand2 _09243_ (
    .a(TM1),
    .b(\DFF_1453.Q ),
    .y(_03562_)
  );
  al_nand3 _09244_ (
    .a(\DFF_1485.Q ),
    .b(_03561_),
    .c(_03562_),
    .y(_03563_)
  );
  al_nand2ft _09245_ (
    .a(TM1),
    .b(\DFF_1453.Q ),
    .y(_03564_)
  );
  al_and2ft _09246_ (
    .a(\DFF_1453.Q ),
    .b(TM1),
    .y(_03565_)
  );
  al_and3fft _09247_ (
    .a(\DFF_1485.Q ),
    .b(_03565_),
    .c(_03564_),
    .y(_03566_)
  );
  al_and2ft _09248_ (
    .a(\DFF_1421.Q ),
    .b(\DFF_1389.Q ),
    .y(_03567_)
  );
  al_nand2ft _09249_ (
    .a(\DFF_1389.Q ),
    .b(\DFF_1421.Q ),
    .y(_03568_)
  );
  al_nand2ft _09250_ (
    .a(_03567_),
    .b(_03568_),
    .y(_03569_)
  );
  al_oai21ftf _09251_ (
    .a(_03563_),
    .b(_03566_),
    .c(_03569_),
    .y(_03570_)
  );
  al_nand3ftt _09252_ (
    .a(_03566_),
    .b(_03563_),
    .c(_03569_),
    .y(_03571_)
  );
  al_nand3 _09253_ (
    .a(_00448_),
    .b(_03570_),
    .c(_03571_),
    .y(_03572_)
  );
  al_aoi21 _09254_ (
    .a(TM0),
    .b(\DFF_1330.Q ),
    .c(TM1),
    .y(_03573_)
  );
  al_nand2 _09255_ (
    .a(_03573_),
    .b(_03572_),
    .y(_03574_)
  );
  al_aoi21ttf _09256_ (
    .a(TM0),
    .b(\DFF_1165.Q ),
    .c(TM1),
    .y(_03575_)
  );
  al_and2 _09257_ (
    .a(_03575_),
    .b(_03083_),
    .y(_03576_)
  );
  al_nor3fft _09258_ (
    .a(RESET),
    .b(_03574_),
    .c(_03576_),
    .y(\DFF_1197.D )
  );
  al_or2 _09259_ (
    .a(TM1),
    .b(\DFF_1454.Q ),
    .y(_03577_)
  );
  al_nand2 _09260_ (
    .a(TM1),
    .b(\DFF_1454.Q ),
    .y(_03578_)
  );
  al_nand3 _09261_ (
    .a(\DFF_1486.Q ),
    .b(_03577_),
    .c(_03578_),
    .y(_03579_)
  );
  al_nand2ft _09262_ (
    .a(TM1),
    .b(\DFF_1454.Q ),
    .y(_03580_)
  );
  al_and2ft _09263_ (
    .a(\DFF_1454.Q ),
    .b(TM1),
    .y(_03581_)
  );
  al_and3fft _09264_ (
    .a(\DFF_1486.Q ),
    .b(_03581_),
    .c(_03580_),
    .y(_03582_)
  );
  al_and2ft _09265_ (
    .a(\DFF_1422.Q ),
    .b(\DFF_1390.Q ),
    .y(_03583_)
  );
  al_nand2ft _09266_ (
    .a(\DFF_1390.Q ),
    .b(\DFF_1422.Q ),
    .y(_03584_)
  );
  al_nand2ft _09267_ (
    .a(_03583_),
    .b(_03584_),
    .y(_03585_)
  );
  al_oai21ftf _09268_ (
    .a(_03579_),
    .b(_03582_),
    .c(_03585_),
    .y(_03586_)
  );
  al_nand3ftt _09269_ (
    .a(_03582_),
    .b(_03579_),
    .c(_03585_),
    .y(_03587_)
  );
  al_nand3 _09270_ (
    .a(_00448_),
    .b(_03586_),
    .c(_03587_),
    .y(_03588_)
  );
  al_aoi21 _09271_ (
    .a(TM0),
    .b(\DFF_1329.Q ),
    .c(TM1),
    .y(_03589_)
  );
  al_nand2 _09272_ (
    .a(_03589_),
    .b(_03588_),
    .y(_03590_)
  );
  al_aoi21ttf _09273_ (
    .a(TM0),
    .b(\DFF_1166.Q ),
    .c(TM1),
    .y(_03591_)
  );
  al_and2 _09274_ (
    .a(_03591_),
    .b(_03099_),
    .y(_03592_)
  );
  al_nor3fft _09275_ (
    .a(RESET),
    .b(_03590_),
    .c(_03592_),
    .y(\DFF_1198.D )
  );
  al_or2 _09276_ (
    .a(TM1),
    .b(\DFF_1455.Q ),
    .y(_03593_)
  );
  al_nand2 _09277_ (
    .a(TM1),
    .b(\DFF_1455.Q ),
    .y(_03594_)
  );
  al_nand3 _09278_ (
    .a(\DFF_1487.Q ),
    .b(_03593_),
    .c(_03594_),
    .y(_03595_)
  );
  al_nand2ft _09279_ (
    .a(TM1),
    .b(\DFF_1455.Q ),
    .y(_03596_)
  );
  al_and2ft _09280_ (
    .a(\DFF_1455.Q ),
    .b(TM1),
    .y(_03597_)
  );
  al_and3fft _09281_ (
    .a(\DFF_1487.Q ),
    .b(_03597_),
    .c(_03596_),
    .y(_03598_)
  );
  al_and2ft _09282_ (
    .a(\DFF_1423.Q ),
    .b(\DFF_1391.Q ),
    .y(_03599_)
  );
  al_nand2ft _09283_ (
    .a(\DFF_1391.Q ),
    .b(\DFF_1423.Q ),
    .y(_03600_)
  );
  al_nand2ft _09284_ (
    .a(_03599_),
    .b(_03600_),
    .y(_03601_)
  );
  al_oai21ftf _09285_ (
    .a(_03595_),
    .b(_03598_),
    .c(_03601_),
    .y(_03602_)
  );
  al_nand3ftt _09286_ (
    .a(_03598_),
    .b(_03595_),
    .c(_03601_),
    .y(_03603_)
  );
  al_nand3 _09287_ (
    .a(_00448_),
    .b(_03602_),
    .c(_03603_),
    .y(_03604_)
  );
  al_aoi21 _09288_ (
    .a(TM0),
    .b(\DFF_1328.Q ),
    .c(TM1),
    .y(_03605_)
  );
  al_nand2 _09289_ (
    .a(_03605_),
    .b(_03604_),
    .y(_03606_)
  );
  al_aoi21ttf _09290_ (
    .a(TM0),
    .b(\DFF_1167.Q ),
    .c(TM1),
    .y(_03607_)
  );
  al_and2 _09291_ (
    .a(_03607_),
    .b(_03115_),
    .y(_03608_)
  );
  al_nor3fft _09292_ (
    .a(RESET),
    .b(_03606_),
    .c(_03608_),
    .y(\DFF_1199.D )
  );
  al_nor2 _09293_ (
    .a(\DFF_1424.Q ),
    .b(\DFF_1456.Q ),
    .y(_03609_)
  );
  al_and2 _09294_ (
    .a(\DFF_1424.Q ),
    .b(\DFF_1456.Q ),
    .y(_03610_)
  );
  al_and2ft _09295_ (
    .a(\DFF_1392.Q ),
    .b(\DFF_1488.Q ),
    .y(_03611_)
  );
  al_nand2ft _09296_ (
    .a(\DFF_1488.Q ),
    .b(\DFF_1392.Q ),
    .y(_03612_)
  );
  al_nand2ft _09297_ (
    .a(_03611_),
    .b(_03612_),
    .y(_03613_)
  );
  al_oa21ttf _09298_ (
    .a(_03609_),
    .b(_03610_),
    .c(_03613_),
    .y(_03614_)
  );
  al_nand3fft _09299_ (
    .a(_03609_),
    .b(_03610_),
    .c(_03613_),
    .y(_03615_)
  );
  al_and3fft _09300_ (
    .a(TM0),
    .b(_03614_),
    .c(_03615_),
    .y(_03616_)
  );
  al_nand2 _09301_ (
    .a(TM0),
    .b(\DFF_1327.Q ),
    .y(_03617_)
  );
  al_or3fft _09302_ (
    .a(_01652_),
    .b(_03617_),
    .c(_03616_),
    .y(_03618_)
  );
  al_and2 _09303_ (
    .a(TM0),
    .b(\DFF_1168.Q ),
    .y(_03619_)
  );
  al_and3fft _09304_ (
    .a(_03619_),
    .b(_03127_),
    .c(TM1),
    .y(_03620_)
  );
  al_nor3fft _09305_ (
    .a(RESET),
    .b(_03618_),
    .c(_03620_),
    .y(\DFF_1200.D )
  );
  al_nor2 _09306_ (
    .a(\DFF_1425.Q ),
    .b(\DFF_1457.Q ),
    .y(_03621_)
  );
  al_and2 _09307_ (
    .a(\DFF_1425.Q ),
    .b(\DFF_1457.Q ),
    .y(_03622_)
  );
  al_and2ft _09308_ (
    .a(\DFF_1393.Q ),
    .b(\DFF_1489.Q ),
    .y(_03623_)
  );
  al_nand2ft _09309_ (
    .a(\DFF_1489.Q ),
    .b(\DFF_1393.Q ),
    .y(_03624_)
  );
  al_nand2ft _09310_ (
    .a(_03623_),
    .b(_03624_),
    .y(_03625_)
  );
  al_oa21ttf _09311_ (
    .a(_03621_),
    .b(_03622_),
    .c(_03625_),
    .y(_03626_)
  );
  al_nand3fft _09312_ (
    .a(_03621_),
    .b(_03622_),
    .c(_03625_),
    .y(_03627_)
  );
  al_and3fft _09313_ (
    .a(TM0),
    .b(_03626_),
    .c(_03627_),
    .y(_03628_)
  );
  al_nand2 _09314_ (
    .a(TM0),
    .b(\DFF_1326.Q ),
    .y(_03629_)
  );
  al_or3fft _09315_ (
    .a(_01652_),
    .b(_03629_),
    .c(_03628_),
    .y(_03630_)
  );
  al_and2 _09316_ (
    .a(TM0),
    .b(\DFF_1169.Q ),
    .y(_03631_)
  );
  al_and3fft _09317_ (
    .a(_03631_),
    .b(_03139_),
    .c(TM1),
    .y(_03632_)
  );
  al_nor3fft _09318_ (
    .a(RESET),
    .b(_03630_),
    .c(_03632_),
    .y(\DFF_1201.D )
  );
  al_nor2 _09319_ (
    .a(\DFF_1426.Q ),
    .b(\DFF_1458.Q ),
    .y(_03633_)
  );
  al_and2 _09320_ (
    .a(\DFF_1426.Q ),
    .b(\DFF_1458.Q ),
    .y(_03634_)
  );
  al_and2ft _09321_ (
    .a(\DFF_1394.Q ),
    .b(\DFF_1490.Q ),
    .y(_03635_)
  );
  al_nand2ft _09322_ (
    .a(\DFF_1490.Q ),
    .b(\DFF_1394.Q ),
    .y(_03636_)
  );
  al_nand2ft _09323_ (
    .a(_03635_),
    .b(_03636_),
    .y(_03637_)
  );
  al_oa21ttf _09324_ (
    .a(_03633_),
    .b(_03634_),
    .c(_03637_),
    .y(_03638_)
  );
  al_nand3fft _09325_ (
    .a(_03633_),
    .b(_03634_),
    .c(_03637_),
    .y(_03639_)
  );
  al_and3fft _09326_ (
    .a(TM0),
    .b(_03638_),
    .c(_03639_),
    .y(_03640_)
  );
  al_nand2 _09327_ (
    .a(TM0),
    .b(\DFF_1325.Q ),
    .y(_03641_)
  );
  al_or3fft _09328_ (
    .a(_01652_),
    .b(_03641_),
    .c(_03640_),
    .y(_03642_)
  );
  al_and2 _09329_ (
    .a(TM0),
    .b(\DFF_1170.Q ),
    .y(_03643_)
  );
  al_and3fft _09330_ (
    .a(_03643_),
    .b(_03151_),
    .c(TM1),
    .y(_03644_)
  );
  al_nor3fft _09331_ (
    .a(RESET),
    .b(_03642_),
    .c(_03644_),
    .y(\DFF_1202.D )
  );
  al_nor2 _09332_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_1459.Q ),
    .y(_03645_)
  );
  al_and2 _09333_ (
    .a(\DFF_1427.Q ),
    .b(\DFF_1459.Q ),
    .y(_03646_)
  );
  al_and2ft _09334_ (
    .a(\DFF_1395.Q ),
    .b(\DFF_1491.Q ),
    .y(_03647_)
  );
  al_nand2ft _09335_ (
    .a(\DFF_1491.Q ),
    .b(\DFF_1395.Q ),
    .y(_03648_)
  );
  al_nand2ft _09336_ (
    .a(_03647_),
    .b(_03648_),
    .y(_03649_)
  );
  al_oa21ttf _09337_ (
    .a(_03645_),
    .b(_03646_),
    .c(_03649_),
    .y(_03650_)
  );
  al_nand3fft _09338_ (
    .a(_03645_),
    .b(_03646_),
    .c(_03649_),
    .y(_03651_)
  );
  al_and3fft _09339_ (
    .a(TM0),
    .b(_03650_),
    .c(_03651_),
    .y(_03652_)
  );
  al_nand2 _09340_ (
    .a(TM0),
    .b(\DFF_1324.Q ),
    .y(_03653_)
  );
  al_or3fft _09341_ (
    .a(_01652_),
    .b(_03653_),
    .c(_03652_),
    .y(_03654_)
  );
  al_and2 _09342_ (
    .a(TM0),
    .b(\DFF_1171.Q ),
    .y(_03655_)
  );
  al_and3fft _09343_ (
    .a(_03655_),
    .b(_03163_),
    .c(TM1),
    .y(_03656_)
  );
  al_nor3fft _09344_ (
    .a(RESET),
    .b(_03654_),
    .c(_03656_),
    .y(\DFF_1203.D )
  );
  al_nor2 _09345_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_1460.Q ),
    .y(_03657_)
  );
  al_and2 _09346_ (
    .a(\DFF_1428.Q ),
    .b(\DFF_1460.Q ),
    .y(_03658_)
  );
  al_and2ft _09347_ (
    .a(\DFF_1396.Q ),
    .b(\DFF_1492.Q ),
    .y(_03659_)
  );
  al_nand2ft _09348_ (
    .a(\DFF_1492.Q ),
    .b(\DFF_1396.Q ),
    .y(_03660_)
  );
  al_nand2ft _09349_ (
    .a(_03659_),
    .b(_03660_),
    .y(_03661_)
  );
  al_oa21ttf _09350_ (
    .a(_03657_),
    .b(_03658_),
    .c(_03661_),
    .y(_03662_)
  );
  al_nand3fft _09351_ (
    .a(_03657_),
    .b(_03658_),
    .c(_03661_),
    .y(_03663_)
  );
  al_and3fft _09352_ (
    .a(TM0),
    .b(_03662_),
    .c(_03663_),
    .y(_03664_)
  );
  al_nand2 _09353_ (
    .a(TM0),
    .b(\DFF_1323.Q ),
    .y(_03665_)
  );
  al_or3fft _09354_ (
    .a(_01652_),
    .b(_03665_),
    .c(_03664_),
    .y(_03666_)
  );
  al_and2 _09355_ (
    .a(TM0),
    .b(\DFF_1172.Q ),
    .y(_03667_)
  );
  al_and3fft _09356_ (
    .a(_03667_),
    .b(_03175_),
    .c(TM1),
    .y(_03668_)
  );
  al_nor3fft _09357_ (
    .a(RESET),
    .b(_03666_),
    .c(_03668_),
    .y(\DFF_1204.D )
  );
  al_nor2 _09358_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_1461.Q ),
    .y(_03669_)
  );
  al_and2 _09359_ (
    .a(\DFF_1429.Q ),
    .b(\DFF_1461.Q ),
    .y(_03670_)
  );
  al_and2ft _09360_ (
    .a(\DFF_1397.Q ),
    .b(\DFF_1493.Q ),
    .y(_03671_)
  );
  al_nand2ft _09361_ (
    .a(\DFF_1493.Q ),
    .b(\DFF_1397.Q ),
    .y(_03672_)
  );
  al_nand2ft _09362_ (
    .a(_03671_),
    .b(_03672_),
    .y(_03673_)
  );
  al_oa21ttf _09363_ (
    .a(_03669_),
    .b(_03670_),
    .c(_03673_),
    .y(_03674_)
  );
  al_nand3fft _09364_ (
    .a(_03669_),
    .b(_03670_),
    .c(_03673_),
    .y(_03675_)
  );
  al_and3fft _09365_ (
    .a(TM0),
    .b(_03674_),
    .c(_03675_),
    .y(_03676_)
  );
  al_nand2 _09366_ (
    .a(TM0),
    .b(\DFF_1322.Q ),
    .y(_03677_)
  );
  al_or3fft _09367_ (
    .a(_01652_),
    .b(_03677_),
    .c(_03676_),
    .y(_03678_)
  );
  al_and2 _09368_ (
    .a(TM0),
    .b(\DFF_1173.Q ),
    .y(_03679_)
  );
  al_and3fft _09369_ (
    .a(_03679_),
    .b(_03187_),
    .c(TM1),
    .y(_03680_)
  );
  al_nor3fft _09370_ (
    .a(RESET),
    .b(_03678_),
    .c(_03680_),
    .y(\DFF_1205.D )
  );
  al_nor2 _09371_ (
    .a(\DFF_1430.Q ),
    .b(\DFF_1462.Q ),
    .y(_03681_)
  );
  al_and2 _09372_ (
    .a(\DFF_1430.Q ),
    .b(\DFF_1462.Q ),
    .y(_03682_)
  );
  al_and2ft _09373_ (
    .a(\DFF_1398.Q ),
    .b(\DFF_1494.Q ),
    .y(_03683_)
  );
  al_nand2ft _09374_ (
    .a(\DFF_1494.Q ),
    .b(\DFF_1398.Q ),
    .y(_03684_)
  );
  al_nand2ft _09375_ (
    .a(_03683_),
    .b(_03684_),
    .y(_03685_)
  );
  al_oa21ttf _09376_ (
    .a(_03681_),
    .b(_03682_),
    .c(_03685_),
    .y(_03686_)
  );
  al_nand3fft _09377_ (
    .a(_03681_),
    .b(_03682_),
    .c(_03685_),
    .y(_03687_)
  );
  al_and3fft _09378_ (
    .a(TM0),
    .b(_03686_),
    .c(_03687_),
    .y(_03688_)
  );
  al_nand2 _09379_ (
    .a(TM0),
    .b(\DFF_1321.Q ),
    .y(_03689_)
  );
  al_or3fft _09380_ (
    .a(_01652_),
    .b(_03689_),
    .c(_03688_),
    .y(_03690_)
  );
  al_and2 _09381_ (
    .a(TM0),
    .b(\DFF_1174.Q ),
    .y(_03691_)
  );
  al_and3fft _09382_ (
    .a(_03691_),
    .b(_03199_),
    .c(TM1),
    .y(_03692_)
  );
  al_nor3fft _09383_ (
    .a(RESET),
    .b(_03690_),
    .c(_03692_),
    .y(\DFF_1206.D )
  );
  al_nor2 _09384_ (
    .a(\DFF_1431.Q ),
    .b(\DFF_1463.Q ),
    .y(_03693_)
  );
  al_and2 _09385_ (
    .a(\DFF_1431.Q ),
    .b(\DFF_1463.Q ),
    .y(_03694_)
  );
  al_and2ft _09386_ (
    .a(\DFF_1399.Q ),
    .b(\DFF_1495.Q ),
    .y(_03695_)
  );
  al_nand2ft _09387_ (
    .a(\DFF_1495.Q ),
    .b(\DFF_1399.Q ),
    .y(_03696_)
  );
  al_nand2ft _09388_ (
    .a(_03695_),
    .b(_03696_),
    .y(_03697_)
  );
  al_oa21ttf _09389_ (
    .a(_03693_),
    .b(_03694_),
    .c(_03697_),
    .y(_03698_)
  );
  al_nand3fft _09390_ (
    .a(_03693_),
    .b(_03694_),
    .c(_03697_),
    .y(_03699_)
  );
  al_and3fft _09391_ (
    .a(TM0),
    .b(_03698_),
    .c(_03699_),
    .y(_03700_)
  );
  al_nand2 _09392_ (
    .a(TM0),
    .b(\DFF_1320.Q ),
    .y(_03701_)
  );
  al_or3fft _09393_ (
    .a(_01652_),
    .b(_03701_),
    .c(_03700_),
    .y(_03702_)
  );
  al_and2 _09394_ (
    .a(TM0),
    .b(\DFF_1175.Q ),
    .y(_03703_)
  );
  al_and3fft _09395_ (
    .a(_03703_),
    .b(_03211_),
    .c(TM1),
    .y(_03704_)
  );
  al_nor3fft _09396_ (
    .a(RESET),
    .b(_03702_),
    .c(_03704_),
    .y(\DFF_1207.D )
  );
  al_nor2 _09397_ (
    .a(\DFF_1432.Q ),
    .b(\DFF_1464.Q ),
    .y(_03705_)
  );
  al_and2 _09398_ (
    .a(\DFF_1432.Q ),
    .b(\DFF_1464.Q ),
    .y(_03706_)
  );
  al_and2ft _09399_ (
    .a(\DFF_1400.Q ),
    .b(\DFF_1496.Q ),
    .y(_03707_)
  );
  al_nand2ft _09400_ (
    .a(\DFF_1496.Q ),
    .b(\DFF_1400.Q ),
    .y(_03708_)
  );
  al_nand2ft _09401_ (
    .a(_03707_),
    .b(_03708_),
    .y(_03709_)
  );
  al_oa21ttf _09402_ (
    .a(_03705_),
    .b(_03706_),
    .c(_03709_),
    .y(_03710_)
  );
  al_nand3fft _09403_ (
    .a(_03705_),
    .b(_03706_),
    .c(_03709_),
    .y(_03711_)
  );
  al_and3fft _09404_ (
    .a(TM0),
    .b(_03710_),
    .c(_03711_),
    .y(_03712_)
  );
  al_nand2 _09405_ (
    .a(TM0),
    .b(\DFF_1319.Q ),
    .y(_03713_)
  );
  al_or3fft _09406_ (
    .a(_01652_),
    .b(_03713_),
    .c(_03712_),
    .y(_03714_)
  );
  al_and2 _09407_ (
    .a(TM0),
    .b(\DFF_1176.Q ),
    .y(_03715_)
  );
  al_and3fft _09408_ (
    .a(_03715_),
    .b(_03223_),
    .c(TM1),
    .y(_03716_)
  );
  al_nor3fft _09409_ (
    .a(RESET),
    .b(_03714_),
    .c(_03716_),
    .y(\DFF_1208.D )
  );
  al_nor2 _09410_ (
    .a(\DFF_1433.Q ),
    .b(\DFF_1465.Q ),
    .y(_03717_)
  );
  al_and2 _09411_ (
    .a(\DFF_1433.Q ),
    .b(\DFF_1465.Q ),
    .y(_03718_)
  );
  al_and2ft _09412_ (
    .a(\DFF_1401.Q ),
    .b(\DFF_1497.Q ),
    .y(_03719_)
  );
  al_nand2ft _09413_ (
    .a(\DFF_1497.Q ),
    .b(\DFF_1401.Q ),
    .y(_03720_)
  );
  al_nand2ft _09414_ (
    .a(_03719_),
    .b(_03720_),
    .y(_03721_)
  );
  al_oa21ttf _09415_ (
    .a(_03717_),
    .b(_03718_),
    .c(_03721_),
    .y(_03722_)
  );
  al_nand3fft _09416_ (
    .a(_03717_),
    .b(_03718_),
    .c(_03721_),
    .y(_03723_)
  );
  al_and3fft _09417_ (
    .a(TM0),
    .b(_03722_),
    .c(_03723_),
    .y(_03724_)
  );
  al_nand2 _09418_ (
    .a(TM0),
    .b(\DFF_1318.Q ),
    .y(_03725_)
  );
  al_or3fft _09419_ (
    .a(_01652_),
    .b(_03725_),
    .c(_03724_),
    .y(_03726_)
  );
  al_and2 _09420_ (
    .a(TM0),
    .b(\DFF_1177.Q ),
    .y(_03727_)
  );
  al_and3fft _09421_ (
    .a(_03727_),
    .b(_03235_),
    .c(TM1),
    .y(_03728_)
  );
  al_nor3fft _09422_ (
    .a(RESET),
    .b(_03726_),
    .c(_03728_),
    .y(\DFF_1209.D )
  );
  al_nor2 _09423_ (
    .a(\DFF_1434.Q ),
    .b(\DFF_1466.Q ),
    .y(_03729_)
  );
  al_and2 _09424_ (
    .a(\DFF_1434.Q ),
    .b(\DFF_1466.Q ),
    .y(_03730_)
  );
  al_and2ft _09425_ (
    .a(\DFF_1402.Q ),
    .b(\DFF_1498.Q ),
    .y(_03731_)
  );
  al_nand2ft _09426_ (
    .a(\DFF_1498.Q ),
    .b(\DFF_1402.Q ),
    .y(_03732_)
  );
  al_nand2ft _09427_ (
    .a(_03731_),
    .b(_03732_),
    .y(_03733_)
  );
  al_oa21ttf _09428_ (
    .a(_03729_),
    .b(_03730_),
    .c(_03733_),
    .y(_03734_)
  );
  al_nand3fft _09429_ (
    .a(_03729_),
    .b(_03730_),
    .c(_03733_),
    .y(_03735_)
  );
  al_and3fft _09430_ (
    .a(TM0),
    .b(_03734_),
    .c(_03735_),
    .y(_03736_)
  );
  al_nand2 _09431_ (
    .a(TM0),
    .b(\DFF_1317.Q ),
    .y(_03737_)
  );
  al_or3fft _09432_ (
    .a(_01652_),
    .b(_03737_),
    .c(_03736_),
    .y(_03738_)
  );
  al_and2 _09433_ (
    .a(TM0),
    .b(\DFF_1178.Q ),
    .y(_03739_)
  );
  al_and3fft _09434_ (
    .a(_03739_),
    .b(_03247_),
    .c(TM1),
    .y(_03740_)
  );
  al_nor3fft _09435_ (
    .a(RESET),
    .b(_03738_),
    .c(_03740_),
    .y(\DFF_1210.D )
  );
  al_nor2 _09436_ (
    .a(\DFF_1435.Q ),
    .b(\DFF_1467.Q ),
    .y(_03741_)
  );
  al_and2 _09437_ (
    .a(\DFF_1435.Q ),
    .b(\DFF_1467.Q ),
    .y(_03742_)
  );
  al_and2ft _09438_ (
    .a(\DFF_1403.Q ),
    .b(\DFF_1499.Q ),
    .y(_03743_)
  );
  al_nand2ft _09439_ (
    .a(\DFF_1499.Q ),
    .b(\DFF_1403.Q ),
    .y(_03744_)
  );
  al_nand2ft _09440_ (
    .a(_03743_),
    .b(_03744_),
    .y(_03745_)
  );
  al_oa21ttf _09441_ (
    .a(_03741_),
    .b(_03742_),
    .c(_03745_),
    .y(_03746_)
  );
  al_nand3fft _09442_ (
    .a(_03741_),
    .b(_03742_),
    .c(_03745_),
    .y(_03747_)
  );
  al_and3fft _09443_ (
    .a(TM0),
    .b(_03746_),
    .c(_03747_),
    .y(_03748_)
  );
  al_nand2 _09444_ (
    .a(TM0),
    .b(\DFF_1316.Q ),
    .y(_03749_)
  );
  al_or3fft _09445_ (
    .a(_01652_),
    .b(_03749_),
    .c(_03748_),
    .y(_03750_)
  );
  al_and2 _09446_ (
    .a(TM0),
    .b(\DFF_1179.Q ),
    .y(_03751_)
  );
  al_and3fft _09447_ (
    .a(_03751_),
    .b(_03259_),
    .c(TM1),
    .y(_03752_)
  );
  al_nor3fft _09448_ (
    .a(RESET),
    .b(_03750_),
    .c(_03752_),
    .y(\DFF_1211.D )
  );
  al_nor2 _09449_ (
    .a(\DFF_1436.Q ),
    .b(\DFF_1468.Q ),
    .y(_03753_)
  );
  al_and2 _09450_ (
    .a(\DFF_1436.Q ),
    .b(\DFF_1468.Q ),
    .y(_03754_)
  );
  al_and2ft _09451_ (
    .a(\DFF_1404.Q ),
    .b(\DFF_1500.Q ),
    .y(_03755_)
  );
  al_nand2ft _09452_ (
    .a(\DFF_1500.Q ),
    .b(\DFF_1404.Q ),
    .y(_03756_)
  );
  al_nand2ft _09453_ (
    .a(_03755_),
    .b(_03756_),
    .y(_03757_)
  );
  al_oa21ttf _09454_ (
    .a(_03753_),
    .b(_03754_),
    .c(_03757_),
    .y(_03758_)
  );
  al_nand3fft _09455_ (
    .a(_03753_),
    .b(_03754_),
    .c(_03757_),
    .y(_03759_)
  );
  al_and3fft _09456_ (
    .a(TM0),
    .b(_03758_),
    .c(_03759_),
    .y(_03760_)
  );
  al_nand2 _09457_ (
    .a(TM0),
    .b(\DFF_1315.Q ),
    .y(_03761_)
  );
  al_or3fft _09458_ (
    .a(_01652_),
    .b(_03761_),
    .c(_03760_),
    .y(_03762_)
  );
  al_and2 _09459_ (
    .a(TM0),
    .b(\DFF_1180.Q ),
    .y(_03763_)
  );
  al_and3fft _09460_ (
    .a(_03763_),
    .b(_03271_),
    .c(TM1),
    .y(_03764_)
  );
  al_nor3fft _09461_ (
    .a(RESET),
    .b(_03762_),
    .c(_03764_),
    .y(\DFF_1212.D )
  );
  al_nor2 _09462_ (
    .a(\DFF_1437.Q ),
    .b(\DFF_1469.Q ),
    .y(_03765_)
  );
  al_and2 _09463_ (
    .a(\DFF_1437.Q ),
    .b(\DFF_1469.Q ),
    .y(_03766_)
  );
  al_and2ft _09464_ (
    .a(\DFF_1405.Q ),
    .b(\DFF_1501.Q ),
    .y(_03767_)
  );
  al_nand2ft _09465_ (
    .a(\DFF_1501.Q ),
    .b(\DFF_1405.Q ),
    .y(_03768_)
  );
  al_nand2ft _09466_ (
    .a(_03767_),
    .b(_03768_),
    .y(_03769_)
  );
  al_oa21ttf _09467_ (
    .a(_03765_),
    .b(_03766_),
    .c(_03769_),
    .y(_03770_)
  );
  al_nand3fft _09468_ (
    .a(_03765_),
    .b(_03766_),
    .c(_03769_),
    .y(_03771_)
  );
  al_and3fft _09469_ (
    .a(TM0),
    .b(_03770_),
    .c(_03771_),
    .y(_03772_)
  );
  al_nand2 _09470_ (
    .a(TM0),
    .b(\DFF_1314.Q ),
    .y(_03773_)
  );
  al_or3fft _09471_ (
    .a(_01652_),
    .b(_03773_),
    .c(_03772_),
    .y(_03774_)
  );
  al_and2 _09472_ (
    .a(TM0),
    .b(\DFF_1181.Q ),
    .y(_03775_)
  );
  al_and3fft _09473_ (
    .a(_03775_),
    .b(_03283_),
    .c(TM1),
    .y(_03776_)
  );
  al_nor3fft _09474_ (
    .a(RESET),
    .b(_03774_),
    .c(_03776_),
    .y(\DFF_1213.D )
  );
  al_nor2 _09475_ (
    .a(\DFF_1438.Q ),
    .b(\DFF_1470.Q ),
    .y(_03777_)
  );
  al_and2 _09476_ (
    .a(\DFF_1438.Q ),
    .b(\DFF_1470.Q ),
    .y(_03778_)
  );
  al_and2ft _09477_ (
    .a(\DFF_1406.Q ),
    .b(\DFF_1502.Q ),
    .y(_03779_)
  );
  al_nand2ft _09478_ (
    .a(\DFF_1502.Q ),
    .b(\DFF_1406.Q ),
    .y(_03780_)
  );
  al_nand2ft _09479_ (
    .a(_03779_),
    .b(_03780_),
    .y(_03781_)
  );
  al_oa21ttf _09480_ (
    .a(_03777_),
    .b(_03778_),
    .c(_03781_),
    .y(_03782_)
  );
  al_nand3fft _09481_ (
    .a(_03777_),
    .b(_03778_),
    .c(_03781_),
    .y(_03783_)
  );
  al_and3fft _09482_ (
    .a(TM0),
    .b(_03782_),
    .c(_03783_),
    .y(_03784_)
  );
  al_nand2 _09483_ (
    .a(TM0),
    .b(\DFF_1313.Q ),
    .y(_03785_)
  );
  al_or3fft _09484_ (
    .a(_01652_),
    .b(_03785_),
    .c(_03784_),
    .y(_03786_)
  );
  al_and2 _09485_ (
    .a(TM0),
    .b(\DFF_1182.Q ),
    .y(_03787_)
  );
  al_and3fft _09486_ (
    .a(_03787_),
    .b(_03295_),
    .c(TM1),
    .y(_03788_)
  );
  al_nor3fft _09487_ (
    .a(RESET),
    .b(_03786_),
    .c(_03788_),
    .y(\DFF_1214.D )
  );
  al_nor2 _09488_ (
    .a(\DFF_1439.Q ),
    .b(\DFF_1471.Q ),
    .y(_03789_)
  );
  al_and2 _09489_ (
    .a(\DFF_1439.Q ),
    .b(\DFF_1471.Q ),
    .y(_03790_)
  );
  al_and2ft _09490_ (
    .a(\DFF_1407.Q ),
    .b(\DFF_1503.Q ),
    .y(_03791_)
  );
  al_nand2ft _09491_ (
    .a(\DFF_1503.Q ),
    .b(\DFF_1407.Q ),
    .y(_03792_)
  );
  al_nand2ft _09492_ (
    .a(_03791_),
    .b(_03792_),
    .y(_03793_)
  );
  al_oa21ttf _09493_ (
    .a(_03789_),
    .b(_03790_),
    .c(_03793_),
    .y(_03794_)
  );
  al_nand3fft _09494_ (
    .a(_03789_),
    .b(_03790_),
    .c(_03793_),
    .y(_03795_)
  );
  al_and3fft _09495_ (
    .a(TM0),
    .b(_03794_),
    .c(_03795_),
    .y(_03796_)
  );
  al_nand2 _09496_ (
    .a(TM0),
    .b(\DFF_1312.Q ),
    .y(_03797_)
  );
  al_or3fft _09497_ (
    .a(_01652_),
    .b(_03797_),
    .c(_03796_),
    .y(_03798_)
  );
  al_and2 _09498_ (
    .a(TM0),
    .b(\DFF_1183.Q ),
    .y(_03799_)
  );
  al_and3fft _09499_ (
    .a(_03799_),
    .b(_03307_),
    .c(TM1),
    .y(_03800_)
  );
  al_nor3fft _09500_ (
    .a(RESET),
    .b(_03798_),
    .c(_03800_),
    .y(\DFF_1215.D )
  );
  al_and2 _09501_ (
    .a(RESET),
    .b(\DFF_1184.Q ),
    .y(\DFF_1216.D )
  );
  al_and2 _09502_ (
    .a(RESET),
    .b(\DFF_1185.Q ),
    .y(\DFF_1217.D )
  );
  al_and2 _09503_ (
    .a(RESET),
    .b(\DFF_1186.Q ),
    .y(\DFF_1218.D )
  );
  al_and2 _09504_ (
    .a(RESET),
    .b(\DFF_1187.Q ),
    .y(\DFF_1219.D )
  );
  al_and2 _09505_ (
    .a(RESET),
    .b(\DFF_1188.Q ),
    .y(\DFF_1220.D )
  );
  al_and2 _09506_ (
    .a(RESET),
    .b(\DFF_1189.Q ),
    .y(\DFF_1221.D )
  );
  al_and2 _09507_ (
    .a(RESET),
    .b(\DFF_1190.Q ),
    .y(\DFF_1222.D )
  );
  al_and2 _09508_ (
    .a(RESET),
    .b(\DFF_1191.Q ),
    .y(\DFF_1223.D )
  );
  al_and2 _09509_ (
    .a(RESET),
    .b(\DFF_1192.Q ),
    .y(\DFF_1224.D )
  );
  al_and2 _09510_ (
    .a(RESET),
    .b(\DFF_1193.Q ),
    .y(\DFF_1225.D )
  );
  al_and2 _09511_ (
    .a(RESET),
    .b(\DFF_1194.Q ),
    .y(\DFF_1226.D )
  );
  al_and2 _09512_ (
    .a(RESET),
    .b(\DFF_1195.Q ),
    .y(\DFF_1227.D )
  );
  al_and2 _09513_ (
    .a(RESET),
    .b(\DFF_1196.Q ),
    .y(\DFF_1228.D )
  );
  al_and2 _09514_ (
    .a(RESET),
    .b(\DFF_1197.Q ),
    .y(\DFF_1229.D )
  );
  al_and2 _09515_ (
    .a(RESET),
    .b(\DFF_1198.Q ),
    .y(\DFF_1230.D )
  );
  al_and2 _09516_ (
    .a(RESET),
    .b(\DFF_1199.Q ),
    .y(\DFF_1231.D )
  );
  al_and2 _09517_ (
    .a(RESET),
    .b(\DFF_1200.Q ),
    .y(\DFF_1232.D )
  );
  al_and2 _09518_ (
    .a(RESET),
    .b(\DFF_1201.Q ),
    .y(\DFF_1233.D )
  );
  al_and2 _09519_ (
    .a(RESET),
    .b(\DFF_1202.Q ),
    .y(\DFF_1234.D )
  );
  al_and2 _09520_ (
    .a(RESET),
    .b(\DFF_1203.Q ),
    .y(\DFF_1235.D )
  );
  al_and2 _09521_ (
    .a(RESET),
    .b(\DFF_1204.Q ),
    .y(\DFF_1236.D )
  );
  al_and2 _09522_ (
    .a(RESET),
    .b(\DFF_1205.Q ),
    .y(\DFF_1237.D )
  );
  al_and2 _09523_ (
    .a(RESET),
    .b(\DFF_1206.Q ),
    .y(\DFF_1238.D )
  );
  al_and2 _09524_ (
    .a(RESET),
    .b(\DFF_1207.Q ),
    .y(\DFF_1239.D )
  );
  al_and2 _09525_ (
    .a(RESET),
    .b(\DFF_1208.Q ),
    .y(\DFF_1240.D )
  );
  al_and2 _09526_ (
    .a(RESET),
    .b(\DFF_1209.Q ),
    .y(\DFF_1241.D )
  );
  al_and2 _09527_ (
    .a(RESET),
    .b(\DFF_1210.Q ),
    .y(\DFF_1242.D )
  );
  al_and2 _09528_ (
    .a(RESET),
    .b(\DFF_1211.Q ),
    .y(\DFF_1243.D )
  );
  al_and2 _09529_ (
    .a(RESET),
    .b(\DFF_1212.Q ),
    .y(\DFF_1244.D )
  );
  al_and2 _09530_ (
    .a(RESET),
    .b(\DFF_1213.Q ),
    .y(\DFF_1245.D )
  );
  al_and2 _09531_ (
    .a(RESET),
    .b(\DFF_1214.Q ),
    .y(\DFF_1246.D )
  );
  al_and2 _09532_ (
    .a(RESET),
    .b(\DFF_1215.Q ),
    .y(\DFF_1247.D )
  );
  al_and2 _09533_ (
    .a(RESET),
    .b(\DFF_1216.Q ),
    .y(\DFF_1248.D )
  );
  al_and2 _09534_ (
    .a(RESET),
    .b(\DFF_1217.Q ),
    .y(\DFF_1249.D )
  );
  al_and2 _09535_ (
    .a(RESET),
    .b(\DFF_1218.Q ),
    .y(\DFF_1250.D )
  );
  al_and2 _09536_ (
    .a(RESET),
    .b(\DFF_1219.Q ),
    .y(\DFF_1251.D )
  );
  al_and2 _09537_ (
    .a(RESET),
    .b(\DFF_1220.Q ),
    .y(\DFF_1252.D )
  );
  al_and2 _09538_ (
    .a(RESET),
    .b(\DFF_1221.Q ),
    .y(\DFF_1253.D )
  );
  al_and2 _09539_ (
    .a(RESET),
    .b(\DFF_1222.Q ),
    .y(\DFF_1254.D )
  );
  al_and2 _09540_ (
    .a(RESET),
    .b(\DFF_1223.Q ),
    .y(\DFF_1255.D )
  );
  al_and2 _09541_ (
    .a(RESET),
    .b(\DFF_1224.Q ),
    .y(\DFF_1256.D )
  );
  al_and2 _09542_ (
    .a(RESET),
    .b(\DFF_1225.Q ),
    .y(\DFF_1257.D )
  );
  al_and2 _09543_ (
    .a(RESET),
    .b(\DFF_1226.Q ),
    .y(\DFF_1258.D )
  );
  al_and2 _09544_ (
    .a(RESET),
    .b(\DFF_1227.Q ),
    .y(\DFF_1259.D )
  );
  al_and2 _09545_ (
    .a(RESET),
    .b(\DFF_1228.Q ),
    .y(\DFF_1260.D )
  );
  al_and2 _09546_ (
    .a(RESET),
    .b(\DFF_1229.Q ),
    .y(\DFF_1261.D )
  );
  al_and2 _09547_ (
    .a(RESET),
    .b(\DFF_1230.Q ),
    .y(\DFF_1262.D )
  );
  al_and2 _09548_ (
    .a(RESET),
    .b(\DFF_1231.Q ),
    .y(\DFF_1263.D )
  );
  al_and2 _09549_ (
    .a(RESET),
    .b(\DFF_1232.Q ),
    .y(\DFF_1264.D )
  );
  al_and2 _09550_ (
    .a(RESET),
    .b(\DFF_1233.Q ),
    .y(\DFF_1265.D )
  );
  al_and2 _09551_ (
    .a(RESET),
    .b(\DFF_1234.Q ),
    .y(\DFF_1266.D )
  );
  al_and2 _09552_ (
    .a(RESET),
    .b(\DFF_1235.Q ),
    .y(\DFF_1267.D )
  );
  al_and2 _09553_ (
    .a(RESET),
    .b(\DFF_1236.Q ),
    .y(\DFF_1268.D )
  );
  al_and2 _09554_ (
    .a(RESET),
    .b(\DFF_1237.Q ),
    .y(\DFF_1269.D )
  );
  al_and2 _09555_ (
    .a(RESET),
    .b(\DFF_1238.Q ),
    .y(\DFF_1270.D )
  );
  al_and2 _09556_ (
    .a(RESET),
    .b(\DFF_1239.Q ),
    .y(\DFF_1271.D )
  );
  al_and2 _09557_ (
    .a(RESET),
    .b(\DFF_1240.Q ),
    .y(\DFF_1272.D )
  );
  al_and2 _09558_ (
    .a(RESET),
    .b(\DFF_1241.Q ),
    .y(\DFF_1273.D )
  );
  al_and2 _09559_ (
    .a(RESET),
    .b(\DFF_1242.Q ),
    .y(\DFF_1274.D )
  );
  al_and2 _09560_ (
    .a(RESET),
    .b(\DFF_1243.Q ),
    .y(\DFF_1275.D )
  );
  al_and2 _09561_ (
    .a(RESET),
    .b(\DFF_1244.Q ),
    .y(\DFF_1276.D )
  );
  al_and2 _09562_ (
    .a(RESET),
    .b(\DFF_1245.Q ),
    .y(\DFF_1277.D )
  );
  al_and2 _09563_ (
    .a(RESET),
    .b(\DFF_1246.Q ),
    .y(\DFF_1278.D )
  );
  al_and2 _09564_ (
    .a(RESET),
    .b(\DFF_1247.Q ),
    .y(\DFF_1279.D )
  );
  al_and2 _09565_ (
    .a(RESET),
    .b(\DFF_1248.Q ),
    .y(\DFF_1280.D )
  );
  al_and2 _09566_ (
    .a(RESET),
    .b(\DFF_1249.Q ),
    .y(\DFF_1281.D )
  );
  al_and2 _09567_ (
    .a(RESET),
    .b(\DFF_1250.Q ),
    .y(\DFF_1282.D )
  );
  al_and2 _09568_ (
    .a(RESET),
    .b(\DFF_1251.Q ),
    .y(\DFF_1283.D )
  );
  al_and2 _09569_ (
    .a(RESET),
    .b(\DFF_1252.Q ),
    .y(\DFF_1284.D )
  );
  al_and2 _09570_ (
    .a(RESET),
    .b(\DFF_1253.Q ),
    .y(\DFF_1285.D )
  );
  al_and2 _09571_ (
    .a(RESET),
    .b(\DFF_1254.Q ),
    .y(\DFF_1286.D )
  );
  al_and2 _09572_ (
    .a(RESET),
    .b(\DFF_1255.Q ),
    .y(\DFF_1287.D )
  );
  al_and2 _09573_ (
    .a(RESET),
    .b(\DFF_1256.Q ),
    .y(\DFF_1288.D )
  );
  al_and2 _09574_ (
    .a(RESET),
    .b(\DFF_1257.Q ),
    .y(\DFF_1289.D )
  );
  al_and2 _09575_ (
    .a(RESET),
    .b(\DFF_1258.Q ),
    .y(\DFF_1290.D )
  );
  al_and2 _09576_ (
    .a(RESET),
    .b(\DFF_1259.Q ),
    .y(\DFF_1291.D )
  );
  al_and2 _09577_ (
    .a(RESET),
    .b(\DFF_1260.Q ),
    .y(\DFF_1292.D )
  );
  al_and2 _09578_ (
    .a(RESET),
    .b(\DFF_1261.Q ),
    .y(\DFF_1293.D )
  );
  al_and2 _09579_ (
    .a(RESET),
    .b(\DFF_1262.Q ),
    .y(\DFF_1294.D )
  );
  al_and2 _09580_ (
    .a(RESET),
    .b(\DFF_1263.Q ),
    .y(\DFF_1295.D )
  );
  al_and2 _09581_ (
    .a(RESET),
    .b(\DFF_1264.Q ),
    .y(\DFF_1296.D )
  );
  al_and2 _09582_ (
    .a(RESET),
    .b(\DFF_1265.Q ),
    .y(\DFF_1297.D )
  );
  al_and2 _09583_ (
    .a(RESET),
    .b(\DFF_1266.Q ),
    .y(\DFF_1298.D )
  );
  al_and2 _09584_ (
    .a(RESET),
    .b(\DFF_1267.Q ),
    .y(\DFF_1299.D )
  );
  al_and2 _09585_ (
    .a(RESET),
    .b(\DFF_1268.Q ),
    .y(\DFF_1300.D )
  );
  al_and2 _09586_ (
    .a(RESET),
    .b(\DFF_1269.Q ),
    .y(\DFF_1301.D )
  );
  al_and2 _09587_ (
    .a(RESET),
    .b(\DFF_1270.Q ),
    .y(\DFF_1302.D )
  );
  al_and2 _09588_ (
    .a(RESET),
    .b(\DFF_1271.Q ),
    .y(\DFF_1303.D )
  );
  al_and2 _09589_ (
    .a(RESET),
    .b(\DFF_1272.Q ),
    .y(\DFF_1304.D )
  );
  al_and2 _09590_ (
    .a(RESET),
    .b(\DFF_1273.Q ),
    .y(\DFF_1305.D )
  );
  al_and2 _09591_ (
    .a(RESET),
    .b(\DFF_1274.Q ),
    .y(\DFF_1306.D )
  );
  al_and2 _09592_ (
    .a(RESET),
    .b(\DFF_1275.Q ),
    .y(\DFF_1307.D )
  );
  al_and2 _09593_ (
    .a(RESET),
    .b(\DFF_1276.Q ),
    .y(\DFF_1308.D )
  );
  al_and2 _09594_ (
    .a(RESET),
    .b(\DFF_1277.Q ),
    .y(\DFF_1309.D )
  );
  al_and2 _09595_ (
    .a(RESET),
    .b(\DFF_1278.Q ),
    .y(\DFF_1310.D )
  );
  al_and2 _09596_ (
    .a(RESET),
    .b(\DFF_1279.Q ),
    .y(\DFF_1311.D )
  );
  al_oa21ftt _09597_ (
    .a(\DFF_1311.Q ),
    .b(\DFF_1343.Q ),
    .c(RESET),
    .y(_03801_)
  );
  al_aoi21ftf _09598_ (
    .a(\DFF_1311.Q ),
    .b(\DFF_1343.Q ),
    .c(_03801_),
    .y(\DFF_1312.D )
  );
  al_oa21ftt _09599_ (
    .a(\DFF_1310.Q ),
    .b(\DFF_1312.Q ),
    .c(RESET),
    .y(_03802_)
  );
  al_aoi21ftf _09600_ (
    .a(\DFF_1310.Q ),
    .b(\DFF_1312.Q ),
    .c(_03802_),
    .y(\DFF_1313.D )
  );
  al_oa21ftt _09601_ (
    .a(\DFF_1309.Q ),
    .b(\DFF_1313.Q ),
    .c(RESET),
    .y(_03803_)
  );
  al_aoi21ftf _09602_ (
    .a(\DFF_1309.Q ),
    .b(\DFF_1313.Q ),
    .c(_03803_),
    .y(\DFF_1314.D )
  );
  al_oa21ftt _09603_ (
    .a(\DFF_1308.Q ),
    .b(\DFF_1314.Q ),
    .c(RESET),
    .y(_03804_)
  );
  al_aoi21ftf _09604_ (
    .a(\DFF_1308.Q ),
    .b(\DFF_1314.Q ),
    .c(_03804_),
    .y(\DFF_1315.D )
  );
  al_nand2ft _09605_ (
    .a(\DFF_1307.Q ),
    .b(\DFF_1315.Q ),
    .y(_03805_)
  );
  al_nand2ft _09606_ (
    .a(\DFF_1315.Q ),
    .b(\DFF_1307.Q ),
    .y(_03806_)
  );
  al_ao21ttf _09607_ (
    .a(_03805_),
    .b(_03806_),
    .c(\DFF_1343.Q ),
    .y(_03807_)
  );
  al_nand3ftt _09608_ (
    .a(\DFF_1343.Q ),
    .b(_03805_),
    .c(_03806_),
    .y(_03808_)
  );
  al_aoi21 _09609_ (
    .a(_03808_),
    .b(_03807_),
    .c(_00451_),
    .y(\DFF_1316.D )
  );
  al_oa21ftt _09610_ (
    .a(\DFF_1306.Q ),
    .b(\DFF_1316.Q ),
    .c(RESET),
    .y(_03809_)
  );
  al_aoi21ftf _09611_ (
    .a(\DFF_1306.Q ),
    .b(\DFF_1316.Q ),
    .c(_03809_),
    .y(\DFF_1317.D )
  );
  al_oa21ftt _09612_ (
    .a(\DFF_1305.Q ),
    .b(\DFF_1317.Q ),
    .c(RESET),
    .y(_03810_)
  );
  al_aoi21ftf _09613_ (
    .a(\DFF_1305.Q ),
    .b(\DFF_1317.Q ),
    .c(_03810_),
    .y(\DFF_1318.D )
  );
  al_oa21ftt _09614_ (
    .a(\DFF_1304.Q ),
    .b(\DFF_1318.Q ),
    .c(RESET),
    .y(_03811_)
  );
  al_aoi21ftf _09615_ (
    .a(\DFF_1304.Q ),
    .b(\DFF_1318.Q ),
    .c(_03811_),
    .y(\DFF_1319.D )
  );
  al_oa21ftt _09616_ (
    .a(\DFF_1303.Q ),
    .b(\DFF_1319.Q ),
    .c(RESET),
    .y(_03812_)
  );
  al_aoi21ftf _09617_ (
    .a(\DFF_1303.Q ),
    .b(\DFF_1319.Q ),
    .c(_03812_),
    .y(\DFF_1320.D )
  );
  al_oa21ftt _09618_ (
    .a(\DFF_1302.Q ),
    .b(\DFF_1320.Q ),
    .c(RESET),
    .y(_03813_)
  );
  al_aoi21ftf _09619_ (
    .a(\DFF_1302.Q ),
    .b(\DFF_1320.Q ),
    .c(_03813_),
    .y(\DFF_1321.D )
  );
  al_oa21ftt _09620_ (
    .a(\DFF_1301.Q ),
    .b(\DFF_1321.Q ),
    .c(RESET),
    .y(_03814_)
  );
  al_aoi21ftf _09621_ (
    .a(\DFF_1301.Q ),
    .b(\DFF_1321.Q ),
    .c(_03814_),
    .y(\DFF_1322.D )
  );
  al_nand2ft _09622_ (
    .a(\DFF_1300.Q ),
    .b(\DFF_1322.Q ),
    .y(_03815_)
  );
  al_nand2ft _09623_ (
    .a(\DFF_1322.Q ),
    .b(\DFF_1300.Q ),
    .y(_03816_)
  );
  al_ao21ttf _09624_ (
    .a(_03815_),
    .b(_03816_),
    .c(\DFF_1343.Q ),
    .y(_03817_)
  );
  al_nand3ftt _09625_ (
    .a(\DFF_1343.Q ),
    .b(_03815_),
    .c(_03816_),
    .y(_03818_)
  );
  al_aoi21 _09626_ (
    .a(_03818_),
    .b(_03817_),
    .c(_00451_),
    .y(\DFF_1323.D )
  );
  al_oa21ftt _09627_ (
    .a(\DFF_1299.Q ),
    .b(\DFF_1323.Q ),
    .c(RESET),
    .y(_03819_)
  );
  al_aoi21ftf _09628_ (
    .a(\DFF_1299.Q ),
    .b(\DFF_1323.Q ),
    .c(_03819_),
    .y(\DFF_1324.D )
  );
  al_oa21ftt _09629_ (
    .a(\DFF_1298.Q ),
    .b(\DFF_1324.Q ),
    .c(RESET),
    .y(_03820_)
  );
  al_aoi21ftf _09630_ (
    .a(\DFF_1298.Q ),
    .b(\DFF_1324.Q ),
    .c(_03820_),
    .y(\DFF_1325.D )
  );
  al_oa21ftt _09631_ (
    .a(\DFF_1297.Q ),
    .b(\DFF_1325.Q ),
    .c(RESET),
    .y(_03821_)
  );
  al_aoi21ftf _09632_ (
    .a(\DFF_1297.Q ),
    .b(\DFF_1325.Q ),
    .c(_03821_),
    .y(\DFF_1326.D )
  );
  al_oa21ftt _09633_ (
    .a(\DFF_1296.Q ),
    .b(\DFF_1326.Q ),
    .c(RESET),
    .y(_03822_)
  );
  al_aoi21ftf _09634_ (
    .a(\DFF_1296.Q ),
    .b(\DFF_1326.Q ),
    .c(_03822_),
    .y(\DFF_1327.D )
  );
  al_nand2ft _09635_ (
    .a(\DFF_1295.Q ),
    .b(\DFF_1327.Q ),
    .y(_03823_)
  );
  al_nand2ft _09636_ (
    .a(\DFF_1327.Q ),
    .b(\DFF_1295.Q ),
    .y(_03824_)
  );
  al_ao21ttf _09637_ (
    .a(_03823_),
    .b(_03824_),
    .c(\DFF_1343.Q ),
    .y(_03825_)
  );
  al_nand3ftt _09638_ (
    .a(\DFF_1343.Q ),
    .b(_03823_),
    .c(_03824_),
    .y(_03826_)
  );
  al_aoi21 _09639_ (
    .a(_03826_),
    .b(_03825_),
    .c(_00451_),
    .y(\DFF_1328.D )
  );
  al_oa21ftt _09640_ (
    .a(\DFF_1294.Q ),
    .b(\DFF_1328.Q ),
    .c(RESET),
    .y(_03827_)
  );
  al_aoi21ftf _09641_ (
    .a(\DFF_1294.Q ),
    .b(\DFF_1328.Q ),
    .c(_03827_),
    .y(\DFF_1329.D )
  );
  al_oa21ftt _09642_ (
    .a(\DFF_1293.Q ),
    .b(\DFF_1329.Q ),
    .c(RESET),
    .y(_03828_)
  );
  al_aoi21ftf _09643_ (
    .a(\DFF_1293.Q ),
    .b(\DFF_1329.Q ),
    .c(_03828_),
    .y(\DFF_1330.D )
  );
  al_oa21ftt _09644_ (
    .a(\DFF_1292.Q ),
    .b(\DFF_1330.Q ),
    .c(RESET),
    .y(_03829_)
  );
  al_aoi21ftf _09645_ (
    .a(\DFF_1292.Q ),
    .b(\DFF_1330.Q ),
    .c(_03829_),
    .y(\DFF_1331.D )
  );
  al_oa21ftt _09646_ (
    .a(\DFF_1291.Q ),
    .b(\DFF_1331.Q ),
    .c(RESET),
    .y(_03830_)
  );
  al_aoi21ftf _09647_ (
    .a(\DFF_1291.Q ),
    .b(\DFF_1331.Q ),
    .c(_03830_),
    .y(\DFF_1332.D )
  );
  al_oa21ftt _09648_ (
    .a(\DFF_1290.Q ),
    .b(\DFF_1332.Q ),
    .c(RESET),
    .y(_03831_)
  );
  al_aoi21ftf _09649_ (
    .a(\DFF_1290.Q ),
    .b(\DFF_1332.Q ),
    .c(_03831_),
    .y(\DFF_1333.D )
  );
  al_oa21ftt _09650_ (
    .a(\DFF_1289.Q ),
    .b(\DFF_1333.Q ),
    .c(RESET),
    .y(_03832_)
  );
  al_aoi21ftf _09651_ (
    .a(\DFF_1289.Q ),
    .b(\DFF_1333.Q ),
    .c(_03832_),
    .y(\DFF_1334.D )
  );
  al_oa21ftt _09652_ (
    .a(\DFF_1288.Q ),
    .b(\DFF_1334.Q ),
    .c(RESET),
    .y(_03833_)
  );
  al_aoi21ftf _09653_ (
    .a(\DFF_1288.Q ),
    .b(\DFF_1334.Q ),
    .c(_03833_),
    .y(\DFF_1335.D )
  );
  al_oa21ftt _09654_ (
    .a(\DFF_1287.Q ),
    .b(\DFF_1335.Q ),
    .c(RESET),
    .y(_03834_)
  );
  al_aoi21ftf _09655_ (
    .a(\DFF_1287.Q ),
    .b(\DFF_1335.Q ),
    .c(_03834_),
    .y(\DFF_1336.D )
  );
  al_oa21ftt _09656_ (
    .a(\DFF_1286.Q ),
    .b(\DFF_1336.Q ),
    .c(RESET),
    .y(_03835_)
  );
  al_aoi21ftf _09657_ (
    .a(\DFF_1286.Q ),
    .b(\DFF_1336.Q ),
    .c(_03835_),
    .y(\DFF_1337.D )
  );
  al_oa21ftt _09658_ (
    .a(\DFF_1285.Q ),
    .b(\DFF_1337.Q ),
    .c(RESET),
    .y(_03836_)
  );
  al_aoi21ftf _09659_ (
    .a(\DFF_1285.Q ),
    .b(\DFF_1337.Q ),
    .c(_03836_),
    .y(\DFF_1338.D )
  );
  al_oa21ftt _09660_ (
    .a(\DFF_1284.Q ),
    .b(\DFF_1338.Q ),
    .c(RESET),
    .y(_03837_)
  );
  al_aoi21ftf _09661_ (
    .a(\DFF_1284.Q ),
    .b(\DFF_1338.Q ),
    .c(_03837_),
    .y(\DFF_1339.D )
  );
  al_oa21ftt _09662_ (
    .a(\DFF_1283.Q ),
    .b(\DFF_1339.Q ),
    .c(RESET),
    .y(_03838_)
  );
  al_aoi21ftf _09663_ (
    .a(\DFF_1283.Q ),
    .b(\DFF_1339.Q ),
    .c(_03838_),
    .y(\DFF_1340.D )
  );
  al_oa21ftt _09664_ (
    .a(\DFF_1282.Q ),
    .b(\DFF_1340.Q ),
    .c(RESET),
    .y(_03839_)
  );
  al_aoi21ftf _09665_ (
    .a(\DFF_1282.Q ),
    .b(\DFF_1340.Q ),
    .c(_03839_),
    .y(\DFF_1341.D )
  );
  al_oa21ftt _09666_ (
    .a(\DFF_1281.Q ),
    .b(\DFF_1341.Q ),
    .c(RESET),
    .y(_03840_)
  );
  al_aoi21ftf _09667_ (
    .a(\DFF_1281.Q ),
    .b(\DFF_1341.Q ),
    .c(_03840_),
    .y(\DFF_1342.D )
  );
  al_oa21ftt _09668_ (
    .a(\DFF_1280.Q ),
    .b(\DFF_1342.Q ),
    .c(RESET),
    .y(_03841_)
  );
  al_aoi21ftf _09669_ (
    .a(\DFF_1280.Q ),
    .b(\DFF_1342.Q ),
    .c(_03841_),
    .y(\DFF_1343.D )
  );
  al_and2 _09670_ (
    .a(RESET),
    .b(\DFF_1345.Q ),
    .y(\DFF_1344.D )
  );
  al_and2 _09671_ (
    .a(RESET),
    .b(\DFF_1346.Q ),
    .y(\DFF_1345.D )
  );
  al_and2 _09672_ (
    .a(RESET),
    .b(\DFF_1347.Q ),
    .y(\DFF_1346.D )
  );
  al_and2 _09673_ (
    .a(RESET),
    .b(\DFF_1348.Q ),
    .y(\DFF_1347.D )
  );
  al_and2 _09674_ (
    .a(RESET),
    .b(\DFF_1349.Q ),
    .y(\DFF_1348.D )
  );
  al_and2 _09675_ (
    .a(RESET),
    .b(\DFF_1350.Q ),
    .y(\DFF_1349.D )
  );
  al_and2 _09676_ (
    .a(RESET),
    .b(\DFF_1351.Q ),
    .y(\DFF_1350.D )
  );
  al_and2 _09677_ (
    .a(RESET),
    .b(\DFF_1352.Q ),
    .y(\DFF_1351.D )
  );
  al_and2 _09678_ (
    .a(RESET),
    .b(\DFF_1353.Q ),
    .y(\DFF_1352.D )
  );
  al_and2 _09679_ (
    .a(RESET),
    .b(\DFF_1354.Q ),
    .y(\DFF_1353.D )
  );
  al_and2 _09680_ (
    .a(RESET),
    .b(\DFF_1355.Q ),
    .y(\DFF_1354.D )
  );
  al_and2 _09681_ (
    .a(RESET),
    .b(\DFF_1356.Q ),
    .y(\DFF_1355.D )
  );
  al_and2 _09682_ (
    .a(RESET),
    .b(\DFF_1357.Q ),
    .y(\DFF_1356.D )
  );
  al_and2 _09683_ (
    .a(RESET),
    .b(\DFF_1358.Q ),
    .y(\DFF_1357.D )
  );
  al_and2 _09684_ (
    .a(RESET),
    .b(\DFF_1359.Q ),
    .y(\DFF_1358.D )
  );
  al_and2 _09685_ (
    .a(RESET),
    .b(\DFF_1360.Q ),
    .y(\DFF_1359.D )
  );
  al_and2 _09686_ (
    .a(RESET),
    .b(\DFF_1361.Q ),
    .y(\DFF_1360.D )
  );
  al_and2 _09687_ (
    .a(RESET),
    .b(\DFF_1362.Q ),
    .y(\DFF_1361.D )
  );
  al_and2 _09688_ (
    .a(RESET),
    .b(\DFF_1363.Q ),
    .y(\DFF_1362.D )
  );
  al_and2 _09689_ (
    .a(RESET),
    .b(\DFF_1364.Q ),
    .y(\DFF_1363.D )
  );
  al_and2 _09690_ (
    .a(RESET),
    .b(\DFF_1365.Q ),
    .y(\DFF_1364.D )
  );
  al_and2 _09691_ (
    .a(RESET),
    .b(\DFF_1366.Q ),
    .y(\DFF_1365.D )
  );
  al_and2 _09692_ (
    .a(RESET),
    .b(\DFF_1367.Q ),
    .y(\DFF_1366.D )
  );
  al_and2 _09693_ (
    .a(RESET),
    .b(\DFF_1368.Q ),
    .y(\DFF_1367.D )
  );
  al_and2 _09694_ (
    .a(RESET),
    .b(\DFF_1369.Q ),
    .y(\DFF_1368.D )
  );
  al_and2 _09695_ (
    .a(RESET),
    .b(\DFF_1370.Q ),
    .y(\DFF_1369.D )
  );
  al_and2 _09696_ (
    .a(RESET),
    .b(\DFF_1371.Q ),
    .y(\DFF_1370.D )
  );
  al_and2 _09697_ (
    .a(RESET),
    .b(\DFF_1372.Q ),
    .y(\DFF_1371.D )
  );
  al_and2 _09698_ (
    .a(RESET),
    .b(\DFF_1373.Q ),
    .y(\DFF_1372.D )
  );
  al_and2 _09699_ (
    .a(RESET),
    .b(\DFF_1374.Q ),
    .y(\DFF_1373.D )
  );
  al_and2 _09700_ (
    .a(RESET),
    .b(\DFF_1375.Q ),
    .y(\DFF_1374.D )
  );
  al_and2ft _09701_ (
    .a(\DFF_1344.Q ),
    .b(RESET),
    .y(\DFF_1375.D )
  );
  al_or2 _09702_ (
    .a(TM1),
    .b(\DFF_1632.Q ),
    .y(_03842_)
  );
  al_nand2 _09703_ (
    .a(TM1),
    .b(\DFF_1632.Q ),
    .y(_03843_)
  );
  al_nand3 _09704_ (
    .a(\DFF_1664.Q ),
    .b(_03842_),
    .c(_03843_),
    .y(_03844_)
  );
  al_nand2ft _09705_ (
    .a(TM1),
    .b(\DFF_1632.Q ),
    .y(_03845_)
  );
  al_and2ft _09706_ (
    .a(\DFF_1632.Q ),
    .b(TM1),
    .y(_03846_)
  );
  al_and3fft _09707_ (
    .a(\DFF_1664.Q ),
    .b(_03846_),
    .c(_03845_),
    .y(_03847_)
  );
  al_and2ft _09708_ (
    .a(\DFF_1600.Q ),
    .b(\DFF_1568.Q ),
    .y(_03848_)
  );
  al_nand2ft _09709_ (
    .a(\DFF_1568.Q ),
    .b(\DFF_1600.Q ),
    .y(_03849_)
  );
  al_nand2ft _09710_ (
    .a(_03848_),
    .b(_03849_),
    .y(_03850_)
  );
  al_oai21ftf _09711_ (
    .a(_03844_),
    .b(_03847_),
    .c(_03850_),
    .y(_03851_)
  );
  al_nand3ftt _09712_ (
    .a(_03847_),
    .b(_03844_),
    .c(_03850_),
    .y(_03852_)
  );
  al_nand3 _09713_ (
    .a(_00448_),
    .b(_03851_),
    .c(_03852_),
    .y(_03853_)
  );
  al_aoi21 _09714_ (
    .a(TM0),
    .b(\DFF_1535.Q ),
    .c(TM1),
    .y(_03854_)
  );
  al_nand2 _09715_ (
    .a(_03854_),
    .b(_03853_),
    .y(_03855_)
  );
  al_aoi21ttf _09716_ (
    .a(\DFF_1344.Q ),
    .b(TM0),
    .c(TM1),
    .y(_03856_)
  );
  al_and2 _09717_ (
    .a(_03856_),
    .b(_03364_),
    .y(_03857_)
  );
  al_nor3fft _09718_ (
    .a(RESET),
    .b(_03855_),
    .c(_03857_),
    .y(\DFF_1376.D )
  );
  al_or2 _09719_ (
    .a(TM1),
    .b(\DFF_1633.Q ),
    .y(_03858_)
  );
  al_nand2 _09720_ (
    .a(TM1),
    .b(\DFF_1633.Q ),
    .y(_03859_)
  );
  al_nand3 _09721_ (
    .a(\DFF_1665.Q ),
    .b(_03858_),
    .c(_03859_),
    .y(_03860_)
  );
  al_nand2ft _09722_ (
    .a(TM1),
    .b(\DFF_1633.Q ),
    .y(_03861_)
  );
  al_and2ft _09723_ (
    .a(\DFF_1633.Q ),
    .b(TM1),
    .y(_03862_)
  );
  al_and3fft _09724_ (
    .a(\DFF_1665.Q ),
    .b(_03862_),
    .c(_03861_),
    .y(_03863_)
  );
  al_and2ft _09725_ (
    .a(\DFF_1601.Q ),
    .b(\DFF_1569.Q ),
    .y(_03864_)
  );
  al_nand2ft _09726_ (
    .a(\DFF_1569.Q ),
    .b(\DFF_1601.Q ),
    .y(_03865_)
  );
  al_nand2ft _09727_ (
    .a(_03864_),
    .b(_03865_),
    .y(_03866_)
  );
  al_oai21ftf _09728_ (
    .a(_03860_),
    .b(_03863_),
    .c(_03866_),
    .y(_03867_)
  );
  al_nand3ftt _09729_ (
    .a(_03863_),
    .b(_03860_),
    .c(_03866_),
    .y(_03868_)
  );
  al_nand3 _09730_ (
    .a(_00448_),
    .b(_03867_),
    .c(_03868_),
    .y(_03869_)
  );
  al_aoi21 _09731_ (
    .a(TM0),
    .b(\DFF_1534.Q ),
    .c(TM1),
    .y(_03870_)
  );
  al_nand2 _09732_ (
    .a(_03870_),
    .b(_03869_),
    .y(_03871_)
  );
  al_aoi21ttf _09733_ (
    .a(TM0),
    .b(\DFF_1345.Q ),
    .c(TM1),
    .y(_03872_)
  );
  al_and2 _09734_ (
    .a(_03872_),
    .b(_03380_),
    .y(_03873_)
  );
  al_nor3fft _09735_ (
    .a(RESET),
    .b(_03871_),
    .c(_03873_),
    .y(\DFF_1377.D )
  );
  al_or2 _09736_ (
    .a(TM1),
    .b(\DFF_1634.Q ),
    .y(_03874_)
  );
  al_nand2 _09737_ (
    .a(TM1),
    .b(\DFF_1634.Q ),
    .y(_03875_)
  );
  al_nand3 _09738_ (
    .a(\DFF_1666.Q ),
    .b(_03874_),
    .c(_03875_),
    .y(_03876_)
  );
  al_nand2ft _09739_ (
    .a(TM1),
    .b(\DFF_1634.Q ),
    .y(_03877_)
  );
  al_and2ft _09740_ (
    .a(\DFF_1634.Q ),
    .b(TM1),
    .y(_03878_)
  );
  al_and3fft _09741_ (
    .a(\DFF_1666.Q ),
    .b(_03878_),
    .c(_03877_),
    .y(_03879_)
  );
  al_and2ft _09742_ (
    .a(\DFF_1602.Q ),
    .b(\DFF_1570.Q ),
    .y(_03880_)
  );
  al_nand2ft _09743_ (
    .a(\DFF_1570.Q ),
    .b(\DFF_1602.Q ),
    .y(_03881_)
  );
  al_nand2ft _09744_ (
    .a(_03880_),
    .b(_03881_),
    .y(_03882_)
  );
  al_oai21ftf _09745_ (
    .a(_03876_),
    .b(_03879_),
    .c(_03882_),
    .y(_03883_)
  );
  al_nand3ftt _09746_ (
    .a(_03879_),
    .b(_03876_),
    .c(_03882_),
    .y(_03884_)
  );
  al_nand3 _09747_ (
    .a(_00448_),
    .b(_03883_),
    .c(_03884_),
    .y(_03885_)
  );
  al_aoi21 _09748_ (
    .a(TM0),
    .b(\DFF_1533.Q ),
    .c(TM1),
    .y(_03886_)
  );
  al_nand2 _09749_ (
    .a(_03886_),
    .b(_03885_),
    .y(_03887_)
  );
  al_aoi21ttf _09750_ (
    .a(TM0),
    .b(\DFF_1346.Q ),
    .c(TM1),
    .y(_03888_)
  );
  al_and2 _09751_ (
    .a(_03888_),
    .b(_03396_),
    .y(_03889_)
  );
  al_nor3fft _09752_ (
    .a(RESET),
    .b(_03887_),
    .c(_03889_),
    .y(\DFF_1378.D )
  );
  al_or2 _09753_ (
    .a(TM1),
    .b(\DFF_1635.Q ),
    .y(_03890_)
  );
  al_nand2 _09754_ (
    .a(TM1),
    .b(\DFF_1635.Q ),
    .y(_03891_)
  );
  al_nand3 _09755_ (
    .a(\DFF_1667.Q ),
    .b(_03890_),
    .c(_03891_),
    .y(_03892_)
  );
  al_nand2ft _09756_ (
    .a(TM1),
    .b(\DFF_1635.Q ),
    .y(_03893_)
  );
  al_and2ft _09757_ (
    .a(\DFF_1635.Q ),
    .b(TM1),
    .y(_03894_)
  );
  al_and3fft _09758_ (
    .a(\DFF_1667.Q ),
    .b(_03894_),
    .c(_03893_),
    .y(_03895_)
  );
  al_and2ft _09759_ (
    .a(\DFF_1603.Q ),
    .b(\DFF_1571.Q ),
    .y(_03896_)
  );
  al_nand2ft _09760_ (
    .a(\DFF_1571.Q ),
    .b(\DFF_1603.Q ),
    .y(_03897_)
  );
  al_nand2ft _09761_ (
    .a(_03896_),
    .b(_03897_),
    .y(_03898_)
  );
  al_oai21ftf _09762_ (
    .a(_03892_),
    .b(_03895_),
    .c(_03898_),
    .y(_03899_)
  );
  al_nand3ftt _09763_ (
    .a(_03895_),
    .b(_03892_),
    .c(_03898_),
    .y(_03900_)
  );
  al_nand3 _09764_ (
    .a(_00448_),
    .b(_03899_),
    .c(_03900_),
    .y(_03901_)
  );
  al_aoi21 _09765_ (
    .a(TM0),
    .b(\DFF_1532.Q ),
    .c(TM1),
    .y(_03902_)
  );
  al_nand2 _09766_ (
    .a(_03902_),
    .b(_03901_),
    .y(_03903_)
  );
  al_aoi21ttf _09767_ (
    .a(TM0),
    .b(\DFF_1347.Q ),
    .c(TM1),
    .y(_03904_)
  );
  al_and2 _09768_ (
    .a(_03904_),
    .b(_03412_),
    .y(_03905_)
  );
  al_nor3fft _09769_ (
    .a(RESET),
    .b(_03903_),
    .c(_03905_),
    .y(\DFF_1379.D )
  );
  al_or2 _09770_ (
    .a(TM1),
    .b(\DFF_1636.Q ),
    .y(_03906_)
  );
  al_nand2 _09771_ (
    .a(TM1),
    .b(\DFF_1636.Q ),
    .y(_03907_)
  );
  al_nand3 _09772_ (
    .a(\DFF_1668.Q ),
    .b(_03906_),
    .c(_03907_),
    .y(_03908_)
  );
  al_nand2ft _09773_ (
    .a(TM1),
    .b(\DFF_1636.Q ),
    .y(_03909_)
  );
  al_and2ft _09774_ (
    .a(\DFF_1636.Q ),
    .b(TM1),
    .y(_03910_)
  );
  al_and3fft _09775_ (
    .a(\DFF_1668.Q ),
    .b(_03910_),
    .c(_03909_),
    .y(_03911_)
  );
  al_and2ft _09776_ (
    .a(\DFF_1604.Q ),
    .b(\DFF_1572.Q ),
    .y(_03912_)
  );
  al_nand2ft _09777_ (
    .a(\DFF_1572.Q ),
    .b(\DFF_1604.Q ),
    .y(_03913_)
  );
  al_nand2ft _09778_ (
    .a(_03912_),
    .b(_03913_),
    .y(_03914_)
  );
  al_oai21ftf _09779_ (
    .a(_03908_),
    .b(_03911_),
    .c(_03914_),
    .y(_03915_)
  );
  al_nand3ftt _09780_ (
    .a(_03911_),
    .b(_03908_),
    .c(_03914_),
    .y(_03916_)
  );
  al_nand3 _09781_ (
    .a(_00448_),
    .b(_03915_),
    .c(_03916_),
    .y(_03917_)
  );
  al_aoi21 _09782_ (
    .a(TM0),
    .b(\DFF_1531.Q ),
    .c(TM1),
    .y(_03918_)
  );
  al_nand2 _09783_ (
    .a(_03918_),
    .b(_03917_),
    .y(_03919_)
  );
  al_aoi21ttf _09784_ (
    .a(TM0),
    .b(\DFF_1348.Q ),
    .c(TM1),
    .y(_03920_)
  );
  al_and2 _09785_ (
    .a(_03920_),
    .b(_03428_),
    .y(_03921_)
  );
  al_nor3fft _09786_ (
    .a(RESET),
    .b(_03919_),
    .c(_03921_),
    .y(\DFF_1380.D )
  );
  al_or2 _09787_ (
    .a(TM1),
    .b(\DFF_1637.Q ),
    .y(_03922_)
  );
  al_nand2 _09788_ (
    .a(TM1),
    .b(\DFF_1637.Q ),
    .y(_03923_)
  );
  al_nand3 _09789_ (
    .a(\DFF_1669.Q ),
    .b(_03922_),
    .c(_03923_),
    .y(_03924_)
  );
  al_nand2ft _09790_ (
    .a(TM1),
    .b(\DFF_1637.Q ),
    .y(_03925_)
  );
  al_and2ft _09791_ (
    .a(\DFF_1637.Q ),
    .b(TM1),
    .y(_03926_)
  );
  al_and3fft _09792_ (
    .a(\DFF_1669.Q ),
    .b(_03926_),
    .c(_03925_),
    .y(_03927_)
  );
  al_and2ft _09793_ (
    .a(\DFF_1605.Q ),
    .b(\DFF_1573.Q ),
    .y(_03928_)
  );
  al_nand2ft _09794_ (
    .a(\DFF_1573.Q ),
    .b(\DFF_1605.Q ),
    .y(_03929_)
  );
  al_nand2ft _09795_ (
    .a(_03928_),
    .b(_03929_),
    .y(_03930_)
  );
  al_oai21ftf _09796_ (
    .a(_03924_),
    .b(_03927_),
    .c(_03930_),
    .y(_03931_)
  );
  al_nand3ftt _09797_ (
    .a(_03927_),
    .b(_03924_),
    .c(_03930_),
    .y(_03932_)
  );
  al_nand3 _09798_ (
    .a(_00448_),
    .b(_03931_),
    .c(_03932_),
    .y(_03933_)
  );
  al_aoi21 _09799_ (
    .a(TM0),
    .b(\DFF_1530.Q ),
    .c(TM1),
    .y(_03934_)
  );
  al_nand2 _09800_ (
    .a(_03934_),
    .b(_03933_),
    .y(_03935_)
  );
  al_aoi21ttf _09801_ (
    .a(TM0),
    .b(\DFF_1349.Q ),
    .c(TM1),
    .y(_03936_)
  );
  al_and2 _09802_ (
    .a(_03936_),
    .b(_03444_),
    .y(_03937_)
  );
  al_nor3fft _09803_ (
    .a(RESET),
    .b(_03935_),
    .c(_03937_),
    .y(\DFF_1381.D )
  );
  al_or2 _09804_ (
    .a(TM1),
    .b(\DFF_1638.Q ),
    .y(_03938_)
  );
  al_nand2 _09805_ (
    .a(TM1),
    .b(\DFF_1638.Q ),
    .y(_03939_)
  );
  al_nand3 _09806_ (
    .a(\DFF_1670.Q ),
    .b(_03938_),
    .c(_03939_),
    .y(_03940_)
  );
  al_nand2ft _09807_ (
    .a(TM1),
    .b(\DFF_1638.Q ),
    .y(_03941_)
  );
  al_and2ft _09808_ (
    .a(\DFF_1638.Q ),
    .b(TM1),
    .y(_03942_)
  );
  al_and3fft _09809_ (
    .a(\DFF_1670.Q ),
    .b(_03942_),
    .c(_03941_),
    .y(_03943_)
  );
  al_and2ft _09810_ (
    .a(\DFF_1606.Q ),
    .b(\DFF_1574.Q ),
    .y(_03944_)
  );
  al_nand2ft _09811_ (
    .a(\DFF_1574.Q ),
    .b(\DFF_1606.Q ),
    .y(_03945_)
  );
  al_nand2ft _09812_ (
    .a(_03944_),
    .b(_03945_),
    .y(_03946_)
  );
  al_oai21ftf _09813_ (
    .a(_03940_),
    .b(_03943_),
    .c(_03946_),
    .y(_03947_)
  );
  al_nand3ftt _09814_ (
    .a(_03943_),
    .b(_03940_),
    .c(_03946_),
    .y(_03948_)
  );
  al_nand3 _09815_ (
    .a(_00448_),
    .b(_03947_),
    .c(_03948_),
    .y(_03949_)
  );
  al_aoi21 _09816_ (
    .a(TM0),
    .b(\DFF_1529.Q ),
    .c(TM1),
    .y(_03950_)
  );
  al_nand2 _09817_ (
    .a(_03950_),
    .b(_03949_),
    .y(_03951_)
  );
  al_aoi21ttf _09818_ (
    .a(TM0),
    .b(\DFF_1350.Q ),
    .c(TM1),
    .y(_03952_)
  );
  al_and2 _09819_ (
    .a(_03952_),
    .b(_03460_),
    .y(_03953_)
  );
  al_nor3fft _09820_ (
    .a(RESET),
    .b(_03951_),
    .c(_03953_),
    .y(\DFF_1382.D )
  );
  al_or2 _09821_ (
    .a(TM1),
    .b(\DFF_1639.Q ),
    .y(_03954_)
  );
  al_nand2 _09822_ (
    .a(TM1),
    .b(\DFF_1639.Q ),
    .y(_03955_)
  );
  al_nand3 _09823_ (
    .a(\DFF_1671.Q ),
    .b(_03954_),
    .c(_03955_),
    .y(_03956_)
  );
  al_nand2ft _09824_ (
    .a(TM1),
    .b(\DFF_1639.Q ),
    .y(_03957_)
  );
  al_and2ft _09825_ (
    .a(\DFF_1639.Q ),
    .b(TM1),
    .y(_03958_)
  );
  al_and3fft _09826_ (
    .a(\DFF_1671.Q ),
    .b(_03958_),
    .c(_03957_),
    .y(_03959_)
  );
  al_and2ft _09827_ (
    .a(\DFF_1607.Q ),
    .b(\DFF_1575.Q ),
    .y(_03960_)
  );
  al_nand2ft _09828_ (
    .a(\DFF_1575.Q ),
    .b(\DFF_1607.Q ),
    .y(_03961_)
  );
  al_nand2ft _09829_ (
    .a(_03960_),
    .b(_03961_),
    .y(_03962_)
  );
  al_oai21ftf _09830_ (
    .a(_03956_),
    .b(_03959_),
    .c(_03962_),
    .y(_03963_)
  );
  al_nand3ftt _09831_ (
    .a(_03959_),
    .b(_03956_),
    .c(_03962_),
    .y(_03964_)
  );
  al_nand3 _09832_ (
    .a(_00448_),
    .b(_03963_),
    .c(_03964_),
    .y(_03965_)
  );
  al_aoi21 _09833_ (
    .a(TM0),
    .b(\DFF_1528.Q ),
    .c(TM1),
    .y(_03966_)
  );
  al_nand2 _09834_ (
    .a(_03966_),
    .b(_03965_),
    .y(_03967_)
  );
  al_aoi21ttf _09835_ (
    .a(TM0),
    .b(\DFF_1351.Q ),
    .c(TM1),
    .y(_03968_)
  );
  al_and2 _09836_ (
    .a(_03968_),
    .b(_03476_),
    .y(_03969_)
  );
  al_nor3fft _09837_ (
    .a(RESET),
    .b(_03967_),
    .c(_03969_),
    .y(\DFF_1383.D )
  );
  al_or2 _09838_ (
    .a(TM1),
    .b(\DFF_1640.Q ),
    .y(_03970_)
  );
  al_nand2 _09839_ (
    .a(TM1),
    .b(\DFF_1640.Q ),
    .y(_03971_)
  );
  al_nand3 _09840_ (
    .a(\DFF_1672.Q ),
    .b(_03970_),
    .c(_03971_),
    .y(_03972_)
  );
  al_nand2ft _09841_ (
    .a(TM1),
    .b(\DFF_1640.Q ),
    .y(_03973_)
  );
  al_and2ft _09842_ (
    .a(\DFF_1640.Q ),
    .b(TM1),
    .y(_03974_)
  );
  al_and3fft _09843_ (
    .a(\DFF_1672.Q ),
    .b(_03974_),
    .c(_03973_),
    .y(_03975_)
  );
  al_and2ft _09844_ (
    .a(\DFF_1608.Q ),
    .b(\DFF_1576.Q ),
    .y(_03976_)
  );
  al_nand2ft _09845_ (
    .a(\DFF_1576.Q ),
    .b(\DFF_1608.Q ),
    .y(_03977_)
  );
  al_nand2ft _09846_ (
    .a(_03976_),
    .b(_03977_),
    .y(_03978_)
  );
  al_oai21ftf _09847_ (
    .a(_03972_),
    .b(_03975_),
    .c(_03978_),
    .y(_03979_)
  );
  al_nand3ftt _09848_ (
    .a(_03975_),
    .b(_03972_),
    .c(_03978_),
    .y(_03980_)
  );
  al_nand3 _09849_ (
    .a(_00448_),
    .b(_03979_),
    .c(_03980_),
    .y(_03981_)
  );
  al_aoi21 _09850_ (
    .a(TM0),
    .b(\DFF_1527.Q ),
    .c(TM1),
    .y(_03982_)
  );
  al_nand2 _09851_ (
    .a(_03982_),
    .b(_03981_),
    .y(_03983_)
  );
  al_aoi21ttf _09852_ (
    .a(TM0),
    .b(\DFF_1352.Q ),
    .c(TM1),
    .y(_03984_)
  );
  al_and2 _09853_ (
    .a(_03984_),
    .b(_03492_),
    .y(_03985_)
  );
  al_nor3fft _09854_ (
    .a(RESET),
    .b(_03983_),
    .c(_03985_),
    .y(\DFF_1384.D )
  );
  al_or2 _09855_ (
    .a(TM1),
    .b(\DFF_1641.Q ),
    .y(_03986_)
  );
  al_nand2 _09856_ (
    .a(TM1),
    .b(\DFF_1641.Q ),
    .y(_03987_)
  );
  al_nand3 _09857_ (
    .a(\DFF_1673.Q ),
    .b(_03986_),
    .c(_03987_),
    .y(_03988_)
  );
  al_nand2ft _09858_ (
    .a(TM1),
    .b(\DFF_1641.Q ),
    .y(_03989_)
  );
  al_and2ft _09859_ (
    .a(\DFF_1641.Q ),
    .b(TM1),
    .y(_03990_)
  );
  al_and3fft _09860_ (
    .a(\DFF_1673.Q ),
    .b(_03990_),
    .c(_03989_),
    .y(_03991_)
  );
  al_and2ft _09861_ (
    .a(\DFF_1609.Q ),
    .b(\DFF_1577.Q ),
    .y(_03992_)
  );
  al_nand2ft _09862_ (
    .a(\DFF_1577.Q ),
    .b(\DFF_1609.Q ),
    .y(_03993_)
  );
  al_nand2ft _09863_ (
    .a(_03992_),
    .b(_03993_),
    .y(_03994_)
  );
  al_oai21ftf _09864_ (
    .a(_03988_),
    .b(_03991_),
    .c(_03994_),
    .y(_03995_)
  );
  al_nand3ftt _09865_ (
    .a(_03991_),
    .b(_03988_),
    .c(_03994_),
    .y(_03996_)
  );
  al_nand3 _09866_ (
    .a(_00448_),
    .b(_03995_),
    .c(_03996_),
    .y(_03997_)
  );
  al_aoi21 _09867_ (
    .a(TM0),
    .b(\DFF_1526.Q ),
    .c(TM1),
    .y(_03998_)
  );
  al_nand2 _09868_ (
    .a(_03998_),
    .b(_03997_),
    .y(_03999_)
  );
  al_aoi21ttf _09869_ (
    .a(TM0),
    .b(\DFF_1353.Q ),
    .c(TM1),
    .y(_04000_)
  );
  al_and2 _09870_ (
    .a(_04000_),
    .b(_03508_),
    .y(_04001_)
  );
  al_nor3fft _09871_ (
    .a(RESET),
    .b(_03999_),
    .c(_04001_),
    .y(\DFF_1385.D )
  );
  al_or2 _09872_ (
    .a(TM1),
    .b(\DFF_1642.Q ),
    .y(_04002_)
  );
  al_nand2 _09873_ (
    .a(TM1),
    .b(\DFF_1642.Q ),
    .y(_04003_)
  );
  al_nand3 _09874_ (
    .a(\DFF_1674.Q ),
    .b(_04002_),
    .c(_04003_),
    .y(_04004_)
  );
  al_nand2ft _09875_ (
    .a(TM1),
    .b(\DFF_1642.Q ),
    .y(_04005_)
  );
  al_and2ft _09876_ (
    .a(\DFF_1642.Q ),
    .b(TM1),
    .y(_04006_)
  );
  al_and3fft _09877_ (
    .a(\DFF_1674.Q ),
    .b(_04006_),
    .c(_04005_),
    .y(_04007_)
  );
  al_and2ft _09878_ (
    .a(\DFF_1610.Q ),
    .b(\DFF_1578.Q ),
    .y(_04008_)
  );
  al_nand2ft _09879_ (
    .a(\DFF_1578.Q ),
    .b(\DFF_1610.Q ),
    .y(_04009_)
  );
  al_nand2ft _09880_ (
    .a(_04008_),
    .b(_04009_),
    .y(_04010_)
  );
  al_oai21ftf _09881_ (
    .a(_04004_),
    .b(_04007_),
    .c(_04010_),
    .y(_04011_)
  );
  al_nand3ftt _09882_ (
    .a(_04007_),
    .b(_04004_),
    .c(_04010_),
    .y(_04012_)
  );
  al_nand3 _09883_ (
    .a(_00448_),
    .b(_04011_),
    .c(_04012_),
    .y(_04013_)
  );
  al_aoi21 _09884_ (
    .a(TM0),
    .b(\DFF_1525.Q ),
    .c(TM1),
    .y(_04014_)
  );
  al_nand2 _09885_ (
    .a(_04014_),
    .b(_04013_),
    .y(_04015_)
  );
  al_aoi21ttf _09886_ (
    .a(TM0),
    .b(\DFF_1354.Q ),
    .c(TM1),
    .y(_04016_)
  );
  al_and2 _09887_ (
    .a(_04016_),
    .b(_03524_),
    .y(_04017_)
  );
  al_nor3fft _09888_ (
    .a(RESET),
    .b(_04015_),
    .c(_04017_),
    .y(\DFF_1386.D )
  );
  al_or2 _09889_ (
    .a(TM1),
    .b(\DFF_1643.Q ),
    .y(_04018_)
  );
  al_nand2 _09890_ (
    .a(TM1),
    .b(\DFF_1643.Q ),
    .y(_04019_)
  );
  al_nand3 _09891_ (
    .a(\DFF_1675.Q ),
    .b(_04018_),
    .c(_04019_),
    .y(_04020_)
  );
  al_nand2ft _09892_ (
    .a(TM1),
    .b(\DFF_1643.Q ),
    .y(_04021_)
  );
  al_and2ft _09893_ (
    .a(\DFF_1643.Q ),
    .b(TM1),
    .y(_04022_)
  );
  al_and3fft _09894_ (
    .a(\DFF_1675.Q ),
    .b(_04022_),
    .c(_04021_),
    .y(_04023_)
  );
  al_and2ft _09895_ (
    .a(\DFF_1611.Q ),
    .b(\DFF_1579.Q ),
    .y(_04024_)
  );
  al_nand2ft _09896_ (
    .a(\DFF_1579.Q ),
    .b(\DFF_1611.Q ),
    .y(_04025_)
  );
  al_nand2ft _09897_ (
    .a(_04024_),
    .b(_04025_),
    .y(_04026_)
  );
  al_oai21ftf _09898_ (
    .a(_04020_),
    .b(_04023_),
    .c(_04026_),
    .y(_04027_)
  );
  al_nand3ftt _09899_ (
    .a(_04023_),
    .b(_04020_),
    .c(_04026_),
    .y(_04028_)
  );
  al_nand3 _09900_ (
    .a(_00448_),
    .b(_04027_),
    .c(_04028_),
    .y(_04029_)
  );
  al_aoi21 _09901_ (
    .a(TM0),
    .b(\DFF_1524.Q ),
    .c(TM1),
    .y(_04030_)
  );
  al_nand2 _09902_ (
    .a(_04030_),
    .b(_04029_),
    .y(_04031_)
  );
  al_aoi21ttf _09903_ (
    .a(TM0),
    .b(\DFF_1355.Q ),
    .c(TM1),
    .y(_04032_)
  );
  al_and2 _09904_ (
    .a(_04032_),
    .b(_03540_),
    .y(_04033_)
  );
  al_nor3fft _09905_ (
    .a(RESET),
    .b(_04031_),
    .c(_04033_),
    .y(\DFF_1387.D )
  );
  al_or2 _09906_ (
    .a(TM1),
    .b(\DFF_1644.Q ),
    .y(_04034_)
  );
  al_nand2 _09907_ (
    .a(TM1),
    .b(\DFF_1644.Q ),
    .y(_04035_)
  );
  al_nand3 _09908_ (
    .a(\DFF_1676.Q ),
    .b(_04034_),
    .c(_04035_),
    .y(_04036_)
  );
  al_nand2ft _09909_ (
    .a(TM1),
    .b(\DFF_1644.Q ),
    .y(_04037_)
  );
  al_and2ft _09910_ (
    .a(\DFF_1644.Q ),
    .b(TM1),
    .y(_04038_)
  );
  al_and3fft _09911_ (
    .a(\DFF_1676.Q ),
    .b(_04038_),
    .c(_04037_),
    .y(_04039_)
  );
  al_and2ft _09912_ (
    .a(\DFF_1612.Q ),
    .b(\DFF_1580.Q ),
    .y(_04040_)
  );
  al_nand2ft _09913_ (
    .a(\DFF_1580.Q ),
    .b(\DFF_1612.Q ),
    .y(_04041_)
  );
  al_nand2ft _09914_ (
    .a(_04040_),
    .b(_04041_),
    .y(_04042_)
  );
  al_oai21ftf _09915_ (
    .a(_04036_),
    .b(_04039_),
    .c(_04042_),
    .y(_04043_)
  );
  al_nand3ftt _09916_ (
    .a(_04039_),
    .b(_04036_),
    .c(_04042_),
    .y(_04044_)
  );
  al_nand3 _09917_ (
    .a(_00448_),
    .b(_04043_),
    .c(_04044_),
    .y(_04045_)
  );
  al_aoi21 _09918_ (
    .a(TM0),
    .b(\DFF_1523.Q ),
    .c(TM1),
    .y(_04046_)
  );
  al_nand2 _09919_ (
    .a(_04046_),
    .b(_04045_),
    .y(_04047_)
  );
  al_aoi21ttf _09920_ (
    .a(TM0),
    .b(\DFF_1356.Q ),
    .c(TM1),
    .y(_04048_)
  );
  al_and2 _09921_ (
    .a(_04048_),
    .b(_03556_),
    .y(_04049_)
  );
  al_nor3fft _09922_ (
    .a(RESET),
    .b(_04047_),
    .c(_04049_),
    .y(\DFF_1388.D )
  );
  al_or2 _09923_ (
    .a(TM1),
    .b(\DFF_1645.Q ),
    .y(_04050_)
  );
  al_nand2 _09924_ (
    .a(TM1),
    .b(\DFF_1645.Q ),
    .y(_04051_)
  );
  al_nand3 _09925_ (
    .a(\DFF_1677.Q ),
    .b(_04050_),
    .c(_04051_),
    .y(_04052_)
  );
  al_nand2ft _09926_ (
    .a(TM1),
    .b(\DFF_1645.Q ),
    .y(_04053_)
  );
  al_and2ft _09927_ (
    .a(\DFF_1645.Q ),
    .b(TM1),
    .y(_04054_)
  );
  al_and3fft _09928_ (
    .a(\DFF_1677.Q ),
    .b(_04054_),
    .c(_04053_),
    .y(_04055_)
  );
  al_and2ft _09929_ (
    .a(\DFF_1613.Q ),
    .b(\DFF_1581.Q ),
    .y(_04056_)
  );
  al_nand2ft _09930_ (
    .a(\DFF_1581.Q ),
    .b(\DFF_1613.Q ),
    .y(_04057_)
  );
  al_nand2ft _09931_ (
    .a(_04056_),
    .b(_04057_),
    .y(_04058_)
  );
  al_oai21ftf _09932_ (
    .a(_04052_),
    .b(_04055_),
    .c(_04058_),
    .y(_04059_)
  );
  al_nand3ftt _09933_ (
    .a(_04055_),
    .b(_04052_),
    .c(_04058_),
    .y(_04060_)
  );
  al_nand3 _09934_ (
    .a(_00448_),
    .b(_04059_),
    .c(_04060_),
    .y(_04061_)
  );
  al_aoi21 _09935_ (
    .a(TM0),
    .b(\DFF_1522.Q ),
    .c(TM1),
    .y(_04062_)
  );
  al_nand2 _09936_ (
    .a(_04062_),
    .b(_04061_),
    .y(_04063_)
  );
  al_aoi21ttf _09937_ (
    .a(TM0),
    .b(\DFF_1357.Q ),
    .c(TM1),
    .y(_04064_)
  );
  al_and2 _09938_ (
    .a(_04064_),
    .b(_03572_),
    .y(_04065_)
  );
  al_nor3fft _09939_ (
    .a(RESET),
    .b(_04063_),
    .c(_04065_),
    .y(\DFF_1389.D )
  );
  al_or2 _09940_ (
    .a(TM1),
    .b(\DFF_1646.Q ),
    .y(_04066_)
  );
  al_nand2 _09941_ (
    .a(TM1),
    .b(\DFF_1646.Q ),
    .y(_04067_)
  );
  al_nand3 _09942_ (
    .a(\DFF_1678.Q ),
    .b(_04066_),
    .c(_04067_),
    .y(_04068_)
  );
  al_nand2ft _09943_ (
    .a(TM1),
    .b(\DFF_1646.Q ),
    .y(_04069_)
  );
  al_and2ft _09944_ (
    .a(\DFF_1646.Q ),
    .b(TM1),
    .y(_04070_)
  );
  al_and3fft _09945_ (
    .a(\DFF_1678.Q ),
    .b(_04070_),
    .c(_04069_),
    .y(_04071_)
  );
  al_and2ft _09946_ (
    .a(\DFF_1614.Q ),
    .b(\DFF_1582.Q ),
    .y(_04072_)
  );
  al_nand2ft _09947_ (
    .a(\DFF_1582.Q ),
    .b(\DFF_1614.Q ),
    .y(_04073_)
  );
  al_nand2ft _09948_ (
    .a(_04072_),
    .b(_04073_),
    .y(_04074_)
  );
  al_oai21ftf _09949_ (
    .a(_04068_),
    .b(_04071_),
    .c(_04074_),
    .y(_04075_)
  );
  al_nand3ftt _09950_ (
    .a(_04071_),
    .b(_04068_),
    .c(_04074_),
    .y(_04076_)
  );
  al_nand3 _09951_ (
    .a(_00448_),
    .b(_04075_),
    .c(_04076_),
    .y(_04077_)
  );
  al_aoi21 _09952_ (
    .a(TM0),
    .b(\DFF_1521.Q ),
    .c(TM1),
    .y(_04078_)
  );
  al_nand2 _09953_ (
    .a(_04078_),
    .b(_04077_),
    .y(_04079_)
  );
  al_aoi21ttf _09954_ (
    .a(TM0),
    .b(\DFF_1358.Q ),
    .c(TM1),
    .y(_04080_)
  );
  al_and2 _09955_ (
    .a(_04080_),
    .b(_03588_),
    .y(_04081_)
  );
  al_nor3fft _09956_ (
    .a(RESET),
    .b(_04079_),
    .c(_04081_),
    .y(\DFF_1390.D )
  );
  al_or2 _09957_ (
    .a(TM1),
    .b(\DFF_1647.Q ),
    .y(_04082_)
  );
  al_nand2 _09958_ (
    .a(TM1),
    .b(\DFF_1647.Q ),
    .y(_04083_)
  );
  al_nand3 _09959_ (
    .a(\DFF_1679.Q ),
    .b(_04082_),
    .c(_04083_),
    .y(_04084_)
  );
  al_nand2ft _09960_ (
    .a(TM1),
    .b(\DFF_1647.Q ),
    .y(_04085_)
  );
  al_and2ft _09961_ (
    .a(\DFF_1647.Q ),
    .b(TM1),
    .y(_04086_)
  );
  al_and3fft _09962_ (
    .a(\DFF_1679.Q ),
    .b(_04086_),
    .c(_04085_),
    .y(_04087_)
  );
  al_and2ft _09963_ (
    .a(\DFF_1615.Q ),
    .b(\DFF_1583.Q ),
    .y(_04088_)
  );
  al_nand2ft _09964_ (
    .a(\DFF_1583.Q ),
    .b(\DFF_1615.Q ),
    .y(_04089_)
  );
  al_nand2ft _09965_ (
    .a(_04088_),
    .b(_04089_),
    .y(_04090_)
  );
  al_oai21ftf _09966_ (
    .a(_04084_),
    .b(_04087_),
    .c(_04090_),
    .y(_04091_)
  );
  al_nand3ftt _09967_ (
    .a(_04087_),
    .b(_04084_),
    .c(_04090_),
    .y(_04092_)
  );
  al_nand3 _09968_ (
    .a(_00448_),
    .b(_04091_),
    .c(_04092_),
    .y(_04093_)
  );
  al_aoi21 _09969_ (
    .a(TM0),
    .b(\DFF_1520.Q ),
    .c(TM1),
    .y(_04094_)
  );
  al_nand2 _09970_ (
    .a(_04094_),
    .b(_04093_),
    .y(_04095_)
  );
  al_aoi21ttf _09971_ (
    .a(TM0),
    .b(\DFF_1359.Q ),
    .c(TM1),
    .y(_04096_)
  );
  al_and2 _09972_ (
    .a(_04096_),
    .b(_03604_),
    .y(_04097_)
  );
  al_nor3fft _09973_ (
    .a(RESET),
    .b(_04095_),
    .c(_04097_),
    .y(\DFF_1391.D )
  );
  al_aoi21ttf _09974_ (
    .a(TM0),
    .b(\DFF_1360.Q ),
    .c(TM1),
    .y(_04098_)
  );
  al_and2ft _09975_ (
    .a(\DFF_1616.Q ),
    .b(\DFF_1648.Q ),
    .y(_04099_)
  );
  al_nand2ft _09976_ (
    .a(\DFF_1648.Q ),
    .b(\DFF_1616.Q ),
    .y(_04100_)
  );
  al_and2ft _09977_ (
    .a(\DFF_1584.Q ),
    .b(\DFF_1680.Q ),
    .y(_04101_)
  );
  al_nand2ft _09978_ (
    .a(\DFF_1680.Q ),
    .b(\DFF_1584.Q ),
    .y(_04102_)
  );
  al_nand2ft _09979_ (
    .a(_04101_),
    .b(_04102_),
    .y(_04103_)
  );
  al_or3ftt _09980_ (
    .a(_04100_),
    .b(_04099_),
    .c(_04103_),
    .y(_04104_)
  );
  al_ao21ftf _09981_ (
    .a(_04099_),
    .b(_04100_),
    .c(_04103_),
    .y(_04105_)
  );
  al_nand3 _09982_ (
    .a(_00448_),
    .b(_04105_),
    .c(_04104_),
    .y(_04106_)
  );
  al_aoi21 _09983_ (
    .a(TM0),
    .b(\DFF_1519.Q ),
    .c(TM1),
    .y(_04107_)
  );
  al_aoi21 _09984_ (
    .a(_04107_),
    .b(_04106_),
    .c(_00451_),
    .y(_04108_)
  );
  al_aoi21ftf _09985_ (
    .a(_03616_),
    .b(_04098_),
    .c(_04108_),
    .y(\DFF_1392.D )
  );
  al_aoi21ttf _09986_ (
    .a(TM0),
    .b(\DFF_1361.Q ),
    .c(TM1),
    .y(_04109_)
  );
  al_and2ft _09987_ (
    .a(\DFF_1617.Q ),
    .b(\DFF_1649.Q ),
    .y(_04110_)
  );
  al_nand2ft _09988_ (
    .a(\DFF_1649.Q ),
    .b(\DFF_1617.Q ),
    .y(_04111_)
  );
  al_and2ft _09989_ (
    .a(\DFF_1585.Q ),
    .b(\DFF_1681.Q ),
    .y(_04112_)
  );
  al_nand2ft _09990_ (
    .a(\DFF_1681.Q ),
    .b(\DFF_1585.Q ),
    .y(_04113_)
  );
  al_nand2ft _09991_ (
    .a(_04112_),
    .b(_04113_),
    .y(_04114_)
  );
  al_or3ftt _09992_ (
    .a(_04111_),
    .b(_04110_),
    .c(_04114_),
    .y(_04115_)
  );
  al_ao21ftf _09993_ (
    .a(_04110_),
    .b(_04111_),
    .c(_04114_),
    .y(_04116_)
  );
  al_nand3 _09994_ (
    .a(_00448_),
    .b(_04116_),
    .c(_04115_),
    .y(_04117_)
  );
  al_aoi21 _09995_ (
    .a(TM0),
    .b(\DFF_1518.Q ),
    .c(TM1),
    .y(_04118_)
  );
  al_aoi21 _09996_ (
    .a(_04118_),
    .b(_04117_),
    .c(_00451_),
    .y(_04119_)
  );
  al_aoi21ftf _09997_ (
    .a(_03628_),
    .b(_04109_),
    .c(_04119_),
    .y(\DFF_1393.D )
  );
  al_aoi21ttf _09998_ (
    .a(TM0),
    .b(\DFF_1362.Q ),
    .c(TM1),
    .y(_04120_)
  );
  al_and2ft _09999_ (
    .a(\DFF_1618.Q ),
    .b(\DFF_1650.Q ),
    .y(_04121_)
  );
  al_nand2ft _10000_ (
    .a(\DFF_1650.Q ),
    .b(\DFF_1618.Q ),
    .y(_04122_)
  );
  al_and2ft _10001_ (
    .a(\DFF_1586.Q ),
    .b(\DFF_1682.Q ),
    .y(_04123_)
  );
  al_nand2ft _10002_ (
    .a(\DFF_1682.Q ),
    .b(\DFF_1586.Q ),
    .y(_04124_)
  );
  al_nand2ft _10003_ (
    .a(_04123_),
    .b(_04124_),
    .y(_04125_)
  );
  al_or3ftt _10004_ (
    .a(_04122_),
    .b(_04121_),
    .c(_04125_),
    .y(_04126_)
  );
  al_ao21ftf _10005_ (
    .a(_04121_),
    .b(_04122_),
    .c(_04125_),
    .y(_04127_)
  );
  al_nand3 _10006_ (
    .a(_00448_),
    .b(_04127_),
    .c(_04126_),
    .y(_04128_)
  );
  al_aoi21 _10007_ (
    .a(TM0),
    .b(\DFF_1517.Q ),
    .c(TM1),
    .y(_04129_)
  );
  al_aoi21 _10008_ (
    .a(_04129_),
    .b(_04128_),
    .c(_00451_),
    .y(_04130_)
  );
  al_aoi21ftf _10009_ (
    .a(_03640_),
    .b(_04120_),
    .c(_04130_),
    .y(\DFF_1394.D )
  );
  al_aoi21ttf _10010_ (
    .a(TM0),
    .b(\DFF_1363.Q ),
    .c(TM1),
    .y(_04131_)
  );
  al_and2ft _10011_ (
    .a(\DFF_1619.Q ),
    .b(\DFF_1651.Q ),
    .y(_04132_)
  );
  al_nand2ft _10012_ (
    .a(\DFF_1651.Q ),
    .b(\DFF_1619.Q ),
    .y(_04133_)
  );
  al_and2ft _10013_ (
    .a(\DFF_1587.Q ),
    .b(\DFF_1683.Q ),
    .y(_04134_)
  );
  al_nand2ft _10014_ (
    .a(\DFF_1683.Q ),
    .b(\DFF_1587.Q ),
    .y(_04135_)
  );
  al_nand2ft _10015_ (
    .a(_04134_),
    .b(_04135_),
    .y(_04136_)
  );
  al_or3ftt _10016_ (
    .a(_04133_),
    .b(_04132_),
    .c(_04136_),
    .y(_04137_)
  );
  al_ao21ftf _10017_ (
    .a(_04132_),
    .b(_04133_),
    .c(_04136_),
    .y(_04138_)
  );
  al_nand3 _10018_ (
    .a(_00448_),
    .b(_04138_),
    .c(_04137_),
    .y(_04139_)
  );
  al_aoi21 _10019_ (
    .a(TM0),
    .b(\DFF_1516.Q ),
    .c(TM1),
    .y(_04140_)
  );
  al_aoi21 _10020_ (
    .a(_04140_),
    .b(_04139_),
    .c(_00451_),
    .y(_04141_)
  );
  al_aoi21ftf _10021_ (
    .a(_03652_),
    .b(_04131_),
    .c(_04141_),
    .y(\DFF_1395.D )
  );
  al_aoi21ttf _10022_ (
    .a(TM0),
    .b(\DFF_1364.Q ),
    .c(TM1),
    .y(_04142_)
  );
  al_and2ft _10023_ (
    .a(\DFF_1620.Q ),
    .b(\DFF_1652.Q ),
    .y(_04143_)
  );
  al_nand2ft _10024_ (
    .a(\DFF_1652.Q ),
    .b(\DFF_1620.Q ),
    .y(_04144_)
  );
  al_and2ft _10025_ (
    .a(\DFF_1588.Q ),
    .b(\DFF_1684.Q ),
    .y(_04145_)
  );
  al_nand2ft _10026_ (
    .a(\DFF_1684.Q ),
    .b(\DFF_1588.Q ),
    .y(_04146_)
  );
  al_nand2ft _10027_ (
    .a(_04145_),
    .b(_04146_),
    .y(_04147_)
  );
  al_or3ftt _10028_ (
    .a(_04144_),
    .b(_04143_),
    .c(_04147_),
    .y(_04148_)
  );
  al_ao21ftf _10029_ (
    .a(_04143_),
    .b(_04144_),
    .c(_04147_),
    .y(_04149_)
  );
  al_nand3 _10030_ (
    .a(_00448_),
    .b(_04149_),
    .c(_04148_),
    .y(_04150_)
  );
  al_aoi21 _10031_ (
    .a(TM0),
    .b(\DFF_1515.Q ),
    .c(TM1),
    .y(_04151_)
  );
  al_aoi21 _10032_ (
    .a(_04151_),
    .b(_04150_),
    .c(_00451_),
    .y(_04152_)
  );
  al_aoi21ftf _10033_ (
    .a(_03664_),
    .b(_04142_),
    .c(_04152_),
    .y(\DFF_1396.D )
  );
  al_aoi21ttf _10034_ (
    .a(TM0),
    .b(\DFF_1365.Q ),
    .c(TM1),
    .y(_04153_)
  );
  al_and2ft _10035_ (
    .a(\DFF_1621.Q ),
    .b(\DFF_1653.Q ),
    .y(_04154_)
  );
  al_nand2ft _10036_ (
    .a(\DFF_1653.Q ),
    .b(\DFF_1621.Q ),
    .y(_04155_)
  );
  al_and2ft _10037_ (
    .a(\DFF_1589.Q ),
    .b(\DFF_1685.Q ),
    .y(_04156_)
  );
  al_nand2ft _10038_ (
    .a(\DFF_1685.Q ),
    .b(\DFF_1589.Q ),
    .y(_04157_)
  );
  al_nand2ft _10039_ (
    .a(_04156_),
    .b(_04157_),
    .y(_04158_)
  );
  al_or3ftt _10040_ (
    .a(_04155_),
    .b(_04154_),
    .c(_04158_),
    .y(_04159_)
  );
  al_ao21ftf _10041_ (
    .a(_04154_),
    .b(_04155_),
    .c(_04158_),
    .y(_04160_)
  );
  al_nand3 _10042_ (
    .a(_00448_),
    .b(_04160_),
    .c(_04159_),
    .y(_04161_)
  );
  al_aoi21 _10043_ (
    .a(TM0),
    .b(\DFF_1514.Q ),
    .c(TM1),
    .y(_04162_)
  );
  al_aoi21 _10044_ (
    .a(_04162_),
    .b(_04161_),
    .c(_00451_),
    .y(_04163_)
  );
  al_aoi21ftf _10045_ (
    .a(_03676_),
    .b(_04153_),
    .c(_04163_),
    .y(\DFF_1397.D )
  );
  al_aoi21ttf _10046_ (
    .a(TM0),
    .b(\DFF_1366.Q ),
    .c(TM1),
    .y(_04164_)
  );
  al_and2ft _10047_ (
    .a(\DFF_1622.Q ),
    .b(\DFF_1654.Q ),
    .y(_04165_)
  );
  al_nand2ft _10048_ (
    .a(\DFF_1654.Q ),
    .b(\DFF_1622.Q ),
    .y(_04166_)
  );
  al_and2ft _10049_ (
    .a(\DFF_1590.Q ),
    .b(\DFF_1686.Q ),
    .y(_04167_)
  );
  al_nand2ft _10050_ (
    .a(\DFF_1686.Q ),
    .b(\DFF_1590.Q ),
    .y(_04168_)
  );
  al_nand2ft _10051_ (
    .a(_04167_),
    .b(_04168_),
    .y(_04169_)
  );
  al_or3ftt _10052_ (
    .a(_04166_),
    .b(_04165_),
    .c(_04169_),
    .y(_04170_)
  );
  al_ao21ftf _10053_ (
    .a(_04165_),
    .b(_04166_),
    .c(_04169_),
    .y(_04171_)
  );
  al_nand3 _10054_ (
    .a(_00448_),
    .b(_04171_),
    .c(_04170_),
    .y(_04172_)
  );
  al_aoi21 _10055_ (
    .a(TM0),
    .b(\DFF_1513.Q ),
    .c(TM1),
    .y(_04173_)
  );
  al_aoi21 _10056_ (
    .a(_04173_),
    .b(_04172_),
    .c(_00451_),
    .y(_04174_)
  );
  al_aoi21ftf _10057_ (
    .a(_03688_),
    .b(_04164_),
    .c(_04174_),
    .y(\DFF_1398.D )
  );
  al_aoi21ttf _10058_ (
    .a(TM0),
    .b(\DFF_1367.Q ),
    .c(TM1),
    .y(_04175_)
  );
  al_and2ft _10059_ (
    .a(\DFF_1623.Q ),
    .b(\DFF_1655.Q ),
    .y(_04176_)
  );
  al_nand2ft _10060_ (
    .a(\DFF_1655.Q ),
    .b(\DFF_1623.Q ),
    .y(_04177_)
  );
  al_and2ft _10061_ (
    .a(\DFF_1591.Q ),
    .b(\DFF_1687.Q ),
    .y(_04178_)
  );
  al_nand2ft _10062_ (
    .a(\DFF_1687.Q ),
    .b(\DFF_1591.Q ),
    .y(_04179_)
  );
  al_nand2ft _10063_ (
    .a(_04178_),
    .b(_04179_),
    .y(_04180_)
  );
  al_or3ftt _10064_ (
    .a(_04177_),
    .b(_04176_),
    .c(_04180_),
    .y(_04181_)
  );
  al_ao21ftf _10065_ (
    .a(_04176_),
    .b(_04177_),
    .c(_04180_),
    .y(_04182_)
  );
  al_nand3 _10066_ (
    .a(_00448_),
    .b(_04182_),
    .c(_04181_),
    .y(_04183_)
  );
  al_aoi21 _10067_ (
    .a(TM0),
    .b(\DFF_1512.Q ),
    .c(TM1),
    .y(_04184_)
  );
  al_aoi21 _10068_ (
    .a(_04184_),
    .b(_04183_),
    .c(_00451_),
    .y(_04185_)
  );
  al_aoi21ftf _10069_ (
    .a(_03700_),
    .b(_04175_),
    .c(_04185_),
    .y(\DFF_1399.D )
  );
  al_aoi21ttf _10070_ (
    .a(TM0),
    .b(\DFF_1368.Q ),
    .c(TM1),
    .y(_04186_)
  );
  al_and2ft _10071_ (
    .a(\DFF_1624.Q ),
    .b(\DFF_1656.Q ),
    .y(_04187_)
  );
  al_nand2ft _10072_ (
    .a(\DFF_1656.Q ),
    .b(\DFF_1624.Q ),
    .y(_04188_)
  );
  al_and2ft _10073_ (
    .a(\DFF_1592.Q ),
    .b(\DFF_1688.Q ),
    .y(_04189_)
  );
  al_nand2ft _10074_ (
    .a(\DFF_1688.Q ),
    .b(\DFF_1592.Q ),
    .y(_04190_)
  );
  al_nand2ft _10075_ (
    .a(_04189_),
    .b(_04190_),
    .y(_04191_)
  );
  al_or3ftt _10076_ (
    .a(_04188_),
    .b(_04187_),
    .c(_04191_),
    .y(_04192_)
  );
  al_ao21ftf _10077_ (
    .a(_04187_),
    .b(_04188_),
    .c(_04191_),
    .y(_04193_)
  );
  al_nand3 _10078_ (
    .a(_00448_),
    .b(_04193_),
    .c(_04192_),
    .y(_04194_)
  );
  al_aoi21 _10079_ (
    .a(TM0),
    .b(\DFF_1511.Q ),
    .c(TM1),
    .y(_04195_)
  );
  al_aoi21 _10080_ (
    .a(_04195_),
    .b(_04194_),
    .c(_00451_),
    .y(_04196_)
  );
  al_aoi21ftf _10081_ (
    .a(_03712_),
    .b(_04186_),
    .c(_04196_),
    .y(\DFF_1400.D )
  );
  al_aoi21ttf _10082_ (
    .a(TM0),
    .b(\DFF_1369.Q ),
    .c(TM1),
    .y(_04197_)
  );
  al_and2ft _10083_ (
    .a(\DFF_1625.Q ),
    .b(\DFF_1657.Q ),
    .y(_04198_)
  );
  al_nand2ft _10084_ (
    .a(\DFF_1657.Q ),
    .b(\DFF_1625.Q ),
    .y(_04199_)
  );
  al_and2ft _10085_ (
    .a(\DFF_1593.Q ),
    .b(\DFF_1689.Q ),
    .y(_04200_)
  );
  al_nand2ft _10086_ (
    .a(\DFF_1689.Q ),
    .b(\DFF_1593.Q ),
    .y(_04201_)
  );
  al_nand2ft _10087_ (
    .a(_04200_),
    .b(_04201_),
    .y(_04202_)
  );
  al_or3ftt _10088_ (
    .a(_04199_),
    .b(_04198_),
    .c(_04202_),
    .y(_04203_)
  );
  al_ao21ftf _10089_ (
    .a(_04198_),
    .b(_04199_),
    .c(_04202_),
    .y(_04204_)
  );
  al_nand3 _10090_ (
    .a(_00448_),
    .b(_04204_),
    .c(_04203_),
    .y(_04205_)
  );
  al_aoi21 _10091_ (
    .a(TM0),
    .b(\DFF_1510.Q ),
    .c(TM1),
    .y(_04206_)
  );
  al_aoi21 _10092_ (
    .a(_04206_),
    .b(_04205_),
    .c(_00451_),
    .y(_04207_)
  );
  al_aoi21ftf _10093_ (
    .a(_03724_),
    .b(_04197_),
    .c(_04207_),
    .y(\DFF_1401.D )
  );
  al_aoi21ttf _10094_ (
    .a(TM0),
    .b(\DFF_1370.Q ),
    .c(TM1),
    .y(_04208_)
  );
  al_and2ft _10095_ (
    .a(\DFF_1626.Q ),
    .b(\DFF_1658.Q ),
    .y(_04209_)
  );
  al_nand2ft _10096_ (
    .a(\DFF_1658.Q ),
    .b(\DFF_1626.Q ),
    .y(_04210_)
  );
  al_and2ft _10097_ (
    .a(\DFF_1594.Q ),
    .b(\DFF_1690.Q ),
    .y(_04211_)
  );
  al_nand2ft _10098_ (
    .a(\DFF_1690.Q ),
    .b(\DFF_1594.Q ),
    .y(_04212_)
  );
  al_nand2ft _10099_ (
    .a(_04211_),
    .b(_04212_),
    .y(_04213_)
  );
  al_or3ftt _10100_ (
    .a(_04210_),
    .b(_04209_),
    .c(_04213_),
    .y(_04214_)
  );
  al_ao21ftf _10101_ (
    .a(_04209_),
    .b(_04210_),
    .c(_04213_),
    .y(_04215_)
  );
  al_nand3 _10102_ (
    .a(_00448_),
    .b(_04215_),
    .c(_04214_),
    .y(_04216_)
  );
  al_aoi21 _10103_ (
    .a(TM0),
    .b(\DFF_1509.Q ),
    .c(TM1),
    .y(_04217_)
  );
  al_aoi21 _10104_ (
    .a(_04217_),
    .b(_04216_),
    .c(_00451_),
    .y(_04218_)
  );
  al_aoi21ftf _10105_ (
    .a(_03736_),
    .b(_04208_),
    .c(_04218_),
    .y(\DFF_1402.D )
  );
  al_aoi21ttf _10106_ (
    .a(TM0),
    .b(\DFF_1371.Q ),
    .c(TM1),
    .y(_04219_)
  );
  al_and2ft _10107_ (
    .a(\DFF_1627.Q ),
    .b(\DFF_1659.Q ),
    .y(_04220_)
  );
  al_nand2ft _10108_ (
    .a(\DFF_1659.Q ),
    .b(\DFF_1627.Q ),
    .y(_04221_)
  );
  al_and2ft _10109_ (
    .a(\DFF_1595.Q ),
    .b(\DFF_1691.Q ),
    .y(_04222_)
  );
  al_nand2ft _10110_ (
    .a(\DFF_1691.Q ),
    .b(\DFF_1595.Q ),
    .y(_04223_)
  );
  al_nand2ft _10111_ (
    .a(_04222_),
    .b(_04223_),
    .y(_04224_)
  );
  al_or3ftt _10112_ (
    .a(_04221_),
    .b(_04220_),
    .c(_04224_),
    .y(_04225_)
  );
  al_ao21ftf _10113_ (
    .a(_04220_),
    .b(_04221_),
    .c(_04224_),
    .y(_04226_)
  );
  al_nand3 _10114_ (
    .a(_00448_),
    .b(_04226_),
    .c(_04225_),
    .y(_04227_)
  );
  al_aoi21 _10115_ (
    .a(TM0),
    .b(\DFF_1508.Q ),
    .c(TM1),
    .y(_04228_)
  );
  al_aoi21 _10116_ (
    .a(_04228_),
    .b(_04227_),
    .c(_00451_),
    .y(_04229_)
  );
  al_aoi21ftf _10117_ (
    .a(_03748_),
    .b(_04219_),
    .c(_04229_),
    .y(\DFF_1403.D )
  );
  al_aoi21ttf _10118_ (
    .a(TM0),
    .b(\DFF_1372.Q ),
    .c(TM1),
    .y(_04230_)
  );
  al_and2ft _10119_ (
    .a(\DFF_1628.Q ),
    .b(\DFF_1660.Q ),
    .y(_04231_)
  );
  al_nand2ft _10120_ (
    .a(\DFF_1660.Q ),
    .b(\DFF_1628.Q ),
    .y(_04232_)
  );
  al_and2ft _10121_ (
    .a(\DFF_1596.Q ),
    .b(\DFF_1692.Q ),
    .y(_04233_)
  );
  al_nand2ft _10122_ (
    .a(\DFF_1692.Q ),
    .b(\DFF_1596.Q ),
    .y(_04234_)
  );
  al_nand2ft _10123_ (
    .a(_04233_),
    .b(_04234_),
    .y(_04235_)
  );
  al_or3ftt _10124_ (
    .a(_04232_),
    .b(_04231_),
    .c(_04235_),
    .y(_04236_)
  );
  al_ao21ftf _10125_ (
    .a(_04231_),
    .b(_04232_),
    .c(_04235_),
    .y(_04237_)
  );
  al_nand3 _10126_ (
    .a(_00448_),
    .b(_04237_),
    .c(_04236_),
    .y(_04238_)
  );
  al_aoi21 _10127_ (
    .a(TM0),
    .b(\DFF_1507.Q ),
    .c(TM1),
    .y(_04239_)
  );
  al_aoi21 _10128_ (
    .a(_04239_),
    .b(_04238_),
    .c(_00451_),
    .y(_04240_)
  );
  al_aoi21ftf _10129_ (
    .a(_03760_),
    .b(_04230_),
    .c(_04240_),
    .y(\DFF_1404.D )
  );
  al_aoi21ttf _10130_ (
    .a(TM0),
    .b(\DFF_1373.Q ),
    .c(TM1),
    .y(_04241_)
  );
  al_and2ft _10131_ (
    .a(\DFF_1629.Q ),
    .b(\DFF_1661.Q ),
    .y(_04242_)
  );
  al_nand2ft _10132_ (
    .a(\DFF_1661.Q ),
    .b(\DFF_1629.Q ),
    .y(_04243_)
  );
  al_and2ft _10133_ (
    .a(\DFF_1597.Q ),
    .b(\DFF_1693.Q ),
    .y(_04244_)
  );
  al_nand2ft _10134_ (
    .a(\DFF_1693.Q ),
    .b(\DFF_1597.Q ),
    .y(_04245_)
  );
  al_nand2ft _10135_ (
    .a(_04244_),
    .b(_04245_),
    .y(_04246_)
  );
  al_or3ftt _10136_ (
    .a(_04243_),
    .b(_04242_),
    .c(_04246_),
    .y(_04247_)
  );
  al_ao21ftf _10137_ (
    .a(_04242_),
    .b(_04243_),
    .c(_04246_),
    .y(_04248_)
  );
  al_nand3 _10138_ (
    .a(_00448_),
    .b(_04248_),
    .c(_04247_),
    .y(_04249_)
  );
  al_aoi21 _10139_ (
    .a(TM0),
    .b(\DFF_1506.Q ),
    .c(TM1),
    .y(_04250_)
  );
  al_aoi21 _10140_ (
    .a(_04250_),
    .b(_04249_),
    .c(_00451_),
    .y(_04251_)
  );
  al_aoi21ftf _10141_ (
    .a(_03772_),
    .b(_04241_),
    .c(_04251_),
    .y(\DFF_1405.D )
  );
  al_aoi21ttf _10142_ (
    .a(TM0),
    .b(\DFF_1374.Q ),
    .c(TM1),
    .y(_04252_)
  );
  al_and2ft _10143_ (
    .a(\DFF_1630.Q ),
    .b(\DFF_1662.Q ),
    .y(_04253_)
  );
  al_nand2ft _10144_ (
    .a(\DFF_1662.Q ),
    .b(\DFF_1630.Q ),
    .y(_04254_)
  );
  al_and2ft _10145_ (
    .a(\DFF_1598.Q ),
    .b(\DFF_1694.Q ),
    .y(_04255_)
  );
  al_nand2ft _10146_ (
    .a(\DFF_1694.Q ),
    .b(\DFF_1598.Q ),
    .y(_04256_)
  );
  al_nand2ft _10147_ (
    .a(_04255_),
    .b(_04256_),
    .y(_04257_)
  );
  al_or3ftt _10148_ (
    .a(_04254_),
    .b(_04253_),
    .c(_04257_),
    .y(_04258_)
  );
  al_ao21ftf _10149_ (
    .a(_04253_),
    .b(_04254_),
    .c(_04257_),
    .y(_04259_)
  );
  al_nand3 _10150_ (
    .a(_00448_),
    .b(_04259_),
    .c(_04258_),
    .y(_04260_)
  );
  al_aoi21 _10151_ (
    .a(TM0),
    .b(\DFF_1505.Q ),
    .c(TM1),
    .y(_04261_)
  );
  al_aoi21 _10152_ (
    .a(_04261_),
    .b(_04260_),
    .c(_00451_),
    .y(_04262_)
  );
  al_aoi21ftf _10153_ (
    .a(_03784_),
    .b(_04252_),
    .c(_04262_),
    .y(\DFF_1406.D )
  );
  al_aoi21ttf _10154_ (
    .a(TM0),
    .b(\DFF_1375.Q ),
    .c(TM1),
    .y(_04263_)
  );
  al_and2ft _10155_ (
    .a(\DFF_1631.Q ),
    .b(\DFF_1663.Q ),
    .y(_04264_)
  );
  al_nand2ft _10156_ (
    .a(\DFF_1663.Q ),
    .b(\DFF_1631.Q ),
    .y(_04265_)
  );
  al_and2ft _10157_ (
    .a(\DFF_1599.Q ),
    .b(\DFF_1695.Q ),
    .y(_04266_)
  );
  al_nand2ft _10158_ (
    .a(\DFF_1695.Q ),
    .b(\DFF_1599.Q ),
    .y(_04267_)
  );
  al_nand2ft _10159_ (
    .a(_04266_),
    .b(_04267_),
    .y(_04268_)
  );
  al_or3ftt _10160_ (
    .a(_04265_),
    .b(_04264_),
    .c(_04268_),
    .y(_04269_)
  );
  al_ao21ftf _10161_ (
    .a(_04264_),
    .b(_04265_),
    .c(_04268_),
    .y(_04270_)
  );
  al_nand3 _10162_ (
    .a(_00448_),
    .b(_04270_),
    .c(_04269_),
    .y(_04271_)
  );
  al_aoi21 _10163_ (
    .a(TM0),
    .b(\DFF_1504.Q ),
    .c(TM1),
    .y(_04272_)
  );
  al_aoi21 _10164_ (
    .a(_04272_),
    .b(_04271_),
    .c(_00451_),
    .y(_04273_)
  );
  al_aoi21ftf _10165_ (
    .a(_03796_),
    .b(_04263_),
    .c(_04273_),
    .y(\DFF_1407.D )
  );
  al_and2 _10166_ (
    .a(RESET),
    .b(\DFF_1376.Q ),
    .y(\DFF_1408.D )
  );
  al_and2 _10167_ (
    .a(RESET),
    .b(\DFF_1377.Q ),
    .y(\DFF_1409.D )
  );
  al_and2 _10168_ (
    .a(RESET),
    .b(\DFF_1378.Q ),
    .y(\DFF_1410.D )
  );
  al_and2 _10169_ (
    .a(RESET),
    .b(\DFF_1379.Q ),
    .y(\DFF_1411.D )
  );
  al_and2 _10170_ (
    .a(RESET),
    .b(\DFF_1380.Q ),
    .y(\DFF_1412.D )
  );
  al_and2 _10171_ (
    .a(RESET),
    .b(\DFF_1381.Q ),
    .y(\DFF_1413.D )
  );
  al_and2 _10172_ (
    .a(RESET),
    .b(\DFF_1382.Q ),
    .y(\DFF_1414.D )
  );
  al_and2 _10173_ (
    .a(RESET),
    .b(\DFF_1383.Q ),
    .y(\DFF_1415.D )
  );
  al_and2 _10174_ (
    .a(RESET),
    .b(\DFF_1384.Q ),
    .y(\DFF_1416.D )
  );
  al_and2 _10175_ (
    .a(RESET),
    .b(\DFF_1385.Q ),
    .y(\DFF_1417.D )
  );
  al_and2 _10176_ (
    .a(RESET),
    .b(\DFF_1386.Q ),
    .y(\DFF_1418.D )
  );
  al_and2 _10177_ (
    .a(RESET),
    .b(\DFF_1387.Q ),
    .y(\DFF_1419.D )
  );
  al_and2 _10178_ (
    .a(RESET),
    .b(\DFF_1388.Q ),
    .y(\DFF_1420.D )
  );
  al_and2 _10179_ (
    .a(RESET),
    .b(\DFF_1389.Q ),
    .y(\DFF_1421.D )
  );
  al_and2 _10180_ (
    .a(RESET),
    .b(\DFF_1390.Q ),
    .y(\DFF_1422.D )
  );
  al_and2 _10181_ (
    .a(RESET),
    .b(\DFF_1391.Q ),
    .y(\DFF_1423.D )
  );
  al_and2 _10182_ (
    .a(RESET),
    .b(\DFF_1392.Q ),
    .y(\DFF_1424.D )
  );
  al_and2 _10183_ (
    .a(RESET),
    .b(\DFF_1393.Q ),
    .y(\DFF_1425.D )
  );
  al_and2 _10184_ (
    .a(RESET),
    .b(\DFF_1394.Q ),
    .y(\DFF_1426.D )
  );
  al_and2 _10185_ (
    .a(RESET),
    .b(\DFF_1395.Q ),
    .y(\DFF_1427.D )
  );
  al_and2 _10186_ (
    .a(RESET),
    .b(\DFF_1396.Q ),
    .y(\DFF_1428.D )
  );
  al_and2 _10187_ (
    .a(RESET),
    .b(\DFF_1397.Q ),
    .y(\DFF_1429.D )
  );
  al_and2 _10188_ (
    .a(RESET),
    .b(\DFF_1398.Q ),
    .y(\DFF_1430.D )
  );
  al_and2 _10189_ (
    .a(RESET),
    .b(\DFF_1399.Q ),
    .y(\DFF_1431.D )
  );
  al_and2 _10190_ (
    .a(RESET),
    .b(\DFF_1400.Q ),
    .y(\DFF_1432.D )
  );
  al_and2 _10191_ (
    .a(RESET),
    .b(\DFF_1401.Q ),
    .y(\DFF_1433.D )
  );
  al_and2 _10192_ (
    .a(RESET),
    .b(\DFF_1402.Q ),
    .y(\DFF_1434.D )
  );
  al_and2 _10193_ (
    .a(RESET),
    .b(\DFF_1403.Q ),
    .y(\DFF_1435.D )
  );
  al_and2 _10194_ (
    .a(RESET),
    .b(\DFF_1404.Q ),
    .y(\DFF_1436.D )
  );
  al_and2 _10195_ (
    .a(RESET),
    .b(\DFF_1405.Q ),
    .y(\DFF_1437.D )
  );
  al_and2 _10196_ (
    .a(RESET),
    .b(\DFF_1406.Q ),
    .y(\DFF_1438.D )
  );
  al_and2 _10197_ (
    .a(RESET),
    .b(\DFF_1407.Q ),
    .y(\DFF_1439.D )
  );
  al_and2 _10198_ (
    .a(RESET),
    .b(\DFF_1408.Q ),
    .y(\DFF_1440.D )
  );
  al_and2 _10199_ (
    .a(RESET),
    .b(\DFF_1409.Q ),
    .y(\DFF_1441.D )
  );
  al_and2 _10200_ (
    .a(RESET),
    .b(\DFF_1410.Q ),
    .y(\DFF_1442.D )
  );
  al_and2 _10201_ (
    .a(RESET),
    .b(\DFF_1411.Q ),
    .y(\DFF_1443.D )
  );
  al_and2 _10202_ (
    .a(RESET),
    .b(\DFF_1412.Q ),
    .y(\DFF_1444.D )
  );
  al_and2 _10203_ (
    .a(RESET),
    .b(\DFF_1413.Q ),
    .y(\DFF_1445.D )
  );
  al_and2 _10204_ (
    .a(RESET),
    .b(\DFF_1414.Q ),
    .y(\DFF_1446.D )
  );
  al_and2 _10205_ (
    .a(RESET),
    .b(\DFF_1415.Q ),
    .y(\DFF_1447.D )
  );
  al_and2 _10206_ (
    .a(RESET),
    .b(\DFF_1416.Q ),
    .y(\DFF_1448.D )
  );
  al_and2 _10207_ (
    .a(RESET),
    .b(\DFF_1417.Q ),
    .y(\DFF_1449.D )
  );
  al_and2 _10208_ (
    .a(RESET),
    .b(\DFF_1418.Q ),
    .y(\DFF_1450.D )
  );
  al_and2 _10209_ (
    .a(RESET),
    .b(\DFF_1419.Q ),
    .y(\DFF_1451.D )
  );
  al_and2 _10210_ (
    .a(RESET),
    .b(\DFF_1420.Q ),
    .y(\DFF_1452.D )
  );
  al_and2 _10211_ (
    .a(RESET),
    .b(\DFF_1421.Q ),
    .y(\DFF_1453.D )
  );
  al_and2 _10212_ (
    .a(RESET),
    .b(\DFF_1422.Q ),
    .y(\DFF_1454.D )
  );
  al_and2 _10213_ (
    .a(RESET),
    .b(\DFF_1423.Q ),
    .y(\DFF_1455.D )
  );
  al_and2 _10214_ (
    .a(RESET),
    .b(\DFF_1424.Q ),
    .y(\DFF_1456.D )
  );
  al_and2 _10215_ (
    .a(RESET),
    .b(\DFF_1425.Q ),
    .y(\DFF_1457.D )
  );
  al_and2 _10216_ (
    .a(RESET),
    .b(\DFF_1426.Q ),
    .y(\DFF_1458.D )
  );
  al_and2 _10217_ (
    .a(RESET),
    .b(\DFF_1427.Q ),
    .y(\DFF_1459.D )
  );
  al_and2 _10218_ (
    .a(RESET),
    .b(\DFF_1428.Q ),
    .y(\DFF_1460.D )
  );
  al_and2 _10219_ (
    .a(RESET),
    .b(\DFF_1429.Q ),
    .y(\DFF_1461.D )
  );
  al_and2 _10220_ (
    .a(RESET),
    .b(\DFF_1430.Q ),
    .y(\DFF_1462.D )
  );
  al_and2 _10221_ (
    .a(RESET),
    .b(\DFF_1431.Q ),
    .y(\DFF_1463.D )
  );
  al_and2 _10222_ (
    .a(RESET),
    .b(\DFF_1432.Q ),
    .y(\DFF_1464.D )
  );
  al_and2 _10223_ (
    .a(RESET),
    .b(\DFF_1433.Q ),
    .y(\DFF_1465.D )
  );
  al_and2 _10224_ (
    .a(RESET),
    .b(\DFF_1434.Q ),
    .y(\DFF_1466.D )
  );
  al_and2 _10225_ (
    .a(RESET),
    .b(\DFF_1435.Q ),
    .y(\DFF_1467.D )
  );
  al_and2 _10226_ (
    .a(RESET),
    .b(\DFF_1436.Q ),
    .y(\DFF_1468.D )
  );
  al_and2 _10227_ (
    .a(RESET),
    .b(\DFF_1437.Q ),
    .y(\DFF_1469.D )
  );
  al_and2 _10228_ (
    .a(RESET),
    .b(\DFF_1438.Q ),
    .y(\DFF_1470.D )
  );
  al_and2 _10229_ (
    .a(RESET),
    .b(\DFF_1439.Q ),
    .y(\DFF_1471.D )
  );
  al_and2 _10230_ (
    .a(RESET),
    .b(\DFF_1440.Q ),
    .y(\DFF_1472.D )
  );
  al_and2 _10231_ (
    .a(RESET),
    .b(\DFF_1441.Q ),
    .y(\DFF_1473.D )
  );
  al_and2 _10232_ (
    .a(RESET),
    .b(\DFF_1442.Q ),
    .y(\DFF_1474.D )
  );
  al_and2 _10233_ (
    .a(RESET),
    .b(\DFF_1443.Q ),
    .y(\DFF_1475.D )
  );
  al_and2 _10234_ (
    .a(RESET),
    .b(\DFF_1444.Q ),
    .y(\DFF_1476.D )
  );
  al_and2 _10235_ (
    .a(RESET),
    .b(\DFF_1445.Q ),
    .y(\DFF_1477.D )
  );
  al_and2 _10236_ (
    .a(RESET),
    .b(\DFF_1446.Q ),
    .y(\DFF_1478.D )
  );
  al_and2 _10237_ (
    .a(RESET),
    .b(\DFF_1447.Q ),
    .y(\DFF_1479.D )
  );
  al_and2 _10238_ (
    .a(RESET),
    .b(\DFF_1448.Q ),
    .y(\DFF_1480.D )
  );
  al_and2 _10239_ (
    .a(RESET),
    .b(\DFF_1449.Q ),
    .y(\DFF_1481.D )
  );
  al_and2 _10240_ (
    .a(RESET),
    .b(\DFF_1450.Q ),
    .y(\DFF_1482.D )
  );
  al_and2 _10241_ (
    .a(RESET),
    .b(\DFF_1451.Q ),
    .y(\DFF_1483.D )
  );
  al_and2 _10242_ (
    .a(RESET),
    .b(\DFF_1452.Q ),
    .y(\DFF_1484.D )
  );
  al_and2 _10243_ (
    .a(RESET),
    .b(\DFF_1453.Q ),
    .y(\DFF_1485.D )
  );
  al_and2 _10244_ (
    .a(RESET),
    .b(\DFF_1454.Q ),
    .y(\DFF_1486.D )
  );
  al_and2 _10245_ (
    .a(RESET),
    .b(\DFF_1455.Q ),
    .y(\DFF_1487.D )
  );
  al_and2 _10246_ (
    .a(RESET),
    .b(\DFF_1456.Q ),
    .y(\DFF_1488.D )
  );
  al_and2 _10247_ (
    .a(RESET),
    .b(\DFF_1457.Q ),
    .y(\DFF_1489.D )
  );
  al_and2 _10248_ (
    .a(RESET),
    .b(\DFF_1458.Q ),
    .y(\DFF_1490.D )
  );
  al_and2 _10249_ (
    .a(RESET),
    .b(\DFF_1459.Q ),
    .y(\DFF_1491.D )
  );
  al_and2 _10250_ (
    .a(RESET),
    .b(\DFF_1460.Q ),
    .y(\DFF_1492.D )
  );
  al_and2 _10251_ (
    .a(RESET),
    .b(\DFF_1461.Q ),
    .y(\DFF_1493.D )
  );
  al_and2 _10252_ (
    .a(RESET),
    .b(\DFF_1462.Q ),
    .y(\DFF_1494.D )
  );
  al_and2 _10253_ (
    .a(RESET),
    .b(\DFF_1463.Q ),
    .y(\DFF_1495.D )
  );
  al_and2 _10254_ (
    .a(RESET),
    .b(\DFF_1464.Q ),
    .y(\DFF_1496.D )
  );
  al_and2 _10255_ (
    .a(RESET),
    .b(\DFF_1465.Q ),
    .y(\DFF_1497.D )
  );
  al_and2 _10256_ (
    .a(RESET),
    .b(\DFF_1466.Q ),
    .y(\DFF_1498.D )
  );
  al_and2 _10257_ (
    .a(RESET),
    .b(\DFF_1467.Q ),
    .y(\DFF_1499.D )
  );
  al_and2 _10258_ (
    .a(RESET),
    .b(\DFF_1468.Q ),
    .y(\DFF_1500.D )
  );
  al_and2 _10259_ (
    .a(RESET),
    .b(\DFF_1469.Q ),
    .y(\DFF_1501.D )
  );
  al_and2 _10260_ (
    .a(RESET),
    .b(\DFF_1470.Q ),
    .y(\DFF_1502.D )
  );
  al_and2 _10261_ (
    .a(RESET),
    .b(\DFF_1471.Q ),
    .y(\DFF_1503.D )
  );
  al_oa21ftt _10262_ (
    .a(\DFF_1503.Q ),
    .b(\DFF_1535.Q ),
    .c(RESET),
    .y(_04274_)
  );
  al_aoi21ftf _10263_ (
    .a(\DFF_1503.Q ),
    .b(\DFF_1535.Q ),
    .c(_04274_),
    .y(\DFF_1504.D )
  );
  al_oa21ftt _10264_ (
    .a(\DFF_1502.Q ),
    .b(\DFF_1504.Q ),
    .c(RESET),
    .y(_04275_)
  );
  al_aoi21ftf _10265_ (
    .a(\DFF_1502.Q ),
    .b(\DFF_1504.Q ),
    .c(_04275_),
    .y(\DFF_1505.D )
  );
  al_oa21ftt _10266_ (
    .a(\DFF_1501.Q ),
    .b(\DFF_1505.Q ),
    .c(RESET),
    .y(_04276_)
  );
  al_aoi21ftf _10267_ (
    .a(\DFF_1501.Q ),
    .b(\DFF_1505.Q ),
    .c(_04276_),
    .y(\DFF_1506.D )
  );
  al_oa21ftt _10268_ (
    .a(\DFF_1500.Q ),
    .b(\DFF_1506.Q ),
    .c(RESET),
    .y(_04277_)
  );
  al_aoi21ftf _10269_ (
    .a(\DFF_1500.Q ),
    .b(\DFF_1506.Q ),
    .c(_04277_),
    .y(\DFF_1507.D )
  );
  al_nand2ft _10270_ (
    .a(\DFF_1499.Q ),
    .b(\DFF_1507.Q ),
    .y(_04278_)
  );
  al_nand2ft _10271_ (
    .a(\DFF_1507.Q ),
    .b(\DFF_1499.Q ),
    .y(_04279_)
  );
  al_ao21ttf _10272_ (
    .a(_04278_),
    .b(_04279_),
    .c(\DFF_1535.Q ),
    .y(_04280_)
  );
  al_nand3ftt _10273_ (
    .a(\DFF_1535.Q ),
    .b(_04278_),
    .c(_04279_),
    .y(_04281_)
  );
  al_aoi21 _10274_ (
    .a(_04281_),
    .b(_04280_),
    .c(_00451_),
    .y(\DFF_1508.D )
  );
  al_oa21ftt _10275_ (
    .a(\DFF_1498.Q ),
    .b(\DFF_1508.Q ),
    .c(RESET),
    .y(_04282_)
  );
  al_aoi21ftf _10276_ (
    .a(\DFF_1498.Q ),
    .b(\DFF_1508.Q ),
    .c(_04282_),
    .y(\DFF_1509.D )
  );
  al_oa21ftt _10277_ (
    .a(\DFF_1497.Q ),
    .b(\DFF_1509.Q ),
    .c(RESET),
    .y(_04283_)
  );
  al_aoi21ftf _10278_ (
    .a(\DFF_1497.Q ),
    .b(\DFF_1509.Q ),
    .c(_04283_),
    .y(\DFF_1510.D )
  );
  al_oa21ftt _10279_ (
    .a(\DFF_1496.Q ),
    .b(\DFF_1510.Q ),
    .c(RESET),
    .y(_04284_)
  );
  al_aoi21ftf _10280_ (
    .a(\DFF_1496.Q ),
    .b(\DFF_1510.Q ),
    .c(_04284_),
    .y(\DFF_1511.D )
  );
  al_oa21ftt _10281_ (
    .a(\DFF_1495.Q ),
    .b(\DFF_1511.Q ),
    .c(RESET),
    .y(_04285_)
  );
  al_aoi21ftf _10282_ (
    .a(\DFF_1495.Q ),
    .b(\DFF_1511.Q ),
    .c(_04285_),
    .y(\DFF_1512.D )
  );
  al_oa21ftt _10283_ (
    .a(\DFF_1494.Q ),
    .b(\DFF_1512.Q ),
    .c(RESET),
    .y(_04286_)
  );
  al_aoi21ftf _10284_ (
    .a(\DFF_1494.Q ),
    .b(\DFF_1512.Q ),
    .c(_04286_),
    .y(\DFF_1513.D )
  );
  al_oa21ftt _10285_ (
    .a(\DFF_1493.Q ),
    .b(\DFF_1513.Q ),
    .c(RESET),
    .y(_04287_)
  );
  al_aoi21ftf _10286_ (
    .a(\DFF_1493.Q ),
    .b(\DFF_1513.Q ),
    .c(_04287_),
    .y(\DFF_1514.D )
  );
  al_nand2ft _10287_ (
    .a(\DFF_1492.Q ),
    .b(\DFF_1514.Q ),
    .y(_04288_)
  );
  al_nand2ft _10288_ (
    .a(\DFF_1514.Q ),
    .b(\DFF_1492.Q ),
    .y(_04289_)
  );
  al_ao21ttf _10289_ (
    .a(_04288_),
    .b(_04289_),
    .c(\DFF_1535.Q ),
    .y(_04290_)
  );
  al_nand3ftt _10290_ (
    .a(\DFF_1535.Q ),
    .b(_04288_),
    .c(_04289_),
    .y(_04291_)
  );
  al_aoi21 _10291_ (
    .a(_04291_),
    .b(_04290_),
    .c(_00451_),
    .y(\DFF_1515.D )
  );
  al_oa21ftt _10292_ (
    .a(\DFF_1491.Q ),
    .b(\DFF_1515.Q ),
    .c(RESET),
    .y(_04292_)
  );
  al_aoi21ftf _10293_ (
    .a(\DFF_1491.Q ),
    .b(\DFF_1515.Q ),
    .c(_04292_),
    .y(\DFF_1516.D )
  );
  al_oa21ftt _10294_ (
    .a(\DFF_1490.Q ),
    .b(\DFF_1516.Q ),
    .c(RESET),
    .y(_04293_)
  );
  al_aoi21ftf _10295_ (
    .a(\DFF_1490.Q ),
    .b(\DFF_1516.Q ),
    .c(_04293_),
    .y(\DFF_1517.D )
  );
  al_oa21ftt _10296_ (
    .a(\DFF_1489.Q ),
    .b(\DFF_1517.Q ),
    .c(RESET),
    .y(_04294_)
  );
  al_aoi21ftf _10297_ (
    .a(\DFF_1489.Q ),
    .b(\DFF_1517.Q ),
    .c(_04294_),
    .y(\DFF_1518.D )
  );
  al_oa21ftt _10298_ (
    .a(\DFF_1488.Q ),
    .b(\DFF_1518.Q ),
    .c(RESET),
    .y(_04295_)
  );
  al_aoi21ftf _10299_ (
    .a(\DFF_1488.Q ),
    .b(\DFF_1518.Q ),
    .c(_04295_),
    .y(\DFF_1519.D )
  );
  al_nand2ft _10300_ (
    .a(\DFF_1487.Q ),
    .b(\DFF_1519.Q ),
    .y(_04296_)
  );
  al_nand2ft _10301_ (
    .a(\DFF_1519.Q ),
    .b(\DFF_1487.Q ),
    .y(_04297_)
  );
  al_ao21ttf _10302_ (
    .a(_04296_),
    .b(_04297_),
    .c(\DFF_1535.Q ),
    .y(_04298_)
  );
  al_nand3ftt _10303_ (
    .a(\DFF_1535.Q ),
    .b(_04296_),
    .c(_04297_),
    .y(_04299_)
  );
  al_aoi21 _10304_ (
    .a(_04299_),
    .b(_04298_),
    .c(_00451_),
    .y(\DFF_1520.D )
  );
  al_oa21ftt _10305_ (
    .a(\DFF_1486.Q ),
    .b(\DFF_1520.Q ),
    .c(RESET),
    .y(_04300_)
  );
  al_aoi21ftf _10306_ (
    .a(\DFF_1486.Q ),
    .b(\DFF_1520.Q ),
    .c(_04300_),
    .y(\DFF_1521.D )
  );
  al_oa21ftt _10307_ (
    .a(\DFF_1485.Q ),
    .b(\DFF_1521.Q ),
    .c(RESET),
    .y(_04301_)
  );
  al_aoi21ftf _10308_ (
    .a(\DFF_1485.Q ),
    .b(\DFF_1521.Q ),
    .c(_04301_),
    .y(\DFF_1522.D )
  );
  al_oa21ftt _10309_ (
    .a(\DFF_1484.Q ),
    .b(\DFF_1522.Q ),
    .c(RESET),
    .y(_04302_)
  );
  al_aoi21ftf _10310_ (
    .a(\DFF_1484.Q ),
    .b(\DFF_1522.Q ),
    .c(_04302_),
    .y(\DFF_1523.D )
  );
  al_oa21ftt _10311_ (
    .a(\DFF_1483.Q ),
    .b(\DFF_1523.Q ),
    .c(RESET),
    .y(_04303_)
  );
  al_aoi21ftf _10312_ (
    .a(\DFF_1483.Q ),
    .b(\DFF_1523.Q ),
    .c(_04303_),
    .y(\DFF_1524.D )
  );
  al_oa21ftt _10313_ (
    .a(\DFF_1482.Q ),
    .b(\DFF_1524.Q ),
    .c(RESET),
    .y(_04304_)
  );
  al_aoi21ftf _10314_ (
    .a(\DFF_1482.Q ),
    .b(\DFF_1524.Q ),
    .c(_04304_),
    .y(\DFF_1525.D )
  );
  al_oa21ftt _10315_ (
    .a(\DFF_1481.Q ),
    .b(\DFF_1525.Q ),
    .c(RESET),
    .y(_04305_)
  );
  al_aoi21ftf _10316_ (
    .a(\DFF_1481.Q ),
    .b(\DFF_1525.Q ),
    .c(_04305_),
    .y(\DFF_1526.D )
  );
  al_oa21ftt _10317_ (
    .a(\DFF_1480.Q ),
    .b(\DFF_1526.Q ),
    .c(RESET),
    .y(_04306_)
  );
  al_aoi21ftf _10318_ (
    .a(\DFF_1480.Q ),
    .b(\DFF_1526.Q ),
    .c(_04306_),
    .y(\DFF_1527.D )
  );
  al_oa21ftt _10319_ (
    .a(\DFF_1479.Q ),
    .b(\DFF_1527.Q ),
    .c(RESET),
    .y(_04307_)
  );
  al_aoi21ftf _10320_ (
    .a(\DFF_1479.Q ),
    .b(\DFF_1527.Q ),
    .c(_04307_),
    .y(\DFF_1528.D )
  );
  al_oa21ftt _10321_ (
    .a(\DFF_1478.Q ),
    .b(\DFF_1528.Q ),
    .c(RESET),
    .y(_04308_)
  );
  al_aoi21ftf _10322_ (
    .a(\DFF_1478.Q ),
    .b(\DFF_1528.Q ),
    .c(_04308_),
    .y(\DFF_1529.D )
  );
  al_oa21ftt _10323_ (
    .a(\DFF_1477.Q ),
    .b(\DFF_1529.Q ),
    .c(RESET),
    .y(_04309_)
  );
  al_aoi21ftf _10324_ (
    .a(\DFF_1477.Q ),
    .b(\DFF_1529.Q ),
    .c(_04309_),
    .y(\DFF_1530.D )
  );
  al_oa21ftt _10325_ (
    .a(\DFF_1476.Q ),
    .b(\DFF_1530.Q ),
    .c(RESET),
    .y(_04310_)
  );
  al_aoi21ftf _10326_ (
    .a(\DFF_1476.Q ),
    .b(\DFF_1530.Q ),
    .c(_04310_),
    .y(\DFF_1531.D )
  );
  al_oa21ftt _10327_ (
    .a(\DFF_1475.Q ),
    .b(\DFF_1531.Q ),
    .c(RESET),
    .y(_04311_)
  );
  al_aoi21ftf _10328_ (
    .a(\DFF_1475.Q ),
    .b(\DFF_1531.Q ),
    .c(_04311_),
    .y(\DFF_1532.D )
  );
  al_oa21ftt _10329_ (
    .a(\DFF_1474.Q ),
    .b(\DFF_1532.Q ),
    .c(RESET),
    .y(_04312_)
  );
  al_aoi21ftf _10330_ (
    .a(\DFF_1474.Q ),
    .b(\DFF_1532.Q ),
    .c(_04312_),
    .y(\DFF_1533.D )
  );
  al_oa21ftt _10331_ (
    .a(\DFF_1473.Q ),
    .b(\DFF_1533.Q ),
    .c(RESET),
    .y(_04313_)
  );
  al_aoi21ftf _10332_ (
    .a(\DFF_1473.Q ),
    .b(\DFF_1533.Q ),
    .c(_04313_),
    .y(\DFF_1534.D )
  );
  al_oa21ftt _10333_ (
    .a(\DFF_1472.Q ),
    .b(\DFF_1534.Q ),
    .c(RESET),
    .y(_04314_)
  );
  al_aoi21ftf _10334_ (
    .a(\DFF_1472.Q ),
    .b(\DFF_1534.Q ),
    .c(_04314_),
    .y(\DFF_1535.D )
  );
  al_and2 _10335_ (
    .a(RESET),
    .b(\DFF_1537.Q ),
    .y(\DFF_1536.D )
  );
  al_and2 _10336_ (
    .a(RESET),
    .b(\DFF_1538.Q ),
    .y(\DFF_1537.D )
  );
  al_and2 _10337_ (
    .a(RESET),
    .b(\DFF_1539.Q ),
    .y(\DFF_1538.D )
  );
  al_and2 _10338_ (
    .a(RESET),
    .b(\DFF_1540.Q ),
    .y(\DFF_1539.D )
  );
  al_and2 _10339_ (
    .a(RESET),
    .b(\DFF_1541.Q ),
    .y(\DFF_1540.D )
  );
  al_and2 _10340_ (
    .a(RESET),
    .b(\DFF_1542.Q ),
    .y(\DFF_1541.D )
  );
  al_and2 _10341_ (
    .a(RESET),
    .b(\DFF_1543.Q ),
    .y(\DFF_1542.D )
  );
  al_and2 _10342_ (
    .a(RESET),
    .b(\DFF_1544.Q ),
    .y(\DFF_1543.D )
  );
  al_and2 _10343_ (
    .a(RESET),
    .b(\DFF_1545.Q ),
    .y(\DFF_1544.D )
  );
  al_and2 _10344_ (
    .a(RESET),
    .b(\DFF_1546.Q ),
    .y(\DFF_1545.D )
  );
  al_and2 _10345_ (
    .a(RESET),
    .b(\DFF_1547.Q ),
    .y(\DFF_1546.D )
  );
  al_and2 _10346_ (
    .a(RESET),
    .b(\DFF_1548.Q ),
    .y(\DFF_1547.D )
  );
  al_and2 _10347_ (
    .a(RESET),
    .b(\DFF_1549.Q ),
    .y(\DFF_1548.D )
  );
  al_and2 _10348_ (
    .a(RESET),
    .b(\DFF_1550.Q ),
    .y(\DFF_1549.D )
  );
  al_and2 _10349_ (
    .a(RESET),
    .b(\DFF_1551.Q ),
    .y(\DFF_1550.D )
  );
  al_and2 _10350_ (
    .a(RESET),
    .b(\DFF_1552.Q ),
    .y(\DFF_1551.D )
  );
  al_and2 _10351_ (
    .a(RESET),
    .b(\DFF_1553.Q ),
    .y(\DFF_1552.D )
  );
  al_and2 _10352_ (
    .a(RESET),
    .b(\DFF_1554.Q ),
    .y(\DFF_1553.D )
  );
  al_and2 _10353_ (
    .a(RESET),
    .b(\DFF_1555.Q ),
    .y(\DFF_1554.D )
  );
  al_and2 _10354_ (
    .a(RESET),
    .b(\DFF_1556.Q ),
    .y(\DFF_1555.D )
  );
  al_and2 _10355_ (
    .a(RESET),
    .b(\DFF_1557.Q ),
    .y(\DFF_1556.D )
  );
  al_and2 _10356_ (
    .a(RESET),
    .b(\DFF_1558.Q ),
    .y(\DFF_1557.D )
  );
  al_and2 _10357_ (
    .a(RESET),
    .b(\DFF_1559.Q ),
    .y(\DFF_1558.D )
  );
  al_and2 _10358_ (
    .a(RESET),
    .b(\DFF_1560.Q ),
    .y(\DFF_1559.D )
  );
  al_and2 _10359_ (
    .a(RESET),
    .b(\DFF_1561.Q ),
    .y(\DFF_1560.D )
  );
  al_and2 _10360_ (
    .a(RESET),
    .b(\DFF_1562.Q ),
    .y(\DFF_1561.D )
  );
  al_and2 _10361_ (
    .a(RESET),
    .b(\DFF_1563.Q ),
    .y(\DFF_1562.D )
  );
  al_and2 _10362_ (
    .a(RESET),
    .b(\DFF_1564.Q ),
    .y(\DFF_1563.D )
  );
  al_and2 _10363_ (
    .a(RESET),
    .b(\DFF_1565.Q ),
    .y(\DFF_1564.D )
  );
  al_and2 _10364_ (
    .a(RESET),
    .b(\DFF_1566.Q ),
    .y(\DFF_1565.D )
  );
  al_and2 _10365_ (
    .a(RESET),
    .b(\DFF_1567.Q ),
    .y(\DFF_1566.D )
  );
  al_and2ft _10366_ (
    .a(\DFF_1536.Q ),
    .b(RESET),
    .y(\DFF_1567.D )
  );
  al_aoi21ttf _10367_ (
    .a(\DFF_1536.Q ),
    .b(TM0),
    .c(TM1),
    .y(_04315_)
  );
  al_mux2l _10368_ (
    .a(\DFF_1727.Q ),
    .b(DATA_0_31),
    .s(TM0),
    .y(_04316_)
  );
  al_oai21ttf _10369_ (
    .a(TM1),
    .b(_04316_),
    .c(_00451_),
    .y(_04317_)
  );
  al_aoi21 _10370_ (
    .a(_04315_),
    .b(_03853_),
    .c(_04317_),
    .y(\DFF_1568.D )
  );
  al_aoi21ttf _10371_ (
    .a(TM0),
    .b(\DFF_1537.Q ),
    .c(TM1),
    .y(_04318_)
  );
  al_mux2l _10372_ (
    .a(\DFF_1726.Q ),
    .b(DATA_0_30),
    .s(TM0),
    .y(_04319_)
  );
  al_oai21ttf _10373_ (
    .a(TM1),
    .b(_04319_),
    .c(_00451_),
    .y(_04320_)
  );
  al_aoi21 _10374_ (
    .a(_04318_),
    .b(_03869_),
    .c(_04320_),
    .y(\DFF_1569.D )
  );
  al_aoi21ttf _10375_ (
    .a(TM0),
    .b(\DFF_1538.Q ),
    .c(TM1),
    .y(_04321_)
  );
  al_mux2l _10376_ (
    .a(\DFF_1725.Q ),
    .b(DATA_0_29),
    .s(TM0),
    .y(_04322_)
  );
  al_oai21ttf _10377_ (
    .a(TM1),
    .b(_04322_),
    .c(_00451_),
    .y(_04323_)
  );
  al_aoi21 _10378_ (
    .a(_04321_),
    .b(_03885_),
    .c(_04323_),
    .y(\DFF_1570.D )
  );
  al_aoi21ttf _10379_ (
    .a(TM0),
    .b(\DFF_1539.Q ),
    .c(TM1),
    .y(_04324_)
  );
  al_mux2l _10380_ (
    .a(\DFF_1724.Q ),
    .b(DATA_0_28),
    .s(TM0),
    .y(_04325_)
  );
  al_oai21ttf _10381_ (
    .a(TM1),
    .b(_04325_),
    .c(_00451_),
    .y(_04326_)
  );
  al_aoi21 _10382_ (
    .a(_04324_),
    .b(_03901_),
    .c(_04326_),
    .y(\DFF_1571.D )
  );
  al_aoi21ttf _10383_ (
    .a(TM0),
    .b(\DFF_1540.Q ),
    .c(TM1),
    .y(_04327_)
  );
  al_mux2l _10384_ (
    .a(\DFF_1723.Q ),
    .b(DATA_0_27),
    .s(TM0),
    .y(_04328_)
  );
  al_oai21ttf _10385_ (
    .a(TM1),
    .b(_04328_),
    .c(_00451_),
    .y(_04329_)
  );
  al_aoi21 _10386_ (
    .a(_04327_),
    .b(_03917_),
    .c(_04329_),
    .y(\DFF_1572.D )
  );
  al_aoi21ttf _10387_ (
    .a(TM0),
    .b(\DFF_1541.Q ),
    .c(TM1),
    .y(_04330_)
  );
  al_mux2l _10388_ (
    .a(\DFF_1722.Q ),
    .b(DATA_0_26),
    .s(TM0),
    .y(_04331_)
  );
  al_oai21ttf _10389_ (
    .a(TM1),
    .b(_04331_),
    .c(_00451_),
    .y(_04332_)
  );
  al_aoi21 _10390_ (
    .a(_04330_),
    .b(_03933_),
    .c(_04332_),
    .y(\DFF_1573.D )
  );
  al_aoi21ttf _10391_ (
    .a(TM0),
    .b(\DFF_1542.Q ),
    .c(TM1),
    .y(_04333_)
  );
  al_mux2l _10392_ (
    .a(\DFF_1721.Q ),
    .b(DATA_0_25),
    .s(TM0),
    .y(_04334_)
  );
  al_oai21ttf _10393_ (
    .a(TM1),
    .b(_04334_),
    .c(_00451_),
    .y(_04335_)
  );
  al_aoi21 _10394_ (
    .a(_04333_),
    .b(_03949_),
    .c(_04335_),
    .y(\DFF_1574.D )
  );
  al_aoi21ttf _10395_ (
    .a(TM0),
    .b(\DFF_1543.Q ),
    .c(TM1),
    .y(_04336_)
  );
  al_mux2l _10396_ (
    .a(\DFF_1720.Q ),
    .b(DATA_0_24),
    .s(TM0),
    .y(_04337_)
  );
  al_oai21ttf _10397_ (
    .a(TM1),
    .b(_04337_),
    .c(_00451_),
    .y(_04338_)
  );
  al_aoi21 _10398_ (
    .a(_04336_),
    .b(_03965_),
    .c(_04338_),
    .y(\DFF_1575.D )
  );
  al_aoi21ttf _10399_ (
    .a(TM0),
    .b(\DFF_1544.Q ),
    .c(TM1),
    .y(_04339_)
  );
  al_mux2l _10400_ (
    .a(\DFF_1719.Q ),
    .b(DATA_0_23),
    .s(TM0),
    .y(_04340_)
  );
  al_oai21ttf _10401_ (
    .a(TM1),
    .b(_04340_),
    .c(_00451_),
    .y(_04341_)
  );
  al_aoi21 _10402_ (
    .a(_04339_),
    .b(_03981_),
    .c(_04341_),
    .y(\DFF_1576.D )
  );
  al_aoi21ttf _10403_ (
    .a(TM0),
    .b(\DFF_1545.Q ),
    .c(TM1),
    .y(_04342_)
  );
  al_mux2l _10404_ (
    .a(\DFF_1718.Q ),
    .b(DATA_0_22),
    .s(TM0),
    .y(_04343_)
  );
  al_oai21ttf _10405_ (
    .a(TM1),
    .b(_04343_),
    .c(_00451_),
    .y(_04344_)
  );
  al_aoi21 _10406_ (
    .a(_04342_),
    .b(_03997_),
    .c(_04344_),
    .y(\DFF_1577.D )
  );
  al_aoi21ttf _10407_ (
    .a(TM0),
    .b(\DFF_1546.Q ),
    .c(TM1),
    .y(_04345_)
  );
  al_mux2l _10408_ (
    .a(\DFF_1717.Q ),
    .b(DATA_0_21),
    .s(TM0),
    .y(_04346_)
  );
  al_oai21ttf _10409_ (
    .a(TM1),
    .b(_04346_),
    .c(_00451_),
    .y(_04347_)
  );
  al_aoi21 _10410_ (
    .a(_04345_),
    .b(_04013_),
    .c(_04347_),
    .y(\DFF_1578.D )
  );
  al_aoi21ttf _10411_ (
    .a(TM0),
    .b(\DFF_1547.Q ),
    .c(TM1),
    .y(_04348_)
  );
  al_mux2l _10412_ (
    .a(\DFF_1716.Q ),
    .b(DATA_0_20),
    .s(TM0),
    .y(_04349_)
  );
  al_oai21ttf _10413_ (
    .a(TM1),
    .b(_04349_),
    .c(_00451_),
    .y(_04350_)
  );
  al_aoi21 _10414_ (
    .a(_04348_),
    .b(_04029_),
    .c(_04350_),
    .y(\DFF_1579.D )
  );
  al_aoi21ttf _10415_ (
    .a(TM0),
    .b(\DFF_1548.Q ),
    .c(TM1),
    .y(_04351_)
  );
  al_mux2l _10416_ (
    .a(\DFF_1715.Q ),
    .b(DATA_0_19),
    .s(TM0),
    .y(_04352_)
  );
  al_oai21ttf _10417_ (
    .a(TM1),
    .b(_04352_),
    .c(_00451_),
    .y(_04353_)
  );
  al_aoi21 _10418_ (
    .a(_04351_),
    .b(_04045_),
    .c(_04353_),
    .y(\DFF_1580.D )
  );
  al_aoi21ttf _10419_ (
    .a(TM0),
    .b(\DFF_1549.Q ),
    .c(TM1),
    .y(_04354_)
  );
  al_mux2l _10420_ (
    .a(\DFF_1714.Q ),
    .b(DATA_0_18),
    .s(TM0),
    .y(_04355_)
  );
  al_oai21ttf _10421_ (
    .a(TM1),
    .b(_04355_),
    .c(_00451_),
    .y(_04356_)
  );
  al_aoi21 _10422_ (
    .a(_04354_),
    .b(_04061_),
    .c(_04356_),
    .y(\DFF_1581.D )
  );
  al_aoi21ttf _10423_ (
    .a(TM0),
    .b(\DFF_1550.Q ),
    .c(TM1),
    .y(_04357_)
  );
  al_mux2l _10424_ (
    .a(\DFF_1713.Q ),
    .b(DATA_0_17),
    .s(TM0),
    .y(_04358_)
  );
  al_oai21ttf _10425_ (
    .a(TM1),
    .b(_04358_),
    .c(_00451_),
    .y(_04359_)
  );
  al_aoi21 _10426_ (
    .a(_04357_),
    .b(_04077_),
    .c(_04359_),
    .y(\DFF_1582.D )
  );
  al_aoi21ttf _10427_ (
    .a(TM0),
    .b(\DFF_1551.Q ),
    .c(TM1),
    .y(_04360_)
  );
  al_mux2l _10428_ (
    .a(\DFF_1712.Q ),
    .b(DATA_0_16),
    .s(TM0),
    .y(_04361_)
  );
  al_oai21ttf _10429_ (
    .a(TM1),
    .b(_04361_),
    .c(_00451_),
    .y(_04362_)
  );
  al_aoi21 _10430_ (
    .a(_04360_),
    .b(_04093_),
    .c(_04362_),
    .y(\DFF_1583.D )
  );
  al_aoi21ttf _10431_ (
    .a(TM0),
    .b(\DFF_1552.Q ),
    .c(TM1),
    .y(_04363_)
  );
  al_mux2l _10432_ (
    .a(\DFF_1711.Q ),
    .b(DATA_0_15),
    .s(TM0),
    .y(_04364_)
  );
  al_oai21ttf _10433_ (
    .a(TM1),
    .b(_04364_),
    .c(_00451_),
    .y(_04365_)
  );
  al_aoi21 _10434_ (
    .a(_04363_),
    .b(_04106_),
    .c(_04365_),
    .y(\DFF_1584.D )
  );
  al_aoi21ttf _10435_ (
    .a(TM0),
    .b(\DFF_1553.Q ),
    .c(TM1),
    .y(_04366_)
  );
  al_mux2l _10436_ (
    .a(\DFF_1710.Q ),
    .b(DATA_0_14),
    .s(TM0),
    .y(_04367_)
  );
  al_oai21ttf _10437_ (
    .a(TM1),
    .b(_04367_),
    .c(_00451_),
    .y(_04368_)
  );
  al_aoi21 _10438_ (
    .a(_04366_),
    .b(_04117_),
    .c(_04368_),
    .y(\DFF_1585.D )
  );
  al_aoi21ttf _10439_ (
    .a(TM0),
    .b(\DFF_1554.Q ),
    .c(TM1),
    .y(_04369_)
  );
  al_mux2l _10440_ (
    .a(\DFF_1709.Q ),
    .b(DATA_0_13),
    .s(TM0),
    .y(_04370_)
  );
  al_oai21ttf _10441_ (
    .a(TM1),
    .b(_04370_),
    .c(_00451_),
    .y(_04371_)
  );
  al_aoi21 _10442_ (
    .a(_04369_),
    .b(_04128_),
    .c(_04371_),
    .y(\DFF_1586.D )
  );
  al_aoi21ttf _10443_ (
    .a(TM0),
    .b(\DFF_1555.Q ),
    .c(TM1),
    .y(_04372_)
  );
  al_mux2l _10444_ (
    .a(\DFF_1708.Q ),
    .b(DATA_0_12),
    .s(TM0),
    .y(_04373_)
  );
  al_oai21ttf _10445_ (
    .a(TM1),
    .b(_04373_),
    .c(_00451_),
    .y(_04374_)
  );
  al_aoi21 _10446_ (
    .a(_04372_),
    .b(_04139_),
    .c(_04374_),
    .y(\DFF_1587.D )
  );
  al_aoi21ttf _10447_ (
    .a(TM0),
    .b(\DFF_1556.Q ),
    .c(TM1),
    .y(_04375_)
  );
  al_mux2l _10448_ (
    .a(\DFF_1707.Q ),
    .b(DATA_0_11),
    .s(TM0),
    .y(_04376_)
  );
  al_oai21ttf _10449_ (
    .a(TM1),
    .b(_04376_),
    .c(_00451_),
    .y(_04377_)
  );
  al_aoi21 _10450_ (
    .a(_04375_),
    .b(_04150_),
    .c(_04377_),
    .y(\DFF_1588.D )
  );
  al_aoi21ttf _10451_ (
    .a(TM0),
    .b(\DFF_1557.Q ),
    .c(TM1),
    .y(_04378_)
  );
  al_mux2l _10452_ (
    .a(\DFF_1706.Q ),
    .b(DATA_0_10),
    .s(TM0),
    .y(_04379_)
  );
  al_oai21ttf _10453_ (
    .a(TM1),
    .b(_04379_),
    .c(_00451_),
    .y(_04380_)
  );
  al_aoi21 _10454_ (
    .a(_04378_),
    .b(_04161_),
    .c(_04380_),
    .y(\DFF_1589.D )
  );
  al_aoi21ttf _10455_ (
    .a(TM0),
    .b(\DFF_1558.Q ),
    .c(TM1),
    .y(_04381_)
  );
  al_mux2l _10456_ (
    .a(\DFF_1705.Q ),
    .b(DATA_0_9),
    .s(TM0),
    .y(_04382_)
  );
  al_oai21ttf _10457_ (
    .a(TM1),
    .b(_04382_),
    .c(_00451_),
    .y(_04383_)
  );
  al_aoi21 _10458_ (
    .a(_04381_),
    .b(_04172_),
    .c(_04383_),
    .y(\DFF_1590.D )
  );
  al_aoi21ttf _10459_ (
    .a(TM0),
    .b(\DFF_1559.Q ),
    .c(TM1),
    .y(_04384_)
  );
  al_mux2l _10460_ (
    .a(\DFF_1704.Q ),
    .b(DATA_0_8),
    .s(TM0),
    .y(_04385_)
  );
  al_oai21ttf _10461_ (
    .a(TM1),
    .b(_04385_),
    .c(_00451_),
    .y(_04386_)
  );
  al_aoi21 _10462_ (
    .a(_04384_),
    .b(_04183_),
    .c(_04386_),
    .y(\DFF_1591.D )
  );
  al_aoi21ttf _10463_ (
    .a(TM0),
    .b(\DFF_1560.Q ),
    .c(TM1),
    .y(_04387_)
  );
  al_mux2l _10464_ (
    .a(\DFF_1703.Q ),
    .b(DATA_0_7),
    .s(TM0),
    .y(_04388_)
  );
  al_oai21ttf _10465_ (
    .a(TM1),
    .b(_04388_),
    .c(_00451_),
    .y(_04389_)
  );
  al_aoi21 _10466_ (
    .a(_04387_),
    .b(_04194_),
    .c(_04389_),
    .y(\DFF_1592.D )
  );
  al_aoi21ttf _10467_ (
    .a(TM0),
    .b(\DFF_1561.Q ),
    .c(TM1),
    .y(_04390_)
  );
  al_mux2l _10468_ (
    .a(\DFF_1702.Q ),
    .b(DATA_0_6),
    .s(TM0),
    .y(_04391_)
  );
  al_oai21ttf _10469_ (
    .a(TM1),
    .b(_04391_),
    .c(_00451_),
    .y(_04392_)
  );
  al_aoi21 _10470_ (
    .a(_04390_),
    .b(_04205_),
    .c(_04392_),
    .y(\DFF_1593.D )
  );
  al_aoi21ttf _10471_ (
    .a(TM0),
    .b(\DFF_1562.Q ),
    .c(TM1),
    .y(_04393_)
  );
  al_mux2l _10472_ (
    .a(\DFF_1701.Q ),
    .b(DATA_0_5),
    .s(TM0),
    .y(_04394_)
  );
  al_oai21ttf _10473_ (
    .a(TM1),
    .b(_04394_),
    .c(_00451_),
    .y(_04395_)
  );
  al_aoi21 _10474_ (
    .a(_04393_),
    .b(_04216_),
    .c(_04395_),
    .y(\DFF_1594.D )
  );
  al_aoi21ttf _10475_ (
    .a(TM0),
    .b(\DFF_1563.Q ),
    .c(TM1),
    .y(_04396_)
  );
  al_mux2l _10476_ (
    .a(\DFF_1700.Q ),
    .b(DATA_0_4),
    .s(TM0),
    .y(_04397_)
  );
  al_oai21ttf _10477_ (
    .a(TM1),
    .b(_04397_),
    .c(_00451_),
    .y(_04398_)
  );
  al_aoi21 _10478_ (
    .a(_04396_),
    .b(_04227_),
    .c(_04398_),
    .y(\DFF_1595.D )
  );
  al_aoi21ttf _10479_ (
    .a(TM0),
    .b(\DFF_1564.Q ),
    .c(TM1),
    .y(_04399_)
  );
  al_mux2l _10480_ (
    .a(\DFF_1699.Q ),
    .b(DATA_0_3),
    .s(TM0),
    .y(_04400_)
  );
  al_oai21ttf _10481_ (
    .a(TM1),
    .b(_04400_),
    .c(_00451_),
    .y(_04401_)
  );
  al_aoi21 _10482_ (
    .a(_04399_),
    .b(_04238_),
    .c(_04401_),
    .y(\DFF_1596.D )
  );
  al_aoi21ttf _10483_ (
    .a(TM0),
    .b(\DFF_1565.Q ),
    .c(TM1),
    .y(_04402_)
  );
  al_mux2l _10484_ (
    .a(\DFF_1698.Q ),
    .b(DATA_0_2),
    .s(TM0),
    .y(_04403_)
  );
  al_oai21ttf _10485_ (
    .a(TM1),
    .b(_04403_),
    .c(_00451_),
    .y(_04404_)
  );
  al_aoi21 _10486_ (
    .a(_04402_),
    .b(_04249_),
    .c(_04404_),
    .y(\DFF_1597.D )
  );
  al_aoi21ttf _10487_ (
    .a(TM0),
    .b(\DFF_1566.Q ),
    .c(TM1),
    .y(_04405_)
  );
  al_mux2l _10488_ (
    .a(\DFF_1697.Q ),
    .b(DATA_0_1),
    .s(TM0),
    .y(_04406_)
  );
  al_oai21ttf _10489_ (
    .a(TM1),
    .b(_04406_),
    .c(_00451_),
    .y(_04407_)
  );
  al_aoi21 _10490_ (
    .a(_04405_),
    .b(_04260_),
    .c(_04407_),
    .y(\DFF_1598.D )
  );
  al_aoi21ttf _10491_ (
    .a(TM0),
    .b(\DFF_1567.Q ),
    .c(TM1),
    .y(_04408_)
  );
  al_mux2l _10492_ (
    .a(\DFF_1696.Q ),
    .b(DATA_0_0),
    .s(TM0),
    .y(_04409_)
  );
  al_oai21ttf _10493_ (
    .a(TM1),
    .b(_04409_),
    .c(_00451_),
    .y(_04410_)
  );
  al_aoi21 _10494_ (
    .a(_04408_),
    .b(_04271_),
    .c(_04410_),
    .y(\DFF_1599.D )
  );
  al_and2 _10495_ (
    .a(RESET),
    .b(\DFF_1568.Q ),
    .y(\DFF_1600.D )
  );
  al_and2 _10496_ (
    .a(RESET),
    .b(\DFF_1569.Q ),
    .y(\DFF_1601.D )
  );
  al_and2 _10497_ (
    .a(RESET),
    .b(\DFF_1570.Q ),
    .y(\DFF_1602.D )
  );
  al_and2 _10498_ (
    .a(RESET),
    .b(\DFF_1571.Q ),
    .y(\DFF_1603.D )
  );
  al_and2 _10499_ (
    .a(RESET),
    .b(\DFF_1572.Q ),
    .y(\DFF_1604.D )
  );
  al_and2 _10500_ (
    .a(RESET),
    .b(\DFF_1573.Q ),
    .y(\DFF_1605.D )
  );
  al_and2 _10501_ (
    .a(RESET),
    .b(\DFF_1574.Q ),
    .y(\DFF_1606.D )
  );
  al_and2 _10502_ (
    .a(RESET),
    .b(\DFF_1575.Q ),
    .y(\DFF_1607.D )
  );
  al_and2 _10503_ (
    .a(RESET),
    .b(\DFF_1576.Q ),
    .y(\DFF_1608.D )
  );
  al_and2 _10504_ (
    .a(RESET),
    .b(\DFF_1577.Q ),
    .y(\DFF_1609.D )
  );
  al_and2 _10505_ (
    .a(RESET),
    .b(\DFF_1578.Q ),
    .y(\DFF_1610.D )
  );
  al_and2 _10506_ (
    .a(RESET),
    .b(\DFF_1579.Q ),
    .y(\DFF_1611.D )
  );
  al_and2 _10507_ (
    .a(RESET),
    .b(\DFF_1580.Q ),
    .y(\DFF_1612.D )
  );
  al_and2 _10508_ (
    .a(RESET),
    .b(\DFF_1581.Q ),
    .y(\DFF_1613.D )
  );
  al_and2 _10509_ (
    .a(RESET),
    .b(\DFF_1582.Q ),
    .y(\DFF_1614.D )
  );
  al_and2 _10510_ (
    .a(RESET),
    .b(\DFF_1583.Q ),
    .y(\DFF_1615.D )
  );
  al_and2 _10511_ (
    .a(RESET),
    .b(\DFF_1584.Q ),
    .y(\DFF_1616.D )
  );
  al_and2 _10512_ (
    .a(RESET),
    .b(\DFF_1585.Q ),
    .y(\DFF_1617.D )
  );
  al_and2 _10513_ (
    .a(RESET),
    .b(\DFF_1586.Q ),
    .y(\DFF_1618.D )
  );
  al_and2 _10514_ (
    .a(RESET),
    .b(\DFF_1587.Q ),
    .y(\DFF_1619.D )
  );
  al_and2 _10515_ (
    .a(RESET),
    .b(\DFF_1588.Q ),
    .y(\DFF_1620.D )
  );
  al_and2 _10516_ (
    .a(RESET),
    .b(\DFF_1589.Q ),
    .y(\DFF_1621.D )
  );
  al_and2 _10517_ (
    .a(RESET),
    .b(\DFF_1590.Q ),
    .y(\DFF_1622.D )
  );
  al_and2 _10518_ (
    .a(RESET),
    .b(\DFF_1591.Q ),
    .y(\DFF_1623.D )
  );
  al_and2 _10519_ (
    .a(RESET),
    .b(\DFF_1592.Q ),
    .y(\DFF_1624.D )
  );
  al_and2 _10520_ (
    .a(RESET),
    .b(\DFF_1593.Q ),
    .y(\DFF_1625.D )
  );
  al_and2 _10521_ (
    .a(RESET),
    .b(\DFF_1594.Q ),
    .y(\DFF_1626.D )
  );
  al_and2 _10522_ (
    .a(RESET),
    .b(\DFF_1595.Q ),
    .y(\DFF_1627.D )
  );
  al_and2 _10523_ (
    .a(RESET),
    .b(\DFF_1596.Q ),
    .y(\DFF_1628.D )
  );
  al_and2 _10524_ (
    .a(RESET),
    .b(\DFF_1597.Q ),
    .y(\DFF_1629.D )
  );
  al_and2 _10525_ (
    .a(RESET),
    .b(\DFF_1598.Q ),
    .y(\DFF_1630.D )
  );
  al_and2 _10526_ (
    .a(RESET),
    .b(\DFF_1599.Q ),
    .y(\DFF_1631.D )
  );
  al_and2 _10527_ (
    .a(RESET),
    .b(\DFF_1600.Q ),
    .y(\DFF_1632.D )
  );
  al_and2 _10528_ (
    .a(RESET),
    .b(\DFF_1601.Q ),
    .y(\DFF_1633.D )
  );
  al_and2 _10529_ (
    .a(RESET),
    .b(\DFF_1602.Q ),
    .y(\DFF_1634.D )
  );
  al_and2 _10530_ (
    .a(RESET),
    .b(\DFF_1603.Q ),
    .y(\DFF_1635.D )
  );
  al_and2 _10531_ (
    .a(RESET),
    .b(\DFF_1604.Q ),
    .y(\DFF_1636.D )
  );
  al_and2 _10532_ (
    .a(RESET),
    .b(\DFF_1605.Q ),
    .y(\DFF_1637.D )
  );
  al_and2 _10533_ (
    .a(RESET),
    .b(\DFF_1606.Q ),
    .y(\DFF_1638.D )
  );
  al_and2 _10534_ (
    .a(RESET),
    .b(\DFF_1607.Q ),
    .y(\DFF_1639.D )
  );
  al_and2 _10535_ (
    .a(RESET),
    .b(\DFF_1608.Q ),
    .y(\DFF_1640.D )
  );
  al_and2 _10536_ (
    .a(RESET),
    .b(\DFF_1609.Q ),
    .y(\DFF_1641.D )
  );
  al_and2 _10537_ (
    .a(RESET),
    .b(\DFF_1610.Q ),
    .y(\DFF_1642.D )
  );
  al_and2 _10538_ (
    .a(RESET),
    .b(\DFF_1611.Q ),
    .y(\DFF_1643.D )
  );
  al_and2 _10539_ (
    .a(RESET),
    .b(\DFF_1612.Q ),
    .y(\DFF_1644.D )
  );
  al_and2 _10540_ (
    .a(RESET),
    .b(\DFF_1613.Q ),
    .y(\DFF_1645.D )
  );
  al_and2 _10541_ (
    .a(RESET),
    .b(\DFF_1614.Q ),
    .y(\DFF_1646.D )
  );
  al_and2 _10542_ (
    .a(RESET),
    .b(\DFF_1615.Q ),
    .y(\DFF_1647.D )
  );
  al_and2 _10543_ (
    .a(RESET),
    .b(\DFF_1616.Q ),
    .y(\DFF_1648.D )
  );
  al_and2 _10544_ (
    .a(RESET),
    .b(\DFF_1617.Q ),
    .y(\DFF_1649.D )
  );
  al_and2 _10545_ (
    .a(RESET),
    .b(\DFF_1618.Q ),
    .y(\DFF_1650.D )
  );
  al_and2 _10546_ (
    .a(RESET),
    .b(\DFF_1619.Q ),
    .y(\DFF_1651.D )
  );
  al_and2 _10547_ (
    .a(RESET),
    .b(\DFF_1620.Q ),
    .y(\DFF_1652.D )
  );
  al_and2 _10548_ (
    .a(RESET),
    .b(\DFF_1621.Q ),
    .y(\DFF_1653.D )
  );
  al_and2 _10549_ (
    .a(RESET),
    .b(\DFF_1622.Q ),
    .y(\DFF_1654.D )
  );
  al_and2 _10550_ (
    .a(RESET),
    .b(\DFF_1623.Q ),
    .y(\DFF_1655.D )
  );
  al_and2 _10551_ (
    .a(RESET),
    .b(\DFF_1624.Q ),
    .y(\DFF_1656.D )
  );
  al_and2 _10552_ (
    .a(RESET),
    .b(\DFF_1625.Q ),
    .y(\DFF_1657.D )
  );
  al_and2 _10553_ (
    .a(RESET),
    .b(\DFF_1626.Q ),
    .y(\DFF_1658.D )
  );
  al_and2 _10554_ (
    .a(RESET),
    .b(\DFF_1627.Q ),
    .y(\DFF_1659.D )
  );
  al_and2 _10555_ (
    .a(RESET),
    .b(\DFF_1628.Q ),
    .y(\DFF_1660.D )
  );
  al_and2 _10556_ (
    .a(RESET),
    .b(\DFF_1629.Q ),
    .y(\DFF_1661.D )
  );
  al_and2 _10557_ (
    .a(RESET),
    .b(\DFF_1630.Q ),
    .y(\DFF_1662.D )
  );
  al_and2 _10558_ (
    .a(RESET),
    .b(\DFF_1631.Q ),
    .y(\DFF_1663.D )
  );
  al_and2 _10559_ (
    .a(RESET),
    .b(\DFF_1632.Q ),
    .y(\DFF_1664.D )
  );
  al_and2 _10560_ (
    .a(RESET),
    .b(\DFF_1633.Q ),
    .y(\DFF_1665.D )
  );
  al_and2 _10561_ (
    .a(RESET),
    .b(\DFF_1634.Q ),
    .y(\DFF_1666.D )
  );
  al_and2 _10562_ (
    .a(RESET),
    .b(\DFF_1635.Q ),
    .y(\DFF_1667.D )
  );
  al_and2 _10563_ (
    .a(RESET),
    .b(\DFF_1636.Q ),
    .y(\DFF_1668.D )
  );
  al_and2 _10564_ (
    .a(RESET),
    .b(\DFF_1637.Q ),
    .y(\DFF_1669.D )
  );
  al_and2 _10565_ (
    .a(RESET),
    .b(\DFF_1638.Q ),
    .y(\DFF_1670.D )
  );
  al_and2 _10566_ (
    .a(RESET),
    .b(\DFF_1639.Q ),
    .y(\DFF_1671.D )
  );
  al_and2 _10567_ (
    .a(RESET),
    .b(\DFF_1640.Q ),
    .y(\DFF_1672.D )
  );
  al_and2 _10568_ (
    .a(RESET),
    .b(\DFF_1641.Q ),
    .y(\DFF_1673.D )
  );
  al_and2 _10569_ (
    .a(RESET),
    .b(\DFF_1642.Q ),
    .y(\DFF_1674.D )
  );
  al_and2 _10570_ (
    .a(RESET),
    .b(\DFF_1643.Q ),
    .y(\DFF_1675.D )
  );
  al_and2 _10571_ (
    .a(RESET),
    .b(\DFF_1644.Q ),
    .y(\DFF_1676.D )
  );
  al_and2 _10572_ (
    .a(RESET),
    .b(\DFF_1645.Q ),
    .y(\DFF_1677.D )
  );
  al_and2 _10573_ (
    .a(RESET),
    .b(\DFF_1646.Q ),
    .y(\DFF_1678.D )
  );
  al_and2 _10574_ (
    .a(RESET),
    .b(\DFF_1647.Q ),
    .y(\DFF_1679.D )
  );
  al_and2 _10575_ (
    .a(RESET),
    .b(\DFF_1648.Q ),
    .y(\DFF_1680.D )
  );
  al_and2 _10576_ (
    .a(RESET),
    .b(\DFF_1649.Q ),
    .y(\DFF_1681.D )
  );
  al_and2 _10577_ (
    .a(RESET),
    .b(\DFF_1650.Q ),
    .y(\DFF_1682.D )
  );
  al_and2 _10578_ (
    .a(RESET),
    .b(\DFF_1651.Q ),
    .y(\DFF_1683.D )
  );
  al_and2 _10579_ (
    .a(RESET),
    .b(\DFF_1652.Q ),
    .y(\DFF_1684.D )
  );
  al_and2 _10580_ (
    .a(RESET),
    .b(\DFF_1653.Q ),
    .y(\DFF_1685.D )
  );
  al_and2 _10581_ (
    .a(RESET),
    .b(\DFF_1654.Q ),
    .y(\DFF_1686.D )
  );
  al_and2 _10582_ (
    .a(RESET),
    .b(\DFF_1655.Q ),
    .y(\DFF_1687.D )
  );
  al_and2 _10583_ (
    .a(RESET),
    .b(\DFF_1656.Q ),
    .y(\DFF_1688.D )
  );
  al_and2 _10584_ (
    .a(RESET),
    .b(\DFF_1657.Q ),
    .y(\DFF_1689.D )
  );
  al_and2 _10585_ (
    .a(RESET),
    .b(\DFF_1658.Q ),
    .y(\DFF_1690.D )
  );
  al_and2 _10586_ (
    .a(RESET),
    .b(\DFF_1659.Q ),
    .y(\DFF_1691.D )
  );
  al_and2 _10587_ (
    .a(RESET),
    .b(\DFF_1660.Q ),
    .y(\DFF_1692.D )
  );
  al_and2 _10588_ (
    .a(RESET),
    .b(\DFF_1661.Q ),
    .y(\DFF_1693.D )
  );
  al_and2 _10589_ (
    .a(RESET),
    .b(\DFF_1662.Q ),
    .y(\DFF_1694.D )
  );
  al_and2 _10590_ (
    .a(RESET),
    .b(\DFF_1663.Q ),
    .y(\DFF_1695.D )
  );
  al_oa21ftt _10591_ (
    .a(\DFF_1695.Q ),
    .b(\DFF_1727.Q ),
    .c(RESET),
    .y(_04411_)
  );
  al_aoi21ftf _10592_ (
    .a(\DFF_1695.Q ),
    .b(\DFF_1727.Q ),
    .c(_04411_),
    .y(\DFF_1696.D )
  );
  al_oa21ftt _10593_ (
    .a(\DFF_1694.Q ),
    .b(\DFF_1696.Q ),
    .c(RESET),
    .y(_04412_)
  );
  al_aoi21ftf _10594_ (
    .a(\DFF_1694.Q ),
    .b(\DFF_1696.Q ),
    .c(_04412_),
    .y(\DFF_1697.D )
  );
  al_oa21ftt _10595_ (
    .a(\DFF_1693.Q ),
    .b(\DFF_1697.Q ),
    .c(RESET),
    .y(_04413_)
  );
  al_aoi21ftf _10596_ (
    .a(\DFF_1693.Q ),
    .b(\DFF_1697.Q ),
    .c(_04413_),
    .y(\DFF_1698.D )
  );
  al_oa21ftt _10597_ (
    .a(\DFF_1692.Q ),
    .b(\DFF_1698.Q ),
    .c(RESET),
    .y(_04414_)
  );
  al_aoi21ftf _10598_ (
    .a(\DFF_1692.Q ),
    .b(\DFF_1698.Q ),
    .c(_04414_),
    .y(\DFF_1699.D )
  );
  al_nand2ft _10599_ (
    .a(\DFF_1691.Q ),
    .b(\DFF_1699.Q ),
    .y(_04415_)
  );
  al_nand2ft _10600_ (
    .a(\DFF_1699.Q ),
    .b(\DFF_1691.Q ),
    .y(_04416_)
  );
  al_ao21ttf _10601_ (
    .a(_04415_),
    .b(_04416_),
    .c(\DFF_1727.Q ),
    .y(_04417_)
  );
  al_nand3ftt _10602_ (
    .a(\DFF_1727.Q ),
    .b(_04415_),
    .c(_04416_),
    .y(_04418_)
  );
  al_aoi21 _10603_ (
    .a(_04418_),
    .b(_04417_),
    .c(_00451_),
    .y(\DFF_1700.D )
  );
  al_oa21ftt _10604_ (
    .a(\DFF_1690.Q ),
    .b(\DFF_1700.Q ),
    .c(RESET),
    .y(_04419_)
  );
  al_aoi21ftf _10605_ (
    .a(\DFF_1690.Q ),
    .b(\DFF_1700.Q ),
    .c(_04419_),
    .y(\DFF_1701.D )
  );
  al_oa21ftt _10606_ (
    .a(\DFF_1689.Q ),
    .b(\DFF_1701.Q ),
    .c(RESET),
    .y(_04420_)
  );
  al_aoi21ftf _10607_ (
    .a(\DFF_1689.Q ),
    .b(\DFF_1701.Q ),
    .c(_04420_),
    .y(\DFF_1702.D )
  );
  al_oa21ftt _10608_ (
    .a(\DFF_1688.Q ),
    .b(\DFF_1702.Q ),
    .c(RESET),
    .y(_04421_)
  );
  al_aoi21ftf _10609_ (
    .a(\DFF_1688.Q ),
    .b(\DFF_1702.Q ),
    .c(_04421_),
    .y(\DFF_1703.D )
  );
  al_oa21ftt _10610_ (
    .a(\DFF_1687.Q ),
    .b(\DFF_1703.Q ),
    .c(RESET),
    .y(_04422_)
  );
  al_aoi21ftf _10611_ (
    .a(\DFF_1687.Q ),
    .b(\DFF_1703.Q ),
    .c(_04422_),
    .y(\DFF_1704.D )
  );
  al_oa21ftt _10612_ (
    .a(\DFF_1686.Q ),
    .b(\DFF_1704.Q ),
    .c(RESET),
    .y(_04423_)
  );
  al_aoi21ftf _10613_ (
    .a(\DFF_1686.Q ),
    .b(\DFF_1704.Q ),
    .c(_04423_),
    .y(\DFF_1705.D )
  );
  al_oa21ftt _10614_ (
    .a(\DFF_1685.Q ),
    .b(\DFF_1705.Q ),
    .c(RESET),
    .y(_04424_)
  );
  al_aoi21ftf _10615_ (
    .a(\DFF_1685.Q ),
    .b(\DFF_1705.Q ),
    .c(_04424_),
    .y(\DFF_1706.D )
  );
  al_nand2ft _10616_ (
    .a(\DFF_1684.Q ),
    .b(\DFF_1706.Q ),
    .y(_04425_)
  );
  al_nand2ft _10617_ (
    .a(\DFF_1706.Q ),
    .b(\DFF_1684.Q ),
    .y(_04426_)
  );
  al_ao21ttf _10618_ (
    .a(_04425_),
    .b(_04426_),
    .c(\DFF_1727.Q ),
    .y(_04427_)
  );
  al_nand3ftt _10619_ (
    .a(\DFF_1727.Q ),
    .b(_04425_),
    .c(_04426_),
    .y(_04428_)
  );
  al_aoi21 _10620_ (
    .a(_04428_),
    .b(_04427_),
    .c(_00451_),
    .y(\DFF_1707.D )
  );
  al_oa21ftt _10621_ (
    .a(\DFF_1683.Q ),
    .b(\DFF_1707.Q ),
    .c(RESET),
    .y(_04429_)
  );
  al_aoi21ftf _10622_ (
    .a(\DFF_1683.Q ),
    .b(\DFF_1707.Q ),
    .c(_04429_),
    .y(\DFF_1708.D )
  );
  al_oa21ftt _10623_ (
    .a(\DFF_1682.Q ),
    .b(\DFF_1708.Q ),
    .c(RESET),
    .y(_04430_)
  );
  al_aoi21ftf _10624_ (
    .a(\DFF_1682.Q ),
    .b(\DFF_1708.Q ),
    .c(_04430_),
    .y(\DFF_1709.D )
  );
  al_oa21ftt _10625_ (
    .a(\DFF_1681.Q ),
    .b(\DFF_1709.Q ),
    .c(RESET),
    .y(_04431_)
  );
  al_aoi21ftf _10626_ (
    .a(\DFF_1681.Q ),
    .b(\DFF_1709.Q ),
    .c(_04431_),
    .y(\DFF_1710.D )
  );
  al_oa21ftt _10627_ (
    .a(\DFF_1680.Q ),
    .b(\DFF_1710.Q ),
    .c(RESET),
    .y(_04432_)
  );
  al_aoi21ftf _10628_ (
    .a(\DFF_1680.Q ),
    .b(\DFF_1710.Q ),
    .c(_04432_),
    .y(\DFF_1711.D )
  );
  al_nand2ft _10629_ (
    .a(\DFF_1679.Q ),
    .b(\DFF_1711.Q ),
    .y(_04433_)
  );
  al_nand2ft _10630_ (
    .a(\DFF_1711.Q ),
    .b(\DFF_1679.Q ),
    .y(_04434_)
  );
  al_ao21ttf _10631_ (
    .a(_04433_),
    .b(_04434_),
    .c(\DFF_1727.Q ),
    .y(_04435_)
  );
  al_nand3ftt _10632_ (
    .a(\DFF_1727.Q ),
    .b(_04433_),
    .c(_04434_),
    .y(_04436_)
  );
  al_aoi21 _10633_ (
    .a(_04436_),
    .b(_04435_),
    .c(_00451_),
    .y(\DFF_1712.D )
  );
  al_oa21ftt _10634_ (
    .a(\DFF_1678.Q ),
    .b(\DFF_1712.Q ),
    .c(RESET),
    .y(_04437_)
  );
  al_aoi21ftf _10635_ (
    .a(\DFF_1678.Q ),
    .b(\DFF_1712.Q ),
    .c(_04437_),
    .y(\DFF_1713.D )
  );
  al_oa21ftt _10636_ (
    .a(\DFF_1677.Q ),
    .b(\DFF_1713.Q ),
    .c(RESET),
    .y(_04438_)
  );
  al_aoi21ftf _10637_ (
    .a(\DFF_1677.Q ),
    .b(\DFF_1713.Q ),
    .c(_04438_),
    .y(\DFF_1714.D )
  );
  al_oa21ftt _10638_ (
    .a(\DFF_1676.Q ),
    .b(\DFF_1714.Q ),
    .c(RESET),
    .y(_04439_)
  );
  al_aoi21ftf _10639_ (
    .a(\DFF_1676.Q ),
    .b(\DFF_1714.Q ),
    .c(_04439_),
    .y(\DFF_1715.D )
  );
  al_oa21ftt _10640_ (
    .a(\DFF_1675.Q ),
    .b(\DFF_1715.Q ),
    .c(RESET),
    .y(_04440_)
  );
  al_aoi21ftf _10641_ (
    .a(\DFF_1675.Q ),
    .b(\DFF_1715.Q ),
    .c(_04440_),
    .y(\DFF_1716.D )
  );
  al_oa21ftt _10642_ (
    .a(\DFF_1674.Q ),
    .b(\DFF_1716.Q ),
    .c(RESET),
    .y(_04441_)
  );
  al_aoi21ftf _10643_ (
    .a(\DFF_1674.Q ),
    .b(\DFF_1716.Q ),
    .c(_04441_),
    .y(\DFF_1717.D )
  );
  al_oa21ftt _10644_ (
    .a(\DFF_1673.Q ),
    .b(\DFF_1717.Q ),
    .c(RESET),
    .y(_04442_)
  );
  al_aoi21ftf _10645_ (
    .a(\DFF_1673.Q ),
    .b(\DFF_1717.Q ),
    .c(_04442_),
    .y(\DFF_1718.D )
  );
  al_oa21ftt _10646_ (
    .a(\DFF_1672.Q ),
    .b(\DFF_1718.Q ),
    .c(RESET),
    .y(_04443_)
  );
  al_aoi21ftf _10647_ (
    .a(\DFF_1672.Q ),
    .b(\DFF_1718.Q ),
    .c(_04443_),
    .y(\DFF_1719.D )
  );
  al_oa21ftt _10648_ (
    .a(\DFF_1671.Q ),
    .b(\DFF_1719.Q ),
    .c(RESET),
    .y(_04444_)
  );
  al_aoi21ftf _10649_ (
    .a(\DFF_1671.Q ),
    .b(\DFF_1719.Q ),
    .c(_04444_),
    .y(\DFF_1720.D )
  );
  al_oa21ftt _10650_ (
    .a(\DFF_1670.Q ),
    .b(\DFF_1720.Q ),
    .c(RESET),
    .y(_04445_)
  );
  al_aoi21ftf _10651_ (
    .a(\DFF_1670.Q ),
    .b(\DFF_1720.Q ),
    .c(_04445_),
    .y(\DFF_1721.D )
  );
  al_oa21ftt _10652_ (
    .a(\DFF_1669.Q ),
    .b(\DFF_1721.Q ),
    .c(RESET),
    .y(_04446_)
  );
  al_aoi21ftf _10653_ (
    .a(\DFF_1669.Q ),
    .b(\DFF_1721.Q ),
    .c(_04446_),
    .y(\DFF_1722.D )
  );
  al_oa21ftt _10654_ (
    .a(\DFF_1668.Q ),
    .b(\DFF_1722.Q ),
    .c(RESET),
    .y(_04447_)
  );
  al_aoi21ftf _10655_ (
    .a(\DFF_1668.Q ),
    .b(\DFF_1722.Q ),
    .c(_04447_),
    .y(\DFF_1723.D )
  );
  al_oa21ftt _10656_ (
    .a(\DFF_1667.Q ),
    .b(\DFF_1723.Q ),
    .c(RESET),
    .y(_04448_)
  );
  al_aoi21ftf _10657_ (
    .a(\DFF_1667.Q ),
    .b(\DFF_1723.Q ),
    .c(_04448_),
    .y(\DFF_1724.D )
  );
  al_oa21ftt _10658_ (
    .a(\DFF_1666.Q ),
    .b(\DFF_1724.Q ),
    .c(RESET),
    .y(_04449_)
  );
  al_aoi21ftf _10659_ (
    .a(\DFF_1666.Q ),
    .b(\DFF_1724.Q ),
    .c(_04449_),
    .y(\DFF_1725.D )
  );
  al_oa21ftt _10660_ (
    .a(\DFF_1665.Q ),
    .b(\DFF_1725.Q ),
    .c(RESET),
    .y(_04450_)
  );
  al_aoi21ftf _10661_ (
    .a(\DFF_1665.Q ),
    .b(\DFF_1725.Q ),
    .c(_04450_),
    .y(\DFF_1726.D )
  );
  al_oa21ftt _10662_ (
    .a(\DFF_1664.Q ),
    .b(\DFF_1726.Q ),
    .c(RESET),
    .y(_04451_)
  );
  al_aoi21ftf _10663_ (
    .a(\DFF_1664.Q ),
    .b(\DFF_1726.Q ),
    .c(_04451_),
    .y(\DFF_1727.D )
  );
  al_dffl _10664_ (
    .clk(CK),
    .d(\DFF_0.D ),
    .q(\DFF_0.Q )
  );
  al_dffl _10665_ (
    .clk(CK),
    .d(\DFF_1.D ),
    .q(\DFF_1.Q )
  );
  al_dffl _10666_ (
    .clk(CK),
    .d(\DFF_2.D ),
    .q(\DFF_2.Q )
  );
  al_dffl _10667_ (
    .clk(CK),
    .d(\DFF_3.D ),
    .q(\DFF_3.Q )
  );
  al_dffl _10668_ (
    .clk(CK),
    .d(\DFF_4.D ),
    .q(\DFF_4.Q )
  );
  al_dffl _10669_ (
    .clk(CK),
    .d(\DFF_5.D ),
    .q(\DFF_5.Q )
  );
  al_dffl _10670_ (
    .clk(CK),
    .d(\DFF_6.D ),
    .q(\DFF_6.Q )
  );
  al_dffl _10671_ (
    .clk(CK),
    .d(\DFF_7.D ),
    .q(\DFF_7.Q )
  );
  al_dffl _10672_ (
    .clk(CK),
    .d(\DFF_8.D ),
    .q(\DFF_8.Q )
  );
  al_dffl _10673_ (
    .clk(CK),
    .d(\DFF_9.D ),
    .q(\DFF_9.Q )
  );
  al_dffl _10674_ (
    .clk(CK),
    .d(\DFF_10.D ),
    .q(\DFF_10.Q )
  );
  al_dffl _10675_ (
    .clk(CK),
    .d(\DFF_11.D ),
    .q(\DFF_11.Q )
  );
  al_dffl _10676_ (
    .clk(CK),
    .d(\DFF_12.D ),
    .q(\DFF_12.Q )
  );
  al_dffl _10677_ (
    .clk(CK),
    .d(\DFF_13.D ),
    .q(\DFF_13.Q )
  );
  al_dffl _10678_ (
    .clk(CK),
    .d(\DFF_14.D ),
    .q(\DFF_14.Q )
  );
  al_dffl _10679_ (
    .clk(CK),
    .d(\DFF_15.D ),
    .q(\DFF_15.Q )
  );
  al_dffl _10680_ (
    .clk(CK),
    .d(\DFF_16.D ),
    .q(\DFF_16.Q )
  );
  al_dffl _10681_ (
    .clk(CK),
    .d(\DFF_17.D ),
    .q(\DFF_17.Q )
  );
  al_dffl _10682_ (
    .clk(CK),
    .d(\DFF_18.D ),
    .q(\DFF_18.Q )
  );
  al_dffl _10683_ (
    .clk(CK),
    .d(\DFF_19.D ),
    .q(\DFF_19.Q )
  );
  al_dffl _10684_ (
    .clk(CK),
    .d(\DFF_20.D ),
    .q(\DFF_20.Q )
  );
  al_dffl _10685_ (
    .clk(CK),
    .d(\DFF_21.D ),
    .q(\DFF_21.Q )
  );
  al_dffl _10686_ (
    .clk(CK),
    .d(\DFF_22.D ),
    .q(\DFF_22.Q )
  );
  al_dffl _10687_ (
    .clk(CK),
    .d(\DFF_23.D ),
    .q(\DFF_23.Q )
  );
  al_dffl _10688_ (
    .clk(CK),
    .d(\DFF_24.D ),
    .q(\DFF_24.Q )
  );
  al_dffl _10689_ (
    .clk(CK),
    .d(\DFF_25.D ),
    .q(\DFF_25.Q )
  );
  al_dffl _10690_ (
    .clk(CK),
    .d(\DFF_26.D ),
    .q(\DFF_26.Q )
  );
  al_dffl _10691_ (
    .clk(CK),
    .d(\DFF_27.D ),
    .q(\DFF_27.Q )
  );
  al_dffl _10692_ (
    .clk(CK),
    .d(\DFF_28.D ),
    .q(\DFF_28.Q )
  );
  al_dffl _10693_ (
    .clk(CK),
    .d(\DFF_29.D ),
    .q(\DFF_29.Q )
  );
  al_dffl _10694_ (
    .clk(CK),
    .d(\DFF_30.D ),
    .q(\DFF_30.Q )
  );
  al_dffl _10695_ (
    .clk(CK),
    .d(\DFF_31.D ),
    .q(\DFF_31.Q )
  );
  al_dffl _10696_ (
    .clk(CK),
    .d(\DFF_32.D ),
    .q(\DFF_32.Q )
  );
  al_dffl _10697_ (
    .clk(CK),
    .d(\DFF_33.D ),
    .q(\DFF_33.Q )
  );
  al_dffl _10698_ (
    .clk(CK),
    .d(\DFF_34.D ),
    .q(\DFF_34.Q )
  );
  al_dffl _10699_ (
    .clk(CK),
    .d(\DFF_35.D ),
    .q(\DFF_35.Q )
  );
  al_dffl _10700_ (
    .clk(CK),
    .d(\DFF_36.D ),
    .q(\DFF_36.Q )
  );
  al_dffl _10701_ (
    .clk(CK),
    .d(\DFF_37.D ),
    .q(\DFF_37.Q )
  );
  al_dffl _10702_ (
    .clk(CK),
    .d(\DFF_38.D ),
    .q(\DFF_38.Q )
  );
  al_dffl _10703_ (
    .clk(CK),
    .d(\DFF_39.D ),
    .q(\DFF_39.Q )
  );
  al_dffl _10704_ (
    .clk(CK),
    .d(\DFF_40.D ),
    .q(\DFF_40.Q )
  );
  al_dffl _10705_ (
    .clk(CK),
    .d(\DFF_41.D ),
    .q(\DFF_41.Q )
  );
  al_dffl _10706_ (
    .clk(CK),
    .d(\DFF_42.D ),
    .q(\DFF_42.Q )
  );
  al_dffl _10707_ (
    .clk(CK),
    .d(\DFF_43.D ),
    .q(\DFF_43.Q )
  );
  al_dffl _10708_ (
    .clk(CK),
    .d(\DFF_44.D ),
    .q(\DFF_44.Q )
  );
  al_dffl _10709_ (
    .clk(CK),
    .d(\DFF_45.D ),
    .q(\DFF_45.Q )
  );
  al_dffl _10710_ (
    .clk(CK),
    .d(\DFF_46.D ),
    .q(\DFF_46.Q )
  );
  al_dffl _10711_ (
    .clk(CK),
    .d(\DFF_47.D ),
    .q(\DFF_47.Q )
  );
  al_dffl _10712_ (
    .clk(CK),
    .d(\DFF_48.D ),
    .q(\DFF_48.Q )
  );
  al_dffl _10713_ (
    .clk(CK),
    .d(\DFF_49.D ),
    .q(\DFF_49.Q )
  );
  al_dffl _10714_ (
    .clk(CK),
    .d(\DFF_50.D ),
    .q(\DFF_50.Q )
  );
  al_dffl _10715_ (
    .clk(CK),
    .d(\DFF_51.D ),
    .q(\DFF_51.Q )
  );
  al_dffl _10716_ (
    .clk(CK),
    .d(\DFF_52.D ),
    .q(\DFF_52.Q )
  );
  al_dffl _10717_ (
    .clk(CK),
    .d(\DFF_53.D ),
    .q(\DFF_53.Q )
  );
  al_dffl _10718_ (
    .clk(CK),
    .d(\DFF_54.D ),
    .q(\DFF_54.Q )
  );
  al_dffl _10719_ (
    .clk(CK),
    .d(\DFF_55.D ),
    .q(\DFF_55.Q )
  );
  al_dffl _10720_ (
    .clk(CK),
    .d(\DFF_56.D ),
    .q(\DFF_56.Q )
  );
  al_dffl _10721_ (
    .clk(CK),
    .d(\DFF_57.D ),
    .q(\DFF_57.Q )
  );
  al_dffl _10722_ (
    .clk(CK),
    .d(\DFF_58.D ),
    .q(\DFF_58.Q )
  );
  al_dffl _10723_ (
    .clk(CK),
    .d(\DFF_59.D ),
    .q(\DFF_59.Q )
  );
  al_dffl _10724_ (
    .clk(CK),
    .d(\DFF_60.D ),
    .q(\DFF_60.Q )
  );
  al_dffl _10725_ (
    .clk(CK),
    .d(\DFF_61.D ),
    .q(\DFF_61.Q )
  );
  al_dffl _10726_ (
    .clk(CK),
    .d(\DFF_62.D ),
    .q(\DFF_62.Q )
  );
  al_dffl _10727_ (
    .clk(CK),
    .d(\DFF_63.D ),
    .q(\DFF_63.Q )
  );
  al_dffl _10728_ (
    .clk(CK),
    .d(\DFF_64.D ),
    .q(\DFF_64.Q )
  );
  al_dffl _10729_ (
    .clk(CK),
    .d(\DFF_65.D ),
    .q(\DFF_65.Q )
  );
  al_dffl _10730_ (
    .clk(CK),
    .d(\DFF_66.D ),
    .q(\DFF_66.Q )
  );
  al_dffl _10731_ (
    .clk(CK),
    .d(\DFF_67.D ),
    .q(\DFF_67.Q )
  );
  al_dffl _10732_ (
    .clk(CK),
    .d(\DFF_68.D ),
    .q(\DFF_68.Q )
  );
  al_dffl _10733_ (
    .clk(CK),
    .d(\DFF_69.D ),
    .q(\DFF_69.Q )
  );
  al_dffl _10734_ (
    .clk(CK),
    .d(\DFF_70.D ),
    .q(\DFF_70.Q )
  );
  al_dffl _10735_ (
    .clk(CK),
    .d(\DFF_71.D ),
    .q(\DFF_71.Q )
  );
  al_dffl _10736_ (
    .clk(CK),
    .d(\DFF_72.D ),
    .q(\DFF_72.Q )
  );
  al_dffl _10737_ (
    .clk(CK),
    .d(\DFF_73.D ),
    .q(\DFF_73.Q )
  );
  al_dffl _10738_ (
    .clk(CK),
    .d(\DFF_74.D ),
    .q(\DFF_74.Q )
  );
  al_dffl _10739_ (
    .clk(CK),
    .d(\DFF_75.D ),
    .q(\DFF_75.Q )
  );
  al_dffl _10740_ (
    .clk(CK),
    .d(\DFF_76.D ),
    .q(\DFF_76.Q )
  );
  al_dffl _10741_ (
    .clk(CK),
    .d(\DFF_77.D ),
    .q(\DFF_77.Q )
  );
  al_dffl _10742_ (
    .clk(CK),
    .d(\DFF_78.D ),
    .q(\DFF_78.Q )
  );
  al_dffl _10743_ (
    .clk(CK),
    .d(\DFF_79.D ),
    .q(\DFF_79.Q )
  );
  al_dffl _10744_ (
    .clk(CK),
    .d(\DFF_80.D ),
    .q(\DFF_80.Q )
  );
  al_dffl _10745_ (
    .clk(CK),
    .d(\DFF_81.D ),
    .q(\DFF_81.Q )
  );
  al_dffl _10746_ (
    .clk(CK),
    .d(\DFF_82.D ),
    .q(\DFF_82.Q )
  );
  al_dffl _10747_ (
    .clk(CK),
    .d(\DFF_83.D ),
    .q(\DFF_83.Q )
  );
  al_dffl _10748_ (
    .clk(CK),
    .d(\DFF_84.D ),
    .q(\DFF_84.Q )
  );
  al_dffl _10749_ (
    .clk(CK),
    .d(\DFF_85.D ),
    .q(\DFF_85.Q )
  );
  al_dffl _10750_ (
    .clk(CK),
    .d(\DFF_86.D ),
    .q(\DFF_86.Q )
  );
  al_dffl _10751_ (
    .clk(CK),
    .d(\DFF_87.D ),
    .q(\DFF_87.Q )
  );
  al_dffl _10752_ (
    .clk(CK),
    .d(\DFF_88.D ),
    .q(\DFF_88.Q )
  );
  al_dffl _10753_ (
    .clk(CK),
    .d(\DFF_89.D ),
    .q(\DFF_89.Q )
  );
  al_dffl _10754_ (
    .clk(CK),
    .d(\DFF_90.D ),
    .q(\DFF_90.Q )
  );
  al_dffl _10755_ (
    .clk(CK),
    .d(\DFF_91.D ),
    .q(\DFF_91.Q )
  );
  al_dffl _10756_ (
    .clk(CK),
    .d(\DFF_92.D ),
    .q(\DFF_92.Q )
  );
  al_dffl _10757_ (
    .clk(CK),
    .d(\DFF_93.D ),
    .q(\DFF_93.Q )
  );
  al_dffl _10758_ (
    .clk(CK),
    .d(\DFF_94.D ),
    .q(\DFF_94.Q )
  );
  al_dffl _10759_ (
    .clk(CK),
    .d(\DFF_95.D ),
    .q(\DFF_95.Q )
  );
  al_dffl _10760_ (
    .clk(CK),
    .d(\DFF_96.D ),
    .q(\DFF_96.Q )
  );
  al_dffl _10761_ (
    .clk(CK),
    .d(\DFF_97.D ),
    .q(\DFF_97.Q )
  );
  al_dffl _10762_ (
    .clk(CK),
    .d(\DFF_98.D ),
    .q(\DFF_98.Q )
  );
  al_dffl _10763_ (
    .clk(CK),
    .d(\DFF_99.D ),
    .q(\DFF_99.Q )
  );
  al_dffl _10764_ (
    .clk(CK),
    .d(\DFF_100.D ),
    .q(\DFF_100.Q )
  );
  al_dffl _10765_ (
    .clk(CK),
    .d(\DFF_101.D ),
    .q(\DFF_101.Q )
  );
  al_dffl _10766_ (
    .clk(CK),
    .d(\DFF_102.D ),
    .q(\DFF_102.Q )
  );
  al_dffl _10767_ (
    .clk(CK),
    .d(\DFF_103.D ),
    .q(\DFF_103.Q )
  );
  al_dffl _10768_ (
    .clk(CK),
    .d(\DFF_104.D ),
    .q(\DFF_104.Q )
  );
  al_dffl _10769_ (
    .clk(CK),
    .d(\DFF_105.D ),
    .q(\DFF_105.Q )
  );
  al_dffl _10770_ (
    .clk(CK),
    .d(\DFF_106.D ),
    .q(\DFF_106.Q )
  );
  al_dffl _10771_ (
    .clk(CK),
    .d(\DFF_107.D ),
    .q(\DFF_107.Q )
  );
  al_dffl _10772_ (
    .clk(CK),
    .d(\DFF_108.D ),
    .q(\DFF_108.Q )
  );
  al_dffl _10773_ (
    .clk(CK),
    .d(\DFF_109.D ),
    .q(\DFF_109.Q )
  );
  al_dffl _10774_ (
    .clk(CK),
    .d(\DFF_110.D ),
    .q(\DFF_110.Q )
  );
  al_dffl _10775_ (
    .clk(CK),
    .d(\DFF_111.D ),
    .q(\DFF_111.Q )
  );
  al_dffl _10776_ (
    .clk(CK),
    .d(\DFF_112.D ),
    .q(\DFF_112.Q )
  );
  al_dffl _10777_ (
    .clk(CK),
    .d(\DFF_113.D ),
    .q(\DFF_113.Q )
  );
  al_dffl _10778_ (
    .clk(CK),
    .d(\DFF_114.D ),
    .q(\DFF_114.Q )
  );
  al_dffl _10779_ (
    .clk(CK),
    .d(\DFF_115.D ),
    .q(\DFF_115.Q )
  );
  al_dffl _10780_ (
    .clk(CK),
    .d(\DFF_116.D ),
    .q(\DFF_116.Q )
  );
  al_dffl _10781_ (
    .clk(CK),
    .d(\DFF_117.D ),
    .q(\DFF_117.Q )
  );
  al_dffl _10782_ (
    .clk(CK),
    .d(\DFF_118.D ),
    .q(\DFF_118.Q )
  );
  al_dffl _10783_ (
    .clk(CK),
    .d(\DFF_119.D ),
    .q(\DFF_119.Q )
  );
  al_dffl _10784_ (
    .clk(CK),
    .d(\DFF_120.D ),
    .q(\DFF_120.Q )
  );
  al_dffl _10785_ (
    .clk(CK),
    .d(\DFF_121.D ),
    .q(\DFF_121.Q )
  );
  al_dffl _10786_ (
    .clk(CK),
    .d(\DFF_122.D ),
    .q(\DFF_122.Q )
  );
  al_dffl _10787_ (
    .clk(CK),
    .d(\DFF_123.D ),
    .q(\DFF_123.Q )
  );
  al_dffl _10788_ (
    .clk(CK),
    .d(\DFF_124.D ),
    .q(\DFF_124.Q )
  );
  al_dffl _10789_ (
    .clk(CK),
    .d(\DFF_125.D ),
    .q(\DFF_125.Q )
  );
  al_dffl _10790_ (
    .clk(CK),
    .d(\DFF_126.D ),
    .q(\DFF_126.Q )
  );
  al_dffl _10791_ (
    .clk(CK),
    .d(\DFF_127.D ),
    .q(\DFF_127.Q )
  );
  al_dffl _10792_ (
    .clk(CK),
    .d(\DFF_128.D ),
    .q(\DFF_128.Q )
  );
  al_dffl _10793_ (
    .clk(CK),
    .d(\DFF_129.D ),
    .q(\DFF_129.Q )
  );
  al_dffl _10794_ (
    .clk(CK),
    .d(\DFF_130.D ),
    .q(\DFF_130.Q )
  );
  al_dffl _10795_ (
    .clk(CK),
    .d(\DFF_131.D ),
    .q(\DFF_131.Q )
  );
  al_dffl _10796_ (
    .clk(CK),
    .d(\DFF_132.D ),
    .q(\DFF_132.Q )
  );
  al_dffl _10797_ (
    .clk(CK),
    .d(\DFF_133.D ),
    .q(\DFF_133.Q )
  );
  al_dffl _10798_ (
    .clk(CK),
    .d(\DFF_134.D ),
    .q(\DFF_134.Q )
  );
  al_dffl _10799_ (
    .clk(CK),
    .d(\DFF_135.D ),
    .q(\DFF_135.Q )
  );
  al_dffl _10800_ (
    .clk(CK),
    .d(\DFF_136.D ),
    .q(\DFF_136.Q )
  );
  al_dffl _10801_ (
    .clk(CK),
    .d(\DFF_137.D ),
    .q(\DFF_137.Q )
  );
  al_dffl _10802_ (
    .clk(CK),
    .d(\DFF_138.D ),
    .q(\DFF_138.Q )
  );
  al_dffl _10803_ (
    .clk(CK),
    .d(\DFF_139.D ),
    .q(\DFF_139.Q )
  );
  al_dffl _10804_ (
    .clk(CK),
    .d(\DFF_140.D ),
    .q(\DFF_140.Q )
  );
  al_dffl _10805_ (
    .clk(CK),
    .d(\DFF_141.D ),
    .q(\DFF_141.Q )
  );
  al_dffl _10806_ (
    .clk(CK),
    .d(\DFF_142.D ),
    .q(\DFF_142.Q )
  );
  al_dffl _10807_ (
    .clk(CK),
    .d(\DFF_143.D ),
    .q(\DFF_143.Q )
  );
  al_dffl _10808_ (
    .clk(CK),
    .d(\DFF_144.D ),
    .q(\DFF_144.Q )
  );
  al_dffl _10809_ (
    .clk(CK),
    .d(\DFF_145.D ),
    .q(\DFF_145.Q )
  );
  al_dffl _10810_ (
    .clk(CK),
    .d(\DFF_146.D ),
    .q(\DFF_146.Q )
  );
  al_dffl _10811_ (
    .clk(CK),
    .d(\DFF_147.D ),
    .q(\DFF_147.Q )
  );
  al_dffl _10812_ (
    .clk(CK),
    .d(\DFF_148.D ),
    .q(\DFF_148.Q )
  );
  al_dffl _10813_ (
    .clk(CK),
    .d(\DFF_149.D ),
    .q(\DFF_149.Q )
  );
  al_dffl _10814_ (
    .clk(CK),
    .d(\DFF_150.D ),
    .q(\DFF_150.Q )
  );
  al_dffl _10815_ (
    .clk(CK),
    .d(\DFF_151.D ),
    .q(\DFF_151.Q )
  );
  al_dffl _10816_ (
    .clk(CK),
    .d(\DFF_152.D ),
    .q(\DFF_152.Q )
  );
  al_dffl _10817_ (
    .clk(CK),
    .d(\DFF_153.D ),
    .q(\DFF_153.Q )
  );
  al_dffl _10818_ (
    .clk(CK),
    .d(\DFF_154.D ),
    .q(\DFF_154.Q )
  );
  al_dffl _10819_ (
    .clk(CK),
    .d(\DFF_155.D ),
    .q(\DFF_155.Q )
  );
  al_dffl _10820_ (
    .clk(CK),
    .d(\DFF_156.D ),
    .q(\DFF_156.Q )
  );
  al_dffl _10821_ (
    .clk(CK),
    .d(\DFF_157.D ),
    .q(\DFF_157.Q )
  );
  al_dffl _10822_ (
    .clk(CK),
    .d(\DFF_158.D ),
    .q(\DFF_158.Q )
  );
  al_dffl _10823_ (
    .clk(CK),
    .d(\DFF_159.D ),
    .q(\DFF_159.Q )
  );
  al_dffl _10824_ (
    .clk(CK),
    .d(\DFF_160.D ),
    .q(\DFF_160.Q )
  );
  al_dffl _10825_ (
    .clk(CK),
    .d(\DFF_161.D ),
    .q(\DFF_161.Q )
  );
  al_dffl _10826_ (
    .clk(CK),
    .d(\DFF_162.D ),
    .q(\DFF_162.Q )
  );
  al_dffl _10827_ (
    .clk(CK),
    .d(\DFF_163.D ),
    .q(\DFF_163.Q )
  );
  al_dffl _10828_ (
    .clk(CK),
    .d(\DFF_164.D ),
    .q(\DFF_164.Q )
  );
  al_dffl _10829_ (
    .clk(CK),
    .d(\DFF_165.D ),
    .q(\DFF_165.Q )
  );
  al_dffl _10830_ (
    .clk(CK),
    .d(\DFF_166.D ),
    .q(\DFF_166.Q )
  );
  al_dffl _10831_ (
    .clk(CK),
    .d(\DFF_167.D ),
    .q(\DFF_167.Q )
  );
  al_dffl _10832_ (
    .clk(CK),
    .d(\DFF_168.D ),
    .q(\DFF_168.Q )
  );
  al_dffl _10833_ (
    .clk(CK),
    .d(\DFF_169.D ),
    .q(\DFF_169.Q )
  );
  al_dffl _10834_ (
    .clk(CK),
    .d(\DFF_170.D ),
    .q(\DFF_170.Q )
  );
  al_dffl _10835_ (
    .clk(CK),
    .d(\DFF_171.D ),
    .q(\DFF_171.Q )
  );
  al_dffl _10836_ (
    .clk(CK),
    .d(\DFF_172.D ),
    .q(\DFF_172.Q )
  );
  al_dffl _10837_ (
    .clk(CK),
    .d(\DFF_173.D ),
    .q(\DFF_173.Q )
  );
  al_dffl _10838_ (
    .clk(CK),
    .d(\DFF_174.D ),
    .q(\DFF_174.Q )
  );
  al_dffl _10839_ (
    .clk(CK),
    .d(\DFF_175.D ),
    .q(\DFF_175.Q )
  );
  al_dffl _10840_ (
    .clk(CK),
    .d(\DFF_176.D ),
    .q(\DFF_176.Q )
  );
  al_dffl _10841_ (
    .clk(CK),
    .d(\DFF_177.D ),
    .q(\DFF_177.Q )
  );
  al_dffl _10842_ (
    .clk(CK),
    .d(\DFF_178.D ),
    .q(\DFF_178.Q )
  );
  al_dffl _10843_ (
    .clk(CK),
    .d(\DFF_179.D ),
    .q(\DFF_179.Q )
  );
  al_dffl _10844_ (
    .clk(CK),
    .d(\DFF_180.D ),
    .q(\DFF_180.Q )
  );
  al_dffl _10845_ (
    .clk(CK),
    .d(\DFF_181.D ),
    .q(\DFF_181.Q )
  );
  al_dffl _10846_ (
    .clk(CK),
    .d(\DFF_182.D ),
    .q(\DFF_182.Q )
  );
  al_dffl _10847_ (
    .clk(CK),
    .d(\DFF_183.D ),
    .q(\DFF_183.Q )
  );
  al_dffl _10848_ (
    .clk(CK),
    .d(\DFF_184.D ),
    .q(\DFF_184.Q )
  );
  al_dffl _10849_ (
    .clk(CK),
    .d(\DFF_185.D ),
    .q(\DFF_185.Q )
  );
  al_dffl _10850_ (
    .clk(CK),
    .d(\DFF_186.D ),
    .q(\DFF_186.Q )
  );
  al_dffl _10851_ (
    .clk(CK),
    .d(\DFF_187.D ),
    .q(\DFF_187.Q )
  );
  al_dffl _10852_ (
    .clk(CK),
    .d(\DFF_188.D ),
    .q(\DFF_188.Q )
  );
  al_dffl _10853_ (
    .clk(CK),
    .d(\DFF_189.D ),
    .q(\DFF_189.Q )
  );
  al_dffl _10854_ (
    .clk(CK),
    .d(\DFF_190.D ),
    .q(\DFF_190.Q )
  );
  al_dffl _10855_ (
    .clk(CK),
    .d(\DFF_191.D ),
    .q(\DFF_191.Q )
  );
  al_dffl _10856_ (
    .clk(CK),
    .d(\DFF_192.D ),
    .q(\DFF_192.Q )
  );
  al_dffl _10857_ (
    .clk(CK),
    .d(\DFF_193.D ),
    .q(\DFF_193.Q )
  );
  al_dffl _10858_ (
    .clk(CK),
    .d(\DFF_194.D ),
    .q(\DFF_194.Q )
  );
  al_dffl _10859_ (
    .clk(CK),
    .d(\DFF_195.D ),
    .q(\DFF_195.Q )
  );
  al_dffl _10860_ (
    .clk(CK),
    .d(\DFF_196.D ),
    .q(\DFF_196.Q )
  );
  al_dffl _10861_ (
    .clk(CK),
    .d(\DFF_197.D ),
    .q(\DFF_197.Q )
  );
  al_dffl _10862_ (
    .clk(CK),
    .d(\DFF_198.D ),
    .q(\DFF_198.Q )
  );
  al_dffl _10863_ (
    .clk(CK),
    .d(\DFF_199.D ),
    .q(\DFF_199.Q )
  );
  al_dffl _10864_ (
    .clk(CK),
    .d(\DFF_200.D ),
    .q(\DFF_200.Q )
  );
  al_dffl _10865_ (
    .clk(CK),
    .d(\DFF_201.D ),
    .q(\DFF_201.Q )
  );
  al_dffl _10866_ (
    .clk(CK),
    .d(\DFF_202.D ),
    .q(\DFF_202.Q )
  );
  al_dffl _10867_ (
    .clk(CK),
    .d(\DFF_203.D ),
    .q(\DFF_203.Q )
  );
  al_dffl _10868_ (
    .clk(CK),
    .d(\DFF_204.D ),
    .q(\DFF_204.Q )
  );
  al_dffl _10869_ (
    .clk(CK),
    .d(\DFF_205.D ),
    .q(\DFF_205.Q )
  );
  al_dffl _10870_ (
    .clk(CK),
    .d(\DFF_206.D ),
    .q(\DFF_206.Q )
  );
  al_dffl _10871_ (
    .clk(CK),
    .d(\DFF_207.D ),
    .q(\DFF_207.Q )
  );
  al_dffl _10872_ (
    .clk(CK),
    .d(\DFF_208.D ),
    .q(\DFF_208.Q )
  );
  al_dffl _10873_ (
    .clk(CK),
    .d(\DFF_209.D ),
    .q(\DFF_209.Q )
  );
  al_dffl _10874_ (
    .clk(CK),
    .d(\DFF_210.D ),
    .q(\DFF_210.Q )
  );
  al_dffl _10875_ (
    .clk(CK),
    .d(\DFF_211.D ),
    .q(\DFF_211.Q )
  );
  al_dffl _10876_ (
    .clk(CK),
    .d(\DFF_212.D ),
    .q(\DFF_212.Q )
  );
  al_dffl _10877_ (
    .clk(CK),
    .d(\DFF_213.D ),
    .q(\DFF_213.Q )
  );
  al_dffl _10878_ (
    .clk(CK),
    .d(\DFF_214.D ),
    .q(\DFF_214.Q )
  );
  al_dffl _10879_ (
    .clk(CK),
    .d(\DFF_215.D ),
    .q(\DFF_215.Q )
  );
  al_dffl _10880_ (
    .clk(CK),
    .d(\DFF_216.D ),
    .q(\DFF_216.Q )
  );
  al_dffl _10881_ (
    .clk(CK),
    .d(\DFF_217.D ),
    .q(\DFF_217.Q )
  );
  al_dffl _10882_ (
    .clk(CK),
    .d(\DFF_218.D ),
    .q(\DFF_218.Q )
  );
  al_dffl _10883_ (
    .clk(CK),
    .d(\DFF_219.D ),
    .q(\DFF_219.Q )
  );
  al_dffl _10884_ (
    .clk(CK),
    .d(\DFF_220.D ),
    .q(\DFF_220.Q )
  );
  al_dffl _10885_ (
    .clk(CK),
    .d(\DFF_221.D ),
    .q(\DFF_221.Q )
  );
  al_dffl _10886_ (
    .clk(CK),
    .d(\DFF_222.D ),
    .q(\DFF_222.Q )
  );
  al_dffl _10887_ (
    .clk(CK),
    .d(\DFF_223.D ),
    .q(\DFF_223.Q )
  );
  al_dffl _10888_ (
    .clk(CK),
    .d(\DFF_224.D ),
    .q(\DFF_224.Q )
  );
  al_dffl _10889_ (
    .clk(CK),
    .d(\DFF_225.D ),
    .q(\DFF_225.Q )
  );
  al_dffl _10890_ (
    .clk(CK),
    .d(\DFF_226.D ),
    .q(\DFF_226.Q )
  );
  al_dffl _10891_ (
    .clk(CK),
    .d(\DFF_227.D ),
    .q(\DFF_227.Q )
  );
  al_dffl _10892_ (
    .clk(CK),
    .d(\DFF_228.D ),
    .q(\DFF_228.Q )
  );
  al_dffl _10893_ (
    .clk(CK),
    .d(\DFF_229.D ),
    .q(\DFF_229.Q )
  );
  al_dffl _10894_ (
    .clk(CK),
    .d(\DFF_230.D ),
    .q(\DFF_230.Q )
  );
  al_dffl _10895_ (
    .clk(CK),
    .d(\DFF_231.D ),
    .q(\DFF_231.Q )
  );
  al_dffl _10896_ (
    .clk(CK),
    .d(\DFF_232.D ),
    .q(\DFF_232.Q )
  );
  al_dffl _10897_ (
    .clk(CK),
    .d(\DFF_233.D ),
    .q(\DFF_233.Q )
  );
  al_dffl _10898_ (
    .clk(CK),
    .d(\DFF_234.D ),
    .q(\DFF_234.Q )
  );
  al_dffl _10899_ (
    .clk(CK),
    .d(\DFF_235.D ),
    .q(\DFF_235.Q )
  );
  al_dffl _10900_ (
    .clk(CK),
    .d(\DFF_236.D ),
    .q(\DFF_236.Q )
  );
  al_dffl _10901_ (
    .clk(CK),
    .d(\DFF_237.D ),
    .q(\DFF_237.Q )
  );
  al_dffl _10902_ (
    .clk(CK),
    .d(\DFF_238.D ),
    .q(\DFF_238.Q )
  );
  al_dffl _10903_ (
    .clk(CK),
    .d(\DFF_239.D ),
    .q(\DFF_239.Q )
  );
  al_dffl _10904_ (
    .clk(CK),
    .d(\DFF_240.D ),
    .q(\DFF_240.Q )
  );
  al_dffl _10905_ (
    .clk(CK),
    .d(\DFF_241.D ),
    .q(\DFF_241.Q )
  );
  al_dffl _10906_ (
    .clk(CK),
    .d(\DFF_242.D ),
    .q(\DFF_242.Q )
  );
  al_dffl _10907_ (
    .clk(CK),
    .d(\DFF_243.D ),
    .q(\DFF_243.Q )
  );
  al_dffl _10908_ (
    .clk(CK),
    .d(\DFF_244.D ),
    .q(\DFF_244.Q )
  );
  al_dffl _10909_ (
    .clk(CK),
    .d(\DFF_245.D ),
    .q(\DFF_245.Q )
  );
  al_dffl _10910_ (
    .clk(CK),
    .d(\DFF_246.D ),
    .q(\DFF_246.Q )
  );
  al_dffl _10911_ (
    .clk(CK),
    .d(\DFF_247.D ),
    .q(\DFF_247.Q )
  );
  al_dffl _10912_ (
    .clk(CK),
    .d(\DFF_248.D ),
    .q(\DFF_248.Q )
  );
  al_dffl _10913_ (
    .clk(CK),
    .d(\DFF_249.D ),
    .q(\DFF_249.Q )
  );
  al_dffl _10914_ (
    .clk(CK),
    .d(\DFF_250.D ),
    .q(\DFF_250.Q )
  );
  al_dffl _10915_ (
    .clk(CK),
    .d(\DFF_251.D ),
    .q(\DFF_251.Q )
  );
  al_dffl _10916_ (
    .clk(CK),
    .d(\DFF_252.D ),
    .q(\DFF_252.Q )
  );
  al_dffl _10917_ (
    .clk(CK),
    .d(\DFF_253.D ),
    .q(\DFF_253.Q )
  );
  al_dffl _10918_ (
    .clk(CK),
    .d(\DFF_254.D ),
    .q(\DFF_254.Q )
  );
  al_dffl _10919_ (
    .clk(CK),
    .d(\DFF_255.D ),
    .q(\DFF_255.Q )
  );
  al_dffl _10920_ (
    .clk(CK),
    .d(\DFF_256.D ),
    .q(\DFF_256.Q )
  );
  al_dffl _10921_ (
    .clk(CK),
    .d(\DFF_257.D ),
    .q(\DFF_257.Q )
  );
  al_dffl _10922_ (
    .clk(CK),
    .d(\DFF_258.D ),
    .q(\DFF_258.Q )
  );
  al_dffl _10923_ (
    .clk(CK),
    .d(\DFF_259.D ),
    .q(\DFF_259.Q )
  );
  al_dffl _10924_ (
    .clk(CK),
    .d(\DFF_260.D ),
    .q(\DFF_260.Q )
  );
  al_dffl _10925_ (
    .clk(CK),
    .d(\DFF_261.D ),
    .q(\DFF_261.Q )
  );
  al_dffl _10926_ (
    .clk(CK),
    .d(\DFF_262.D ),
    .q(\DFF_262.Q )
  );
  al_dffl _10927_ (
    .clk(CK),
    .d(\DFF_263.D ),
    .q(\DFF_263.Q )
  );
  al_dffl _10928_ (
    .clk(CK),
    .d(\DFF_264.D ),
    .q(\DFF_264.Q )
  );
  al_dffl _10929_ (
    .clk(CK),
    .d(\DFF_265.D ),
    .q(\DFF_265.Q )
  );
  al_dffl _10930_ (
    .clk(CK),
    .d(\DFF_266.D ),
    .q(\DFF_266.Q )
  );
  al_dffl _10931_ (
    .clk(CK),
    .d(\DFF_267.D ),
    .q(\DFF_267.Q )
  );
  al_dffl _10932_ (
    .clk(CK),
    .d(\DFF_268.D ),
    .q(\DFF_268.Q )
  );
  al_dffl _10933_ (
    .clk(CK),
    .d(\DFF_269.D ),
    .q(\DFF_269.Q )
  );
  al_dffl _10934_ (
    .clk(CK),
    .d(\DFF_270.D ),
    .q(\DFF_270.Q )
  );
  al_dffl _10935_ (
    .clk(CK),
    .d(\DFF_271.D ),
    .q(\DFF_271.Q )
  );
  al_dffl _10936_ (
    .clk(CK),
    .d(\DFF_272.D ),
    .q(\DFF_272.Q )
  );
  al_dffl _10937_ (
    .clk(CK),
    .d(\DFF_273.D ),
    .q(\DFF_273.Q )
  );
  al_dffl _10938_ (
    .clk(CK),
    .d(\DFF_274.D ),
    .q(\DFF_274.Q )
  );
  al_dffl _10939_ (
    .clk(CK),
    .d(\DFF_275.D ),
    .q(\DFF_275.Q )
  );
  al_dffl _10940_ (
    .clk(CK),
    .d(\DFF_276.D ),
    .q(\DFF_276.Q )
  );
  al_dffl _10941_ (
    .clk(CK),
    .d(\DFF_277.D ),
    .q(\DFF_277.Q )
  );
  al_dffl _10942_ (
    .clk(CK),
    .d(\DFF_278.D ),
    .q(\DFF_278.Q )
  );
  al_dffl _10943_ (
    .clk(CK),
    .d(\DFF_279.D ),
    .q(\DFF_279.Q )
  );
  al_dffl _10944_ (
    .clk(CK),
    .d(\DFF_280.D ),
    .q(\DFF_280.Q )
  );
  al_dffl _10945_ (
    .clk(CK),
    .d(\DFF_281.D ),
    .q(\DFF_281.Q )
  );
  al_dffl _10946_ (
    .clk(CK),
    .d(\DFF_282.D ),
    .q(\DFF_282.Q )
  );
  al_dffl _10947_ (
    .clk(CK),
    .d(\DFF_283.D ),
    .q(\DFF_283.Q )
  );
  al_dffl _10948_ (
    .clk(CK),
    .d(\DFF_284.D ),
    .q(\DFF_284.Q )
  );
  al_dffl _10949_ (
    .clk(CK),
    .d(\DFF_285.D ),
    .q(\DFF_285.Q )
  );
  al_dffl _10950_ (
    .clk(CK),
    .d(\DFF_286.D ),
    .q(\DFF_286.Q )
  );
  al_dffl _10951_ (
    .clk(CK),
    .d(\DFF_287.D ),
    .q(\DFF_287.Q )
  );
  al_dffl _10952_ (
    .clk(CK),
    .d(\DFF_288.D ),
    .q(\DFF_288.Q )
  );
  al_dffl _10953_ (
    .clk(CK),
    .d(\DFF_289.D ),
    .q(\DFF_289.Q )
  );
  al_dffl _10954_ (
    .clk(CK),
    .d(\DFF_290.D ),
    .q(\DFF_290.Q )
  );
  al_dffl _10955_ (
    .clk(CK),
    .d(\DFF_291.D ),
    .q(\DFF_291.Q )
  );
  al_dffl _10956_ (
    .clk(CK),
    .d(\DFF_292.D ),
    .q(\DFF_292.Q )
  );
  al_dffl _10957_ (
    .clk(CK),
    .d(\DFF_293.D ),
    .q(\DFF_293.Q )
  );
  al_dffl _10958_ (
    .clk(CK),
    .d(\DFF_294.D ),
    .q(\DFF_294.Q )
  );
  al_dffl _10959_ (
    .clk(CK),
    .d(\DFF_295.D ),
    .q(\DFF_295.Q )
  );
  al_dffl _10960_ (
    .clk(CK),
    .d(\DFF_296.D ),
    .q(\DFF_296.Q )
  );
  al_dffl _10961_ (
    .clk(CK),
    .d(\DFF_297.D ),
    .q(\DFF_297.Q )
  );
  al_dffl _10962_ (
    .clk(CK),
    .d(\DFF_298.D ),
    .q(\DFF_298.Q )
  );
  al_dffl _10963_ (
    .clk(CK),
    .d(\DFF_299.D ),
    .q(\DFF_299.Q )
  );
  al_dffl _10964_ (
    .clk(CK),
    .d(\DFF_300.D ),
    .q(\DFF_300.Q )
  );
  al_dffl _10965_ (
    .clk(CK),
    .d(\DFF_301.D ),
    .q(\DFF_301.Q )
  );
  al_dffl _10966_ (
    .clk(CK),
    .d(\DFF_302.D ),
    .q(\DFF_302.Q )
  );
  al_dffl _10967_ (
    .clk(CK),
    .d(\DFF_303.D ),
    .q(\DFF_303.Q )
  );
  al_dffl _10968_ (
    .clk(CK),
    .d(\DFF_304.D ),
    .q(\DFF_304.Q )
  );
  al_dffl _10969_ (
    .clk(CK),
    .d(\DFF_305.D ),
    .q(\DFF_305.Q )
  );
  al_dffl _10970_ (
    .clk(CK),
    .d(\DFF_306.D ),
    .q(\DFF_306.Q )
  );
  al_dffl _10971_ (
    .clk(CK),
    .d(\DFF_307.D ),
    .q(\DFF_307.Q )
  );
  al_dffl _10972_ (
    .clk(CK),
    .d(\DFF_308.D ),
    .q(\DFF_308.Q )
  );
  al_dffl _10973_ (
    .clk(CK),
    .d(\DFF_309.D ),
    .q(\DFF_309.Q )
  );
  al_dffl _10974_ (
    .clk(CK),
    .d(\DFF_310.D ),
    .q(\DFF_310.Q )
  );
  al_dffl _10975_ (
    .clk(CK),
    .d(\DFF_311.D ),
    .q(\DFF_311.Q )
  );
  al_dffl _10976_ (
    .clk(CK),
    .d(\DFF_312.D ),
    .q(\DFF_312.Q )
  );
  al_dffl _10977_ (
    .clk(CK),
    .d(\DFF_313.D ),
    .q(\DFF_313.Q )
  );
  al_dffl _10978_ (
    .clk(CK),
    .d(\DFF_314.D ),
    .q(\DFF_314.Q )
  );
  al_dffl _10979_ (
    .clk(CK),
    .d(\DFF_315.D ),
    .q(\DFF_315.Q )
  );
  al_dffl _10980_ (
    .clk(CK),
    .d(\DFF_316.D ),
    .q(\DFF_316.Q )
  );
  al_dffl _10981_ (
    .clk(CK),
    .d(\DFF_317.D ),
    .q(\DFF_317.Q )
  );
  al_dffl _10982_ (
    .clk(CK),
    .d(\DFF_318.D ),
    .q(\DFF_318.Q )
  );
  al_dffl _10983_ (
    .clk(CK),
    .d(\DFF_319.D ),
    .q(\DFF_319.Q )
  );
  al_dffl _10984_ (
    .clk(CK),
    .d(\DFF_320.D ),
    .q(\DFF_320.Q )
  );
  al_dffl _10985_ (
    .clk(CK),
    .d(\DFF_321.D ),
    .q(\DFF_321.Q )
  );
  al_dffl _10986_ (
    .clk(CK),
    .d(\DFF_322.D ),
    .q(\DFF_322.Q )
  );
  al_dffl _10987_ (
    .clk(CK),
    .d(\DFF_323.D ),
    .q(\DFF_323.Q )
  );
  al_dffl _10988_ (
    .clk(CK),
    .d(\DFF_324.D ),
    .q(\DFF_324.Q )
  );
  al_dffl _10989_ (
    .clk(CK),
    .d(\DFF_325.D ),
    .q(\DFF_325.Q )
  );
  al_dffl _10990_ (
    .clk(CK),
    .d(\DFF_326.D ),
    .q(\DFF_326.Q )
  );
  al_dffl _10991_ (
    .clk(CK),
    .d(\DFF_327.D ),
    .q(\DFF_327.Q )
  );
  al_dffl _10992_ (
    .clk(CK),
    .d(\DFF_328.D ),
    .q(\DFF_328.Q )
  );
  al_dffl _10993_ (
    .clk(CK),
    .d(\DFF_329.D ),
    .q(\DFF_329.Q )
  );
  al_dffl _10994_ (
    .clk(CK),
    .d(\DFF_330.D ),
    .q(\DFF_330.Q )
  );
  al_dffl _10995_ (
    .clk(CK),
    .d(\DFF_331.D ),
    .q(\DFF_331.Q )
  );
  al_dffl _10996_ (
    .clk(CK),
    .d(\DFF_332.D ),
    .q(\DFF_332.Q )
  );
  al_dffl _10997_ (
    .clk(CK),
    .d(\DFF_333.D ),
    .q(\DFF_333.Q )
  );
  al_dffl _10998_ (
    .clk(CK),
    .d(\DFF_334.D ),
    .q(\DFF_334.Q )
  );
  al_dffl _10999_ (
    .clk(CK),
    .d(\DFF_335.D ),
    .q(\DFF_335.Q )
  );
  al_dffl _11000_ (
    .clk(CK),
    .d(\DFF_336.D ),
    .q(\DFF_336.Q )
  );
  al_dffl _11001_ (
    .clk(CK),
    .d(\DFF_337.D ),
    .q(\DFF_337.Q )
  );
  al_dffl _11002_ (
    .clk(CK),
    .d(\DFF_338.D ),
    .q(\DFF_338.Q )
  );
  al_dffl _11003_ (
    .clk(CK),
    .d(\DFF_339.D ),
    .q(\DFF_339.Q )
  );
  al_dffl _11004_ (
    .clk(CK),
    .d(\DFF_340.D ),
    .q(\DFF_340.Q )
  );
  al_dffl _11005_ (
    .clk(CK),
    .d(\DFF_341.D ),
    .q(\DFF_341.Q )
  );
  al_dffl _11006_ (
    .clk(CK),
    .d(\DFF_342.D ),
    .q(\DFF_342.Q )
  );
  al_dffl _11007_ (
    .clk(CK),
    .d(\DFF_343.D ),
    .q(\DFF_343.Q )
  );
  al_dffl _11008_ (
    .clk(CK),
    .d(\DFF_344.D ),
    .q(\DFF_344.Q )
  );
  al_dffl _11009_ (
    .clk(CK),
    .d(\DFF_345.D ),
    .q(\DFF_345.Q )
  );
  al_dffl _11010_ (
    .clk(CK),
    .d(\DFF_346.D ),
    .q(\DFF_346.Q )
  );
  al_dffl _11011_ (
    .clk(CK),
    .d(\DFF_347.D ),
    .q(\DFF_347.Q )
  );
  al_dffl _11012_ (
    .clk(CK),
    .d(\DFF_348.D ),
    .q(\DFF_348.Q )
  );
  al_dffl _11013_ (
    .clk(CK),
    .d(\DFF_349.D ),
    .q(\DFF_349.Q )
  );
  al_dffl _11014_ (
    .clk(CK),
    .d(\DFF_350.D ),
    .q(\DFF_350.Q )
  );
  al_dffl _11015_ (
    .clk(CK),
    .d(\DFF_351.D ),
    .q(\DFF_351.Q )
  );
  al_dffl _11016_ (
    .clk(CK),
    .d(\DFF_352.D ),
    .q(\DFF_352.Q )
  );
  al_dffl _11017_ (
    .clk(CK),
    .d(\DFF_353.D ),
    .q(\DFF_353.Q )
  );
  al_dffl _11018_ (
    .clk(CK),
    .d(\DFF_354.D ),
    .q(\DFF_354.Q )
  );
  al_dffl _11019_ (
    .clk(CK),
    .d(\DFF_355.D ),
    .q(\DFF_355.Q )
  );
  al_dffl _11020_ (
    .clk(CK),
    .d(\DFF_356.D ),
    .q(\DFF_356.Q )
  );
  al_dffl _11021_ (
    .clk(CK),
    .d(\DFF_357.D ),
    .q(\DFF_357.Q )
  );
  al_dffl _11022_ (
    .clk(CK),
    .d(\DFF_358.D ),
    .q(\DFF_358.Q )
  );
  al_dffl _11023_ (
    .clk(CK),
    .d(\DFF_359.D ),
    .q(\DFF_359.Q )
  );
  al_dffl _11024_ (
    .clk(CK),
    .d(\DFF_360.D ),
    .q(\DFF_360.Q )
  );
  al_dffl _11025_ (
    .clk(CK),
    .d(\DFF_361.D ),
    .q(\DFF_361.Q )
  );
  al_dffl _11026_ (
    .clk(CK),
    .d(\DFF_362.D ),
    .q(\DFF_362.Q )
  );
  al_dffl _11027_ (
    .clk(CK),
    .d(\DFF_363.D ),
    .q(\DFF_363.Q )
  );
  al_dffl _11028_ (
    .clk(CK),
    .d(\DFF_364.D ),
    .q(\DFF_364.Q )
  );
  al_dffl _11029_ (
    .clk(CK),
    .d(\DFF_365.D ),
    .q(\DFF_365.Q )
  );
  al_dffl _11030_ (
    .clk(CK),
    .d(\DFF_366.D ),
    .q(\DFF_366.Q )
  );
  al_dffl _11031_ (
    .clk(CK),
    .d(\DFF_367.D ),
    .q(\DFF_367.Q )
  );
  al_dffl _11032_ (
    .clk(CK),
    .d(\DFF_368.D ),
    .q(\DFF_368.Q )
  );
  al_dffl _11033_ (
    .clk(CK),
    .d(\DFF_369.D ),
    .q(\DFF_369.Q )
  );
  al_dffl _11034_ (
    .clk(CK),
    .d(\DFF_370.D ),
    .q(\DFF_370.Q )
  );
  al_dffl _11035_ (
    .clk(CK),
    .d(\DFF_371.D ),
    .q(\DFF_371.Q )
  );
  al_dffl _11036_ (
    .clk(CK),
    .d(\DFF_372.D ),
    .q(\DFF_372.Q )
  );
  al_dffl _11037_ (
    .clk(CK),
    .d(\DFF_373.D ),
    .q(\DFF_373.Q )
  );
  al_dffl _11038_ (
    .clk(CK),
    .d(\DFF_374.D ),
    .q(\DFF_374.Q )
  );
  al_dffl _11039_ (
    .clk(CK),
    .d(\DFF_375.D ),
    .q(\DFF_375.Q )
  );
  al_dffl _11040_ (
    .clk(CK),
    .d(\DFF_376.D ),
    .q(\DFF_376.Q )
  );
  al_dffl _11041_ (
    .clk(CK),
    .d(\DFF_377.D ),
    .q(\DFF_377.Q )
  );
  al_dffl _11042_ (
    .clk(CK),
    .d(\DFF_378.D ),
    .q(\DFF_378.Q )
  );
  al_dffl _11043_ (
    .clk(CK),
    .d(\DFF_379.D ),
    .q(\DFF_379.Q )
  );
  al_dffl _11044_ (
    .clk(CK),
    .d(\DFF_380.D ),
    .q(\DFF_380.Q )
  );
  al_dffl _11045_ (
    .clk(CK),
    .d(\DFF_381.D ),
    .q(\DFF_381.Q )
  );
  al_dffl _11046_ (
    .clk(CK),
    .d(\DFF_382.D ),
    .q(\DFF_382.Q )
  );
  al_dffl _11047_ (
    .clk(CK),
    .d(\DFF_383.D ),
    .q(\DFF_383.Q )
  );
  al_dffl _11048_ (
    .clk(CK),
    .d(\DFF_384.D ),
    .q(\DFF_384.Q )
  );
  al_dffl _11049_ (
    .clk(CK),
    .d(\DFF_385.D ),
    .q(\DFF_385.Q )
  );
  al_dffl _11050_ (
    .clk(CK),
    .d(\DFF_386.D ),
    .q(\DFF_386.Q )
  );
  al_dffl _11051_ (
    .clk(CK),
    .d(\DFF_387.D ),
    .q(\DFF_387.Q )
  );
  al_dffl _11052_ (
    .clk(CK),
    .d(\DFF_388.D ),
    .q(\DFF_388.Q )
  );
  al_dffl _11053_ (
    .clk(CK),
    .d(\DFF_389.D ),
    .q(\DFF_389.Q )
  );
  al_dffl _11054_ (
    .clk(CK),
    .d(\DFF_390.D ),
    .q(\DFF_390.Q )
  );
  al_dffl _11055_ (
    .clk(CK),
    .d(\DFF_391.D ),
    .q(\DFF_391.Q )
  );
  al_dffl _11056_ (
    .clk(CK),
    .d(\DFF_392.D ),
    .q(\DFF_392.Q )
  );
  al_dffl _11057_ (
    .clk(CK),
    .d(\DFF_393.D ),
    .q(\DFF_393.Q )
  );
  al_dffl _11058_ (
    .clk(CK),
    .d(\DFF_394.D ),
    .q(\DFF_394.Q )
  );
  al_dffl _11059_ (
    .clk(CK),
    .d(\DFF_395.D ),
    .q(\DFF_395.Q )
  );
  al_dffl _11060_ (
    .clk(CK),
    .d(\DFF_396.D ),
    .q(\DFF_396.Q )
  );
  al_dffl _11061_ (
    .clk(CK),
    .d(\DFF_397.D ),
    .q(\DFF_397.Q )
  );
  al_dffl _11062_ (
    .clk(CK),
    .d(\DFF_398.D ),
    .q(\DFF_398.Q )
  );
  al_dffl _11063_ (
    .clk(CK),
    .d(\DFF_399.D ),
    .q(\DFF_399.Q )
  );
  al_dffl _11064_ (
    .clk(CK),
    .d(\DFF_400.D ),
    .q(\DFF_400.Q )
  );
  al_dffl _11065_ (
    .clk(CK),
    .d(\DFF_401.D ),
    .q(\DFF_401.Q )
  );
  al_dffl _11066_ (
    .clk(CK),
    .d(\DFF_402.D ),
    .q(\DFF_402.Q )
  );
  al_dffl _11067_ (
    .clk(CK),
    .d(\DFF_403.D ),
    .q(\DFF_403.Q )
  );
  al_dffl _11068_ (
    .clk(CK),
    .d(\DFF_404.D ),
    .q(\DFF_404.Q )
  );
  al_dffl _11069_ (
    .clk(CK),
    .d(\DFF_405.D ),
    .q(\DFF_405.Q )
  );
  al_dffl _11070_ (
    .clk(CK),
    .d(\DFF_406.D ),
    .q(\DFF_406.Q )
  );
  al_dffl _11071_ (
    .clk(CK),
    .d(\DFF_407.D ),
    .q(\DFF_407.Q )
  );
  al_dffl _11072_ (
    .clk(CK),
    .d(\DFF_408.D ),
    .q(\DFF_408.Q )
  );
  al_dffl _11073_ (
    .clk(CK),
    .d(\DFF_409.D ),
    .q(\DFF_409.Q )
  );
  al_dffl _11074_ (
    .clk(CK),
    .d(\DFF_410.D ),
    .q(\DFF_410.Q )
  );
  al_dffl _11075_ (
    .clk(CK),
    .d(\DFF_411.D ),
    .q(\DFF_411.Q )
  );
  al_dffl _11076_ (
    .clk(CK),
    .d(\DFF_412.D ),
    .q(\DFF_412.Q )
  );
  al_dffl _11077_ (
    .clk(CK),
    .d(\DFF_413.D ),
    .q(\DFF_413.Q )
  );
  al_dffl _11078_ (
    .clk(CK),
    .d(\DFF_414.D ),
    .q(\DFF_414.Q )
  );
  al_dffl _11079_ (
    .clk(CK),
    .d(\DFF_415.D ),
    .q(\DFF_415.Q )
  );
  al_dffl _11080_ (
    .clk(CK),
    .d(\DFF_416.D ),
    .q(\DFF_416.Q )
  );
  al_dffl _11081_ (
    .clk(CK),
    .d(\DFF_417.D ),
    .q(\DFF_417.Q )
  );
  al_dffl _11082_ (
    .clk(CK),
    .d(\DFF_418.D ),
    .q(\DFF_418.Q )
  );
  al_dffl _11083_ (
    .clk(CK),
    .d(\DFF_419.D ),
    .q(\DFF_419.Q )
  );
  al_dffl _11084_ (
    .clk(CK),
    .d(\DFF_420.D ),
    .q(\DFF_420.Q )
  );
  al_dffl _11085_ (
    .clk(CK),
    .d(\DFF_421.D ),
    .q(\DFF_421.Q )
  );
  al_dffl _11086_ (
    .clk(CK),
    .d(\DFF_422.D ),
    .q(\DFF_422.Q )
  );
  al_dffl _11087_ (
    .clk(CK),
    .d(\DFF_423.D ),
    .q(\DFF_423.Q )
  );
  al_dffl _11088_ (
    .clk(CK),
    .d(\DFF_424.D ),
    .q(\DFF_424.Q )
  );
  al_dffl _11089_ (
    .clk(CK),
    .d(\DFF_425.D ),
    .q(\DFF_425.Q )
  );
  al_dffl _11090_ (
    .clk(CK),
    .d(\DFF_426.D ),
    .q(\DFF_426.Q )
  );
  al_dffl _11091_ (
    .clk(CK),
    .d(\DFF_427.D ),
    .q(\DFF_427.Q )
  );
  al_dffl _11092_ (
    .clk(CK),
    .d(\DFF_428.D ),
    .q(\DFF_428.Q )
  );
  al_dffl _11093_ (
    .clk(CK),
    .d(\DFF_429.D ),
    .q(\DFF_429.Q )
  );
  al_dffl _11094_ (
    .clk(CK),
    .d(\DFF_430.D ),
    .q(\DFF_430.Q )
  );
  al_dffl _11095_ (
    .clk(CK),
    .d(\DFF_431.D ),
    .q(\DFF_431.Q )
  );
  al_dffl _11096_ (
    .clk(CK),
    .d(\DFF_432.D ),
    .q(\DFF_432.Q )
  );
  al_dffl _11097_ (
    .clk(CK),
    .d(\DFF_433.D ),
    .q(\DFF_433.Q )
  );
  al_dffl _11098_ (
    .clk(CK),
    .d(\DFF_434.D ),
    .q(\DFF_434.Q )
  );
  al_dffl _11099_ (
    .clk(CK),
    .d(\DFF_435.D ),
    .q(\DFF_435.Q )
  );
  al_dffl _11100_ (
    .clk(CK),
    .d(\DFF_436.D ),
    .q(\DFF_436.Q )
  );
  al_dffl _11101_ (
    .clk(CK),
    .d(\DFF_437.D ),
    .q(\DFF_437.Q )
  );
  al_dffl _11102_ (
    .clk(CK),
    .d(\DFF_438.D ),
    .q(\DFF_438.Q )
  );
  al_dffl _11103_ (
    .clk(CK),
    .d(\DFF_439.D ),
    .q(\DFF_439.Q )
  );
  al_dffl _11104_ (
    .clk(CK),
    .d(\DFF_440.D ),
    .q(\DFF_440.Q )
  );
  al_dffl _11105_ (
    .clk(CK),
    .d(\DFF_441.D ),
    .q(\DFF_441.Q )
  );
  al_dffl _11106_ (
    .clk(CK),
    .d(\DFF_442.D ),
    .q(\DFF_442.Q )
  );
  al_dffl _11107_ (
    .clk(CK),
    .d(\DFF_443.D ),
    .q(\DFF_443.Q )
  );
  al_dffl _11108_ (
    .clk(CK),
    .d(\DFF_444.D ),
    .q(\DFF_444.Q )
  );
  al_dffl _11109_ (
    .clk(CK),
    .d(\DFF_445.D ),
    .q(\DFF_445.Q )
  );
  al_dffl _11110_ (
    .clk(CK),
    .d(\DFF_446.D ),
    .q(\DFF_446.Q )
  );
  al_dffl _11111_ (
    .clk(CK),
    .d(\DFF_447.D ),
    .q(\DFF_447.Q )
  );
  al_dffl _11112_ (
    .clk(CK),
    .d(\DFF_448.D ),
    .q(\DFF_448.Q )
  );
  al_dffl _11113_ (
    .clk(CK),
    .d(\DFF_449.D ),
    .q(\DFF_449.Q )
  );
  al_dffl _11114_ (
    .clk(CK),
    .d(\DFF_450.D ),
    .q(\DFF_450.Q )
  );
  al_dffl _11115_ (
    .clk(CK),
    .d(\DFF_451.D ),
    .q(\DFF_451.Q )
  );
  al_dffl _11116_ (
    .clk(CK),
    .d(\DFF_452.D ),
    .q(\DFF_452.Q )
  );
  al_dffl _11117_ (
    .clk(CK),
    .d(\DFF_453.D ),
    .q(\DFF_453.Q )
  );
  al_dffl _11118_ (
    .clk(CK),
    .d(\DFF_454.D ),
    .q(\DFF_454.Q )
  );
  al_dffl _11119_ (
    .clk(CK),
    .d(\DFF_455.D ),
    .q(\DFF_455.Q )
  );
  al_dffl _11120_ (
    .clk(CK),
    .d(\DFF_456.D ),
    .q(\DFF_456.Q )
  );
  al_dffl _11121_ (
    .clk(CK),
    .d(\DFF_457.D ),
    .q(\DFF_457.Q )
  );
  al_dffl _11122_ (
    .clk(CK),
    .d(\DFF_458.D ),
    .q(\DFF_458.Q )
  );
  al_dffl _11123_ (
    .clk(CK),
    .d(\DFF_459.D ),
    .q(\DFF_459.Q )
  );
  al_dffl _11124_ (
    .clk(CK),
    .d(\DFF_460.D ),
    .q(\DFF_460.Q )
  );
  al_dffl _11125_ (
    .clk(CK),
    .d(\DFF_461.D ),
    .q(\DFF_461.Q )
  );
  al_dffl _11126_ (
    .clk(CK),
    .d(\DFF_462.D ),
    .q(\DFF_462.Q )
  );
  al_dffl _11127_ (
    .clk(CK),
    .d(\DFF_463.D ),
    .q(\DFF_463.Q )
  );
  al_dffl _11128_ (
    .clk(CK),
    .d(\DFF_464.D ),
    .q(\DFF_464.Q )
  );
  al_dffl _11129_ (
    .clk(CK),
    .d(\DFF_465.D ),
    .q(\DFF_465.Q )
  );
  al_dffl _11130_ (
    .clk(CK),
    .d(\DFF_466.D ),
    .q(\DFF_466.Q )
  );
  al_dffl _11131_ (
    .clk(CK),
    .d(\DFF_467.D ),
    .q(\DFF_467.Q )
  );
  al_dffl _11132_ (
    .clk(CK),
    .d(\DFF_468.D ),
    .q(\DFF_468.Q )
  );
  al_dffl _11133_ (
    .clk(CK),
    .d(\DFF_469.D ),
    .q(\DFF_469.Q )
  );
  al_dffl _11134_ (
    .clk(CK),
    .d(\DFF_470.D ),
    .q(\DFF_470.Q )
  );
  al_dffl _11135_ (
    .clk(CK),
    .d(\DFF_471.D ),
    .q(\DFF_471.Q )
  );
  al_dffl _11136_ (
    .clk(CK),
    .d(\DFF_472.D ),
    .q(\DFF_472.Q )
  );
  al_dffl _11137_ (
    .clk(CK),
    .d(\DFF_473.D ),
    .q(\DFF_473.Q )
  );
  al_dffl _11138_ (
    .clk(CK),
    .d(\DFF_474.D ),
    .q(\DFF_474.Q )
  );
  al_dffl _11139_ (
    .clk(CK),
    .d(\DFF_475.D ),
    .q(\DFF_475.Q )
  );
  al_dffl _11140_ (
    .clk(CK),
    .d(\DFF_476.D ),
    .q(\DFF_476.Q )
  );
  al_dffl _11141_ (
    .clk(CK),
    .d(\DFF_477.D ),
    .q(\DFF_477.Q )
  );
  al_dffl _11142_ (
    .clk(CK),
    .d(\DFF_478.D ),
    .q(\DFF_478.Q )
  );
  al_dffl _11143_ (
    .clk(CK),
    .d(\DFF_479.D ),
    .q(\DFF_479.Q )
  );
  al_dffl _11144_ (
    .clk(CK),
    .d(\DFF_480.D ),
    .q(\DFF_480.Q )
  );
  al_dffl _11145_ (
    .clk(CK),
    .d(\DFF_481.D ),
    .q(\DFF_481.Q )
  );
  al_dffl _11146_ (
    .clk(CK),
    .d(\DFF_482.D ),
    .q(\DFF_482.Q )
  );
  al_dffl _11147_ (
    .clk(CK),
    .d(\DFF_483.D ),
    .q(\DFF_483.Q )
  );
  al_dffl _11148_ (
    .clk(CK),
    .d(\DFF_484.D ),
    .q(\DFF_484.Q )
  );
  al_dffl _11149_ (
    .clk(CK),
    .d(\DFF_485.D ),
    .q(\DFF_485.Q )
  );
  al_dffl _11150_ (
    .clk(CK),
    .d(\DFF_486.D ),
    .q(\DFF_486.Q )
  );
  al_dffl _11151_ (
    .clk(CK),
    .d(\DFF_487.D ),
    .q(\DFF_487.Q )
  );
  al_dffl _11152_ (
    .clk(CK),
    .d(\DFF_488.D ),
    .q(\DFF_488.Q )
  );
  al_dffl _11153_ (
    .clk(CK),
    .d(\DFF_489.D ),
    .q(\DFF_489.Q )
  );
  al_dffl _11154_ (
    .clk(CK),
    .d(\DFF_490.D ),
    .q(\DFF_490.Q )
  );
  al_dffl _11155_ (
    .clk(CK),
    .d(\DFF_491.D ),
    .q(\DFF_491.Q )
  );
  al_dffl _11156_ (
    .clk(CK),
    .d(\DFF_492.D ),
    .q(\DFF_492.Q )
  );
  al_dffl _11157_ (
    .clk(CK),
    .d(\DFF_493.D ),
    .q(\DFF_493.Q )
  );
  al_dffl _11158_ (
    .clk(CK),
    .d(\DFF_494.D ),
    .q(\DFF_494.Q )
  );
  al_dffl _11159_ (
    .clk(CK),
    .d(\DFF_495.D ),
    .q(\DFF_495.Q )
  );
  al_dffl _11160_ (
    .clk(CK),
    .d(\DFF_496.D ),
    .q(\DFF_496.Q )
  );
  al_dffl _11161_ (
    .clk(CK),
    .d(\DFF_497.D ),
    .q(\DFF_497.Q )
  );
  al_dffl _11162_ (
    .clk(CK),
    .d(\DFF_498.D ),
    .q(\DFF_498.Q )
  );
  al_dffl _11163_ (
    .clk(CK),
    .d(\DFF_499.D ),
    .q(\DFF_499.Q )
  );
  al_dffl _11164_ (
    .clk(CK),
    .d(\DFF_500.D ),
    .q(\DFF_500.Q )
  );
  al_dffl _11165_ (
    .clk(CK),
    .d(\DFF_501.D ),
    .q(\DFF_501.Q )
  );
  al_dffl _11166_ (
    .clk(CK),
    .d(\DFF_502.D ),
    .q(\DFF_502.Q )
  );
  al_dffl _11167_ (
    .clk(CK),
    .d(\DFF_503.D ),
    .q(\DFF_503.Q )
  );
  al_dffl _11168_ (
    .clk(CK),
    .d(\DFF_504.D ),
    .q(\DFF_504.Q )
  );
  al_dffl _11169_ (
    .clk(CK),
    .d(\DFF_505.D ),
    .q(\DFF_505.Q )
  );
  al_dffl _11170_ (
    .clk(CK),
    .d(\DFF_506.D ),
    .q(\DFF_506.Q )
  );
  al_dffl _11171_ (
    .clk(CK),
    .d(\DFF_507.D ),
    .q(\DFF_507.Q )
  );
  al_dffl _11172_ (
    .clk(CK),
    .d(\DFF_508.D ),
    .q(\DFF_508.Q )
  );
  al_dffl _11173_ (
    .clk(CK),
    .d(\DFF_509.D ),
    .q(\DFF_509.Q )
  );
  al_dffl _11174_ (
    .clk(CK),
    .d(\DFF_510.D ),
    .q(\DFF_510.Q )
  );
  al_dffl _11175_ (
    .clk(CK),
    .d(\DFF_511.D ),
    .q(\DFF_511.Q )
  );
  al_dffl _11176_ (
    .clk(CK),
    .d(\DFF_512.D ),
    .q(\DFF_512.Q )
  );
  al_dffl _11177_ (
    .clk(CK),
    .d(\DFF_513.D ),
    .q(\DFF_513.Q )
  );
  al_dffl _11178_ (
    .clk(CK),
    .d(\DFF_514.D ),
    .q(\DFF_514.Q )
  );
  al_dffl _11179_ (
    .clk(CK),
    .d(\DFF_515.D ),
    .q(\DFF_515.Q )
  );
  al_dffl _11180_ (
    .clk(CK),
    .d(\DFF_516.D ),
    .q(\DFF_516.Q )
  );
  al_dffl _11181_ (
    .clk(CK),
    .d(\DFF_517.D ),
    .q(\DFF_517.Q )
  );
  al_dffl _11182_ (
    .clk(CK),
    .d(\DFF_518.D ),
    .q(\DFF_518.Q )
  );
  al_dffl _11183_ (
    .clk(CK),
    .d(\DFF_519.D ),
    .q(\DFF_519.Q )
  );
  al_dffl _11184_ (
    .clk(CK),
    .d(\DFF_520.D ),
    .q(\DFF_520.Q )
  );
  al_dffl _11185_ (
    .clk(CK),
    .d(\DFF_521.D ),
    .q(\DFF_521.Q )
  );
  al_dffl _11186_ (
    .clk(CK),
    .d(\DFF_522.D ),
    .q(\DFF_522.Q )
  );
  al_dffl _11187_ (
    .clk(CK),
    .d(\DFF_523.D ),
    .q(\DFF_523.Q )
  );
  al_dffl _11188_ (
    .clk(CK),
    .d(\DFF_524.D ),
    .q(\DFF_524.Q )
  );
  al_dffl _11189_ (
    .clk(CK),
    .d(\DFF_525.D ),
    .q(\DFF_525.Q )
  );
  al_dffl _11190_ (
    .clk(CK),
    .d(\DFF_526.D ),
    .q(\DFF_526.Q )
  );
  al_dffl _11191_ (
    .clk(CK),
    .d(\DFF_527.D ),
    .q(\DFF_527.Q )
  );
  al_dffl _11192_ (
    .clk(CK),
    .d(\DFF_528.D ),
    .q(\DFF_528.Q )
  );
  al_dffl _11193_ (
    .clk(CK),
    .d(\DFF_529.D ),
    .q(\DFF_529.Q )
  );
  al_dffl _11194_ (
    .clk(CK),
    .d(\DFF_530.D ),
    .q(\DFF_530.Q )
  );
  al_dffl _11195_ (
    .clk(CK),
    .d(\DFF_531.D ),
    .q(\DFF_531.Q )
  );
  al_dffl _11196_ (
    .clk(CK),
    .d(\DFF_532.D ),
    .q(\DFF_532.Q )
  );
  al_dffl _11197_ (
    .clk(CK),
    .d(\DFF_533.D ),
    .q(\DFF_533.Q )
  );
  al_dffl _11198_ (
    .clk(CK),
    .d(\DFF_534.D ),
    .q(\DFF_534.Q )
  );
  al_dffl _11199_ (
    .clk(CK),
    .d(\DFF_535.D ),
    .q(\DFF_535.Q )
  );
  al_dffl _11200_ (
    .clk(CK),
    .d(\DFF_536.D ),
    .q(\DFF_536.Q )
  );
  al_dffl _11201_ (
    .clk(CK),
    .d(\DFF_537.D ),
    .q(\DFF_537.Q )
  );
  al_dffl _11202_ (
    .clk(CK),
    .d(\DFF_538.D ),
    .q(\DFF_538.Q )
  );
  al_dffl _11203_ (
    .clk(CK),
    .d(\DFF_539.D ),
    .q(\DFF_539.Q )
  );
  al_dffl _11204_ (
    .clk(CK),
    .d(\DFF_540.D ),
    .q(\DFF_540.Q )
  );
  al_dffl _11205_ (
    .clk(CK),
    .d(\DFF_541.D ),
    .q(\DFF_541.Q )
  );
  al_dffl _11206_ (
    .clk(CK),
    .d(\DFF_542.D ),
    .q(\DFF_542.Q )
  );
  al_dffl _11207_ (
    .clk(CK),
    .d(\DFF_543.D ),
    .q(\DFF_543.Q )
  );
  al_dffl _11208_ (
    .clk(CK),
    .d(\DFF_544.D ),
    .q(\DFF_544.Q )
  );
  al_dffl _11209_ (
    .clk(CK),
    .d(\DFF_545.D ),
    .q(\DFF_545.Q )
  );
  al_dffl _11210_ (
    .clk(CK),
    .d(\DFF_546.D ),
    .q(\DFF_546.Q )
  );
  al_dffl _11211_ (
    .clk(CK),
    .d(\DFF_547.D ),
    .q(\DFF_547.Q )
  );
  al_dffl _11212_ (
    .clk(CK),
    .d(\DFF_548.D ),
    .q(\DFF_548.Q )
  );
  al_dffl _11213_ (
    .clk(CK),
    .d(\DFF_549.D ),
    .q(\DFF_549.Q )
  );
  al_dffl _11214_ (
    .clk(CK),
    .d(\DFF_550.D ),
    .q(\DFF_550.Q )
  );
  al_dffl _11215_ (
    .clk(CK),
    .d(\DFF_551.D ),
    .q(\DFF_551.Q )
  );
  al_dffl _11216_ (
    .clk(CK),
    .d(\DFF_552.D ),
    .q(\DFF_552.Q )
  );
  al_dffl _11217_ (
    .clk(CK),
    .d(\DFF_553.D ),
    .q(\DFF_553.Q )
  );
  al_dffl _11218_ (
    .clk(CK),
    .d(\DFF_554.D ),
    .q(\DFF_554.Q )
  );
  al_dffl _11219_ (
    .clk(CK),
    .d(\DFF_555.D ),
    .q(\DFF_555.Q )
  );
  al_dffl _11220_ (
    .clk(CK),
    .d(\DFF_556.D ),
    .q(\DFF_556.Q )
  );
  al_dffl _11221_ (
    .clk(CK),
    .d(\DFF_557.D ),
    .q(\DFF_557.Q )
  );
  al_dffl _11222_ (
    .clk(CK),
    .d(\DFF_558.D ),
    .q(\DFF_558.Q )
  );
  al_dffl _11223_ (
    .clk(CK),
    .d(\DFF_559.D ),
    .q(\DFF_559.Q )
  );
  al_dffl _11224_ (
    .clk(CK),
    .d(\DFF_560.D ),
    .q(\DFF_560.Q )
  );
  al_dffl _11225_ (
    .clk(CK),
    .d(\DFF_561.D ),
    .q(\DFF_561.Q )
  );
  al_dffl _11226_ (
    .clk(CK),
    .d(\DFF_562.D ),
    .q(\DFF_562.Q )
  );
  al_dffl _11227_ (
    .clk(CK),
    .d(\DFF_563.D ),
    .q(\DFF_563.Q )
  );
  al_dffl _11228_ (
    .clk(CK),
    .d(\DFF_564.D ),
    .q(\DFF_564.Q )
  );
  al_dffl _11229_ (
    .clk(CK),
    .d(\DFF_565.D ),
    .q(\DFF_565.Q )
  );
  al_dffl _11230_ (
    .clk(CK),
    .d(\DFF_566.D ),
    .q(\DFF_566.Q )
  );
  al_dffl _11231_ (
    .clk(CK),
    .d(\DFF_567.D ),
    .q(\DFF_567.Q )
  );
  al_dffl _11232_ (
    .clk(CK),
    .d(\DFF_568.D ),
    .q(\DFF_568.Q )
  );
  al_dffl _11233_ (
    .clk(CK),
    .d(\DFF_569.D ),
    .q(\DFF_569.Q )
  );
  al_dffl _11234_ (
    .clk(CK),
    .d(\DFF_570.D ),
    .q(\DFF_570.Q )
  );
  al_dffl _11235_ (
    .clk(CK),
    .d(\DFF_571.D ),
    .q(\DFF_571.Q )
  );
  al_dffl _11236_ (
    .clk(CK),
    .d(\DFF_572.D ),
    .q(\DFF_572.Q )
  );
  al_dffl _11237_ (
    .clk(CK),
    .d(\DFF_573.D ),
    .q(\DFF_573.Q )
  );
  al_dffl _11238_ (
    .clk(CK),
    .d(\DFF_574.D ),
    .q(\DFF_574.Q )
  );
  al_dffl _11239_ (
    .clk(CK),
    .d(\DFF_575.D ),
    .q(\DFF_575.Q )
  );
  al_dffl _11240_ (
    .clk(CK),
    .d(\DFF_576.D ),
    .q(\DFF_576.Q )
  );
  al_dffl _11241_ (
    .clk(CK),
    .d(\DFF_577.D ),
    .q(\DFF_577.Q )
  );
  al_dffl _11242_ (
    .clk(CK),
    .d(\DFF_578.D ),
    .q(\DFF_578.Q )
  );
  al_dffl _11243_ (
    .clk(CK),
    .d(\DFF_579.D ),
    .q(\DFF_579.Q )
  );
  al_dffl _11244_ (
    .clk(CK),
    .d(\DFF_580.D ),
    .q(\DFF_580.Q )
  );
  al_dffl _11245_ (
    .clk(CK),
    .d(\DFF_581.D ),
    .q(\DFF_581.Q )
  );
  al_dffl _11246_ (
    .clk(CK),
    .d(\DFF_582.D ),
    .q(\DFF_582.Q )
  );
  al_dffl _11247_ (
    .clk(CK),
    .d(\DFF_583.D ),
    .q(\DFF_583.Q )
  );
  al_dffl _11248_ (
    .clk(CK),
    .d(\DFF_584.D ),
    .q(\DFF_584.Q )
  );
  al_dffl _11249_ (
    .clk(CK),
    .d(\DFF_585.D ),
    .q(\DFF_585.Q )
  );
  al_dffl _11250_ (
    .clk(CK),
    .d(\DFF_586.D ),
    .q(\DFF_586.Q )
  );
  al_dffl _11251_ (
    .clk(CK),
    .d(\DFF_587.D ),
    .q(\DFF_587.Q )
  );
  al_dffl _11252_ (
    .clk(CK),
    .d(\DFF_588.D ),
    .q(\DFF_588.Q )
  );
  al_dffl _11253_ (
    .clk(CK),
    .d(\DFF_589.D ),
    .q(\DFF_589.Q )
  );
  al_dffl _11254_ (
    .clk(CK),
    .d(\DFF_590.D ),
    .q(\DFF_590.Q )
  );
  al_dffl _11255_ (
    .clk(CK),
    .d(\DFF_591.D ),
    .q(\DFF_591.Q )
  );
  al_dffl _11256_ (
    .clk(CK),
    .d(\DFF_592.D ),
    .q(\DFF_592.Q )
  );
  al_dffl _11257_ (
    .clk(CK),
    .d(\DFF_593.D ),
    .q(\DFF_593.Q )
  );
  al_dffl _11258_ (
    .clk(CK),
    .d(\DFF_594.D ),
    .q(\DFF_594.Q )
  );
  al_dffl _11259_ (
    .clk(CK),
    .d(\DFF_595.D ),
    .q(\DFF_595.Q )
  );
  al_dffl _11260_ (
    .clk(CK),
    .d(\DFF_596.D ),
    .q(\DFF_596.Q )
  );
  al_dffl _11261_ (
    .clk(CK),
    .d(\DFF_597.D ),
    .q(\DFF_597.Q )
  );
  al_dffl _11262_ (
    .clk(CK),
    .d(\DFF_598.D ),
    .q(\DFF_598.Q )
  );
  al_dffl _11263_ (
    .clk(CK),
    .d(\DFF_599.D ),
    .q(\DFF_599.Q )
  );
  al_dffl _11264_ (
    .clk(CK),
    .d(\DFF_600.D ),
    .q(\DFF_600.Q )
  );
  al_dffl _11265_ (
    .clk(CK),
    .d(\DFF_601.D ),
    .q(\DFF_601.Q )
  );
  al_dffl _11266_ (
    .clk(CK),
    .d(\DFF_602.D ),
    .q(\DFF_602.Q )
  );
  al_dffl _11267_ (
    .clk(CK),
    .d(\DFF_603.D ),
    .q(\DFF_603.Q )
  );
  al_dffl _11268_ (
    .clk(CK),
    .d(\DFF_604.D ),
    .q(\DFF_604.Q )
  );
  al_dffl _11269_ (
    .clk(CK),
    .d(\DFF_605.D ),
    .q(\DFF_605.Q )
  );
  al_dffl _11270_ (
    .clk(CK),
    .d(\DFF_606.D ),
    .q(\DFF_606.Q )
  );
  al_dffl _11271_ (
    .clk(CK),
    .d(\DFF_607.D ),
    .q(\DFF_607.Q )
  );
  al_dffl _11272_ (
    .clk(CK),
    .d(\DFF_608.D ),
    .q(\DFF_608.Q )
  );
  al_dffl _11273_ (
    .clk(CK),
    .d(\DFF_609.D ),
    .q(\DFF_609.Q )
  );
  al_dffl _11274_ (
    .clk(CK),
    .d(\DFF_610.D ),
    .q(\DFF_610.Q )
  );
  al_dffl _11275_ (
    .clk(CK),
    .d(\DFF_611.D ),
    .q(\DFF_611.Q )
  );
  al_dffl _11276_ (
    .clk(CK),
    .d(\DFF_612.D ),
    .q(\DFF_612.Q )
  );
  al_dffl _11277_ (
    .clk(CK),
    .d(\DFF_613.D ),
    .q(\DFF_613.Q )
  );
  al_dffl _11278_ (
    .clk(CK),
    .d(\DFF_614.D ),
    .q(\DFF_614.Q )
  );
  al_dffl _11279_ (
    .clk(CK),
    .d(\DFF_615.D ),
    .q(\DFF_615.Q )
  );
  al_dffl _11280_ (
    .clk(CK),
    .d(\DFF_616.D ),
    .q(\DFF_616.Q )
  );
  al_dffl _11281_ (
    .clk(CK),
    .d(\DFF_617.D ),
    .q(\DFF_617.Q )
  );
  al_dffl _11282_ (
    .clk(CK),
    .d(\DFF_618.D ),
    .q(\DFF_618.Q )
  );
  al_dffl _11283_ (
    .clk(CK),
    .d(\DFF_619.D ),
    .q(\DFF_619.Q )
  );
  al_dffl _11284_ (
    .clk(CK),
    .d(\DFF_620.D ),
    .q(\DFF_620.Q )
  );
  al_dffl _11285_ (
    .clk(CK),
    .d(\DFF_621.D ),
    .q(\DFF_621.Q )
  );
  al_dffl _11286_ (
    .clk(CK),
    .d(\DFF_622.D ),
    .q(\DFF_622.Q )
  );
  al_dffl _11287_ (
    .clk(CK),
    .d(\DFF_623.D ),
    .q(\DFF_623.Q )
  );
  al_dffl _11288_ (
    .clk(CK),
    .d(\DFF_624.D ),
    .q(\DFF_624.Q )
  );
  al_dffl _11289_ (
    .clk(CK),
    .d(\DFF_625.D ),
    .q(\DFF_625.Q )
  );
  al_dffl _11290_ (
    .clk(CK),
    .d(\DFF_626.D ),
    .q(\DFF_626.Q )
  );
  al_dffl _11291_ (
    .clk(CK),
    .d(\DFF_627.D ),
    .q(\DFF_627.Q )
  );
  al_dffl _11292_ (
    .clk(CK),
    .d(\DFF_628.D ),
    .q(\DFF_628.Q )
  );
  al_dffl _11293_ (
    .clk(CK),
    .d(\DFF_629.D ),
    .q(\DFF_629.Q )
  );
  al_dffl _11294_ (
    .clk(CK),
    .d(\DFF_630.D ),
    .q(\DFF_630.Q )
  );
  al_dffl _11295_ (
    .clk(CK),
    .d(\DFF_631.D ),
    .q(\DFF_631.Q )
  );
  al_dffl _11296_ (
    .clk(CK),
    .d(\DFF_632.D ),
    .q(\DFF_632.Q )
  );
  al_dffl _11297_ (
    .clk(CK),
    .d(\DFF_633.D ),
    .q(\DFF_633.Q )
  );
  al_dffl _11298_ (
    .clk(CK),
    .d(\DFF_634.D ),
    .q(\DFF_634.Q )
  );
  al_dffl _11299_ (
    .clk(CK),
    .d(\DFF_635.D ),
    .q(\DFF_635.Q )
  );
  al_dffl _11300_ (
    .clk(CK),
    .d(\DFF_636.D ),
    .q(\DFF_636.Q )
  );
  al_dffl _11301_ (
    .clk(CK),
    .d(\DFF_637.D ),
    .q(\DFF_637.Q )
  );
  al_dffl _11302_ (
    .clk(CK),
    .d(\DFF_638.D ),
    .q(\DFF_638.Q )
  );
  al_dffl _11303_ (
    .clk(CK),
    .d(\DFF_639.D ),
    .q(\DFF_639.Q )
  );
  al_dffl _11304_ (
    .clk(CK),
    .d(\DFF_640.D ),
    .q(\DFF_640.Q )
  );
  al_dffl _11305_ (
    .clk(CK),
    .d(\DFF_641.D ),
    .q(\DFF_641.Q )
  );
  al_dffl _11306_ (
    .clk(CK),
    .d(\DFF_642.D ),
    .q(\DFF_642.Q )
  );
  al_dffl _11307_ (
    .clk(CK),
    .d(\DFF_643.D ),
    .q(\DFF_643.Q )
  );
  al_dffl _11308_ (
    .clk(CK),
    .d(\DFF_644.D ),
    .q(\DFF_644.Q )
  );
  al_dffl _11309_ (
    .clk(CK),
    .d(\DFF_645.D ),
    .q(\DFF_645.Q )
  );
  al_dffl _11310_ (
    .clk(CK),
    .d(\DFF_646.D ),
    .q(\DFF_646.Q )
  );
  al_dffl _11311_ (
    .clk(CK),
    .d(\DFF_647.D ),
    .q(\DFF_647.Q )
  );
  al_dffl _11312_ (
    .clk(CK),
    .d(\DFF_648.D ),
    .q(\DFF_648.Q )
  );
  al_dffl _11313_ (
    .clk(CK),
    .d(\DFF_649.D ),
    .q(\DFF_649.Q )
  );
  al_dffl _11314_ (
    .clk(CK),
    .d(\DFF_650.D ),
    .q(\DFF_650.Q )
  );
  al_dffl _11315_ (
    .clk(CK),
    .d(\DFF_651.D ),
    .q(\DFF_651.Q )
  );
  al_dffl _11316_ (
    .clk(CK),
    .d(\DFF_652.D ),
    .q(\DFF_652.Q )
  );
  al_dffl _11317_ (
    .clk(CK),
    .d(\DFF_653.D ),
    .q(\DFF_653.Q )
  );
  al_dffl _11318_ (
    .clk(CK),
    .d(\DFF_654.D ),
    .q(\DFF_654.Q )
  );
  al_dffl _11319_ (
    .clk(CK),
    .d(\DFF_655.D ),
    .q(\DFF_655.Q )
  );
  al_dffl _11320_ (
    .clk(CK),
    .d(\DFF_656.D ),
    .q(\DFF_656.Q )
  );
  al_dffl _11321_ (
    .clk(CK),
    .d(\DFF_657.D ),
    .q(\DFF_657.Q )
  );
  al_dffl _11322_ (
    .clk(CK),
    .d(\DFF_658.D ),
    .q(\DFF_658.Q )
  );
  al_dffl _11323_ (
    .clk(CK),
    .d(\DFF_659.D ),
    .q(\DFF_659.Q )
  );
  al_dffl _11324_ (
    .clk(CK),
    .d(\DFF_660.D ),
    .q(\DFF_660.Q )
  );
  al_dffl _11325_ (
    .clk(CK),
    .d(\DFF_661.D ),
    .q(\DFF_661.Q )
  );
  al_dffl _11326_ (
    .clk(CK),
    .d(\DFF_662.D ),
    .q(\DFF_662.Q )
  );
  al_dffl _11327_ (
    .clk(CK),
    .d(\DFF_663.D ),
    .q(\DFF_663.Q )
  );
  al_dffl _11328_ (
    .clk(CK),
    .d(\DFF_664.D ),
    .q(\DFF_664.Q )
  );
  al_dffl _11329_ (
    .clk(CK),
    .d(\DFF_665.D ),
    .q(\DFF_665.Q )
  );
  al_dffl _11330_ (
    .clk(CK),
    .d(\DFF_666.D ),
    .q(\DFF_666.Q )
  );
  al_dffl _11331_ (
    .clk(CK),
    .d(\DFF_667.D ),
    .q(\DFF_667.Q )
  );
  al_dffl _11332_ (
    .clk(CK),
    .d(\DFF_668.D ),
    .q(\DFF_668.Q )
  );
  al_dffl _11333_ (
    .clk(CK),
    .d(\DFF_669.D ),
    .q(\DFF_669.Q )
  );
  al_dffl _11334_ (
    .clk(CK),
    .d(\DFF_670.D ),
    .q(\DFF_670.Q )
  );
  al_dffl _11335_ (
    .clk(CK),
    .d(\DFF_671.D ),
    .q(\DFF_671.Q )
  );
  al_dffl _11336_ (
    .clk(CK),
    .d(\DFF_672.D ),
    .q(\DFF_672.Q )
  );
  al_dffl _11337_ (
    .clk(CK),
    .d(\DFF_673.D ),
    .q(\DFF_673.Q )
  );
  al_dffl _11338_ (
    .clk(CK),
    .d(\DFF_674.D ),
    .q(\DFF_674.Q )
  );
  al_dffl _11339_ (
    .clk(CK),
    .d(\DFF_675.D ),
    .q(\DFF_675.Q )
  );
  al_dffl _11340_ (
    .clk(CK),
    .d(\DFF_676.D ),
    .q(\DFF_676.Q )
  );
  al_dffl _11341_ (
    .clk(CK),
    .d(\DFF_677.D ),
    .q(\DFF_677.Q )
  );
  al_dffl _11342_ (
    .clk(CK),
    .d(\DFF_678.D ),
    .q(\DFF_678.Q )
  );
  al_dffl _11343_ (
    .clk(CK),
    .d(\DFF_679.D ),
    .q(\DFF_679.Q )
  );
  al_dffl _11344_ (
    .clk(CK),
    .d(\DFF_680.D ),
    .q(\DFF_680.Q )
  );
  al_dffl _11345_ (
    .clk(CK),
    .d(\DFF_681.D ),
    .q(\DFF_681.Q )
  );
  al_dffl _11346_ (
    .clk(CK),
    .d(\DFF_682.D ),
    .q(\DFF_682.Q )
  );
  al_dffl _11347_ (
    .clk(CK),
    .d(\DFF_683.D ),
    .q(\DFF_683.Q )
  );
  al_dffl _11348_ (
    .clk(CK),
    .d(\DFF_684.D ),
    .q(\DFF_684.Q )
  );
  al_dffl _11349_ (
    .clk(CK),
    .d(\DFF_685.D ),
    .q(\DFF_685.Q )
  );
  al_dffl _11350_ (
    .clk(CK),
    .d(\DFF_686.D ),
    .q(\DFF_686.Q )
  );
  al_dffl _11351_ (
    .clk(CK),
    .d(\DFF_687.D ),
    .q(\DFF_687.Q )
  );
  al_dffl _11352_ (
    .clk(CK),
    .d(\DFF_688.D ),
    .q(\DFF_688.Q )
  );
  al_dffl _11353_ (
    .clk(CK),
    .d(\DFF_689.D ),
    .q(\DFF_689.Q )
  );
  al_dffl _11354_ (
    .clk(CK),
    .d(\DFF_690.D ),
    .q(\DFF_690.Q )
  );
  al_dffl _11355_ (
    .clk(CK),
    .d(\DFF_691.D ),
    .q(\DFF_691.Q )
  );
  al_dffl _11356_ (
    .clk(CK),
    .d(\DFF_692.D ),
    .q(\DFF_692.Q )
  );
  al_dffl _11357_ (
    .clk(CK),
    .d(\DFF_693.D ),
    .q(\DFF_693.Q )
  );
  al_dffl _11358_ (
    .clk(CK),
    .d(\DFF_694.D ),
    .q(\DFF_694.Q )
  );
  al_dffl _11359_ (
    .clk(CK),
    .d(\DFF_695.D ),
    .q(\DFF_695.Q )
  );
  al_dffl _11360_ (
    .clk(CK),
    .d(\DFF_696.D ),
    .q(\DFF_696.Q )
  );
  al_dffl _11361_ (
    .clk(CK),
    .d(\DFF_697.D ),
    .q(\DFF_697.Q )
  );
  al_dffl _11362_ (
    .clk(CK),
    .d(\DFF_698.D ),
    .q(\DFF_698.Q )
  );
  al_dffl _11363_ (
    .clk(CK),
    .d(\DFF_699.D ),
    .q(\DFF_699.Q )
  );
  al_dffl _11364_ (
    .clk(CK),
    .d(\DFF_700.D ),
    .q(\DFF_700.Q )
  );
  al_dffl _11365_ (
    .clk(CK),
    .d(\DFF_701.D ),
    .q(\DFF_701.Q )
  );
  al_dffl _11366_ (
    .clk(CK),
    .d(\DFF_702.D ),
    .q(\DFF_702.Q )
  );
  al_dffl _11367_ (
    .clk(CK),
    .d(\DFF_703.D ),
    .q(\DFF_703.Q )
  );
  al_dffl _11368_ (
    .clk(CK),
    .d(\DFF_704.D ),
    .q(\DFF_704.Q )
  );
  al_dffl _11369_ (
    .clk(CK),
    .d(\DFF_705.D ),
    .q(\DFF_705.Q )
  );
  al_dffl _11370_ (
    .clk(CK),
    .d(\DFF_706.D ),
    .q(\DFF_706.Q )
  );
  al_dffl _11371_ (
    .clk(CK),
    .d(\DFF_707.D ),
    .q(\DFF_707.Q )
  );
  al_dffl _11372_ (
    .clk(CK),
    .d(\DFF_708.D ),
    .q(\DFF_708.Q )
  );
  al_dffl _11373_ (
    .clk(CK),
    .d(\DFF_709.D ),
    .q(\DFF_709.Q )
  );
  al_dffl _11374_ (
    .clk(CK),
    .d(\DFF_710.D ),
    .q(\DFF_710.Q )
  );
  al_dffl _11375_ (
    .clk(CK),
    .d(\DFF_711.D ),
    .q(\DFF_711.Q )
  );
  al_dffl _11376_ (
    .clk(CK),
    .d(\DFF_712.D ),
    .q(\DFF_712.Q )
  );
  al_dffl _11377_ (
    .clk(CK),
    .d(\DFF_713.D ),
    .q(\DFF_713.Q )
  );
  al_dffl _11378_ (
    .clk(CK),
    .d(\DFF_714.D ),
    .q(\DFF_714.Q )
  );
  al_dffl _11379_ (
    .clk(CK),
    .d(\DFF_715.D ),
    .q(\DFF_715.Q )
  );
  al_dffl _11380_ (
    .clk(CK),
    .d(\DFF_716.D ),
    .q(\DFF_716.Q )
  );
  al_dffl _11381_ (
    .clk(CK),
    .d(\DFF_717.D ),
    .q(\DFF_717.Q )
  );
  al_dffl _11382_ (
    .clk(CK),
    .d(\DFF_718.D ),
    .q(\DFF_718.Q )
  );
  al_dffl _11383_ (
    .clk(CK),
    .d(\DFF_719.D ),
    .q(\DFF_719.Q )
  );
  al_dffl _11384_ (
    .clk(CK),
    .d(\DFF_720.D ),
    .q(\DFF_720.Q )
  );
  al_dffl _11385_ (
    .clk(CK),
    .d(\DFF_721.D ),
    .q(\DFF_721.Q )
  );
  al_dffl _11386_ (
    .clk(CK),
    .d(\DFF_722.D ),
    .q(\DFF_722.Q )
  );
  al_dffl _11387_ (
    .clk(CK),
    .d(\DFF_723.D ),
    .q(\DFF_723.Q )
  );
  al_dffl _11388_ (
    .clk(CK),
    .d(\DFF_724.D ),
    .q(\DFF_724.Q )
  );
  al_dffl _11389_ (
    .clk(CK),
    .d(\DFF_725.D ),
    .q(\DFF_725.Q )
  );
  al_dffl _11390_ (
    .clk(CK),
    .d(\DFF_726.D ),
    .q(\DFF_726.Q )
  );
  al_dffl _11391_ (
    .clk(CK),
    .d(\DFF_727.D ),
    .q(\DFF_727.Q )
  );
  al_dffl _11392_ (
    .clk(CK),
    .d(\DFF_728.D ),
    .q(\DFF_728.Q )
  );
  al_dffl _11393_ (
    .clk(CK),
    .d(\DFF_729.D ),
    .q(\DFF_729.Q )
  );
  al_dffl _11394_ (
    .clk(CK),
    .d(\DFF_730.D ),
    .q(\DFF_730.Q )
  );
  al_dffl _11395_ (
    .clk(CK),
    .d(\DFF_731.D ),
    .q(\DFF_731.Q )
  );
  al_dffl _11396_ (
    .clk(CK),
    .d(\DFF_732.D ),
    .q(\DFF_732.Q )
  );
  al_dffl _11397_ (
    .clk(CK),
    .d(\DFF_733.D ),
    .q(\DFF_733.Q )
  );
  al_dffl _11398_ (
    .clk(CK),
    .d(\DFF_734.D ),
    .q(\DFF_734.Q )
  );
  al_dffl _11399_ (
    .clk(CK),
    .d(\DFF_735.D ),
    .q(\DFF_735.Q )
  );
  al_dffl _11400_ (
    .clk(CK),
    .d(\DFF_736.D ),
    .q(\DFF_736.Q )
  );
  al_dffl _11401_ (
    .clk(CK),
    .d(\DFF_737.D ),
    .q(\DFF_737.Q )
  );
  al_dffl _11402_ (
    .clk(CK),
    .d(\DFF_738.D ),
    .q(\DFF_738.Q )
  );
  al_dffl _11403_ (
    .clk(CK),
    .d(\DFF_739.D ),
    .q(\DFF_739.Q )
  );
  al_dffl _11404_ (
    .clk(CK),
    .d(\DFF_740.D ),
    .q(\DFF_740.Q )
  );
  al_dffl _11405_ (
    .clk(CK),
    .d(\DFF_741.D ),
    .q(\DFF_741.Q )
  );
  al_dffl _11406_ (
    .clk(CK),
    .d(\DFF_742.D ),
    .q(\DFF_742.Q )
  );
  al_dffl _11407_ (
    .clk(CK),
    .d(\DFF_743.D ),
    .q(\DFF_743.Q )
  );
  al_dffl _11408_ (
    .clk(CK),
    .d(\DFF_744.D ),
    .q(\DFF_744.Q )
  );
  al_dffl _11409_ (
    .clk(CK),
    .d(\DFF_745.D ),
    .q(\DFF_745.Q )
  );
  al_dffl _11410_ (
    .clk(CK),
    .d(\DFF_746.D ),
    .q(\DFF_746.Q )
  );
  al_dffl _11411_ (
    .clk(CK),
    .d(\DFF_747.D ),
    .q(\DFF_747.Q )
  );
  al_dffl _11412_ (
    .clk(CK),
    .d(\DFF_748.D ),
    .q(\DFF_748.Q )
  );
  al_dffl _11413_ (
    .clk(CK),
    .d(\DFF_749.D ),
    .q(\DFF_749.Q )
  );
  al_dffl _11414_ (
    .clk(CK),
    .d(\DFF_750.D ),
    .q(\DFF_750.Q )
  );
  al_dffl _11415_ (
    .clk(CK),
    .d(\DFF_751.D ),
    .q(\DFF_751.Q )
  );
  al_dffl _11416_ (
    .clk(CK),
    .d(\DFF_752.D ),
    .q(\DFF_752.Q )
  );
  al_dffl _11417_ (
    .clk(CK),
    .d(\DFF_753.D ),
    .q(\DFF_753.Q )
  );
  al_dffl _11418_ (
    .clk(CK),
    .d(\DFF_754.D ),
    .q(\DFF_754.Q )
  );
  al_dffl _11419_ (
    .clk(CK),
    .d(\DFF_755.D ),
    .q(\DFF_755.Q )
  );
  al_dffl _11420_ (
    .clk(CK),
    .d(\DFF_756.D ),
    .q(\DFF_756.Q )
  );
  al_dffl _11421_ (
    .clk(CK),
    .d(\DFF_757.D ),
    .q(\DFF_757.Q )
  );
  al_dffl _11422_ (
    .clk(CK),
    .d(\DFF_758.D ),
    .q(\DFF_758.Q )
  );
  al_dffl _11423_ (
    .clk(CK),
    .d(\DFF_759.D ),
    .q(\DFF_759.Q )
  );
  al_dffl _11424_ (
    .clk(CK),
    .d(\DFF_760.D ),
    .q(\DFF_760.Q )
  );
  al_dffl _11425_ (
    .clk(CK),
    .d(\DFF_761.D ),
    .q(\DFF_761.Q )
  );
  al_dffl _11426_ (
    .clk(CK),
    .d(\DFF_762.D ),
    .q(\DFF_762.Q )
  );
  al_dffl _11427_ (
    .clk(CK),
    .d(\DFF_763.D ),
    .q(\DFF_763.Q )
  );
  al_dffl _11428_ (
    .clk(CK),
    .d(\DFF_764.D ),
    .q(\DFF_764.Q )
  );
  al_dffl _11429_ (
    .clk(CK),
    .d(\DFF_765.D ),
    .q(\DFF_765.Q )
  );
  al_dffl _11430_ (
    .clk(CK),
    .d(\DFF_766.D ),
    .q(\DFF_766.Q )
  );
  al_dffl _11431_ (
    .clk(CK),
    .d(\DFF_767.D ),
    .q(\DFF_767.Q )
  );
  al_dffl _11432_ (
    .clk(CK),
    .d(\DFF_768.D ),
    .q(\DFF_768.Q )
  );
  al_dffl _11433_ (
    .clk(CK),
    .d(\DFF_769.D ),
    .q(\DFF_769.Q )
  );
  al_dffl _11434_ (
    .clk(CK),
    .d(\DFF_770.D ),
    .q(\DFF_770.Q )
  );
  al_dffl _11435_ (
    .clk(CK),
    .d(\DFF_771.D ),
    .q(\DFF_771.Q )
  );
  al_dffl _11436_ (
    .clk(CK),
    .d(\DFF_772.D ),
    .q(\DFF_772.Q )
  );
  al_dffl _11437_ (
    .clk(CK),
    .d(\DFF_773.D ),
    .q(\DFF_773.Q )
  );
  al_dffl _11438_ (
    .clk(CK),
    .d(\DFF_774.D ),
    .q(\DFF_774.Q )
  );
  al_dffl _11439_ (
    .clk(CK),
    .d(\DFF_775.D ),
    .q(\DFF_775.Q )
  );
  al_dffl _11440_ (
    .clk(CK),
    .d(\DFF_776.D ),
    .q(\DFF_776.Q )
  );
  al_dffl _11441_ (
    .clk(CK),
    .d(\DFF_777.D ),
    .q(\DFF_777.Q )
  );
  al_dffl _11442_ (
    .clk(CK),
    .d(\DFF_778.D ),
    .q(\DFF_778.Q )
  );
  al_dffl _11443_ (
    .clk(CK),
    .d(\DFF_779.D ),
    .q(\DFF_779.Q )
  );
  al_dffl _11444_ (
    .clk(CK),
    .d(\DFF_780.D ),
    .q(\DFF_780.Q )
  );
  al_dffl _11445_ (
    .clk(CK),
    .d(\DFF_781.D ),
    .q(\DFF_781.Q )
  );
  al_dffl _11446_ (
    .clk(CK),
    .d(\DFF_782.D ),
    .q(\DFF_782.Q )
  );
  al_dffl _11447_ (
    .clk(CK),
    .d(\DFF_783.D ),
    .q(\DFF_783.Q )
  );
  al_dffl _11448_ (
    .clk(CK),
    .d(\DFF_784.D ),
    .q(\DFF_784.Q )
  );
  al_dffl _11449_ (
    .clk(CK),
    .d(\DFF_785.D ),
    .q(\DFF_785.Q )
  );
  al_dffl _11450_ (
    .clk(CK),
    .d(\DFF_786.D ),
    .q(\DFF_786.Q )
  );
  al_dffl _11451_ (
    .clk(CK),
    .d(\DFF_787.D ),
    .q(\DFF_787.Q )
  );
  al_dffl _11452_ (
    .clk(CK),
    .d(\DFF_788.D ),
    .q(\DFF_788.Q )
  );
  al_dffl _11453_ (
    .clk(CK),
    .d(\DFF_789.D ),
    .q(\DFF_789.Q )
  );
  al_dffl _11454_ (
    .clk(CK),
    .d(\DFF_790.D ),
    .q(\DFF_790.Q )
  );
  al_dffl _11455_ (
    .clk(CK),
    .d(\DFF_791.D ),
    .q(\DFF_791.Q )
  );
  al_dffl _11456_ (
    .clk(CK),
    .d(\DFF_792.D ),
    .q(\DFF_792.Q )
  );
  al_dffl _11457_ (
    .clk(CK),
    .d(\DFF_793.D ),
    .q(\DFF_793.Q )
  );
  al_dffl _11458_ (
    .clk(CK),
    .d(\DFF_794.D ),
    .q(\DFF_794.Q )
  );
  al_dffl _11459_ (
    .clk(CK),
    .d(\DFF_795.D ),
    .q(\DFF_795.Q )
  );
  al_dffl _11460_ (
    .clk(CK),
    .d(\DFF_796.D ),
    .q(\DFF_796.Q )
  );
  al_dffl _11461_ (
    .clk(CK),
    .d(\DFF_797.D ),
    .q(\DFF_797.Q )
  );
  al_dffl _11462_ (
    .clk(CK),
    .d(\DFF_798.D ),
    .q(\DFF_798.Q )
  );
  al_dffl _11463_ (
    .clk(CK),
    .d(\DFF_799.D ),
    .q(\DFF_799.Q )
  );
  al_dffl _11464_ (
    .clk(CK),
    .d(\DFF_800.D ),
    .q(\DFF_800.Q )
  );
  al_dffl _11465_ (
    .clk(CK),
    .d(\DFF_801.D ),
    .q(\DFF_801.Q )
  );
  al_dffl _11466_ (
    .clk(CK),
    .d(\DFF_802.D ),
    .q(\DFF_802.Q )
  );
  al_dffl _11467_ (
    .clk(CK),
    .d(\DFF_803.D ),
    .q(\DFF_803.Q )
  );
  al_dffl _11468_ (
    .clk(CK),
    .d(\DFF_804.D ),
    .q(\DFF_804.Q )
  );
  al_dffl _11469_ (
    .clk(CK),
    .d(\DFF_805.D ),
    .q(\DFF_805.Q )
  );
  al_dffl _11470_ (
    .clk(CK),
    .d(\DFF_806.D ),
    .q(\DFF_806.Q )
  );
  al_dffl _11471_ (
    .clk(CK),
    .d(\DFF_807.D ),
    .q(\DFF_807.Q )
  );
  al_dffl _11472_ (
    .clk(CK),
    .d(\DFF_808.D ),
    .q(\DFF_808.Q )
  );
  al_dffl _11473_ (
    .clk(CK),
    .d(\DFF_809.D ),
    .q(\DFF_809.Q )
  );
  al_dffl _11474_ (
    .clk(CK),
    .d(\DFF_810.D ),
    .q(\DFF_810.Q )
  );
  al_dffl _11475_ (
    .clk(CK),
    .d(\DFF_811.D ),
    .q(\DFF_811.Q )
  );
  al_dffl _11476_ (
    .clk(CK),
    .d(\DFF_812.D ),
    .q(\DFF_812.Q )
  );
  al_dffl _11477_ (
    .clk(CK),
    .d(\DFF_813.D ),
    .q(\DFF_813.Q )
  );
  al_dffl _11478_ (
    .clk(CK),
    .d(\DFF_814.D ),
    .q(\DFF_814.Q )
  );
  al_dffl _11479_ (
    .clk(CK),
    .d(\DFF_815.D ),
    .q(\DFF_815.Q )
  );
  al_dffl _11480_ (
    .clk(CK),
    .d(\DFF_816.D ),
    .q(\DFF_816.Q )
  );
  al_dffl _11481_ (
    .clk(CK),
    .d(\DFF_817.D ),
    .q(\DFF_817.Q )
  );
  al_dffl _11482_ (
    .clk(CK),
    .d(\DFF_818.D ),
    .q(\DFF_818.Q )
  );
  al_dffl _11483_ (
    .clk(CK),
    .d(\DFF_819.D ),
    .q(\DFF_819.Q )
  );
  al_dffl _11484_ (
    .clk(CK),
    .d(\DFF_820.D ),
    .q(\DFF_820.Q )
  );
  al_dffl _11485_ (
    .clk(CK),
    .d(\DFF_821.D ),
    .q(\DFF_821.Q )
  );
  al_dffl _11486_ (
    .clk(CK),
    .d(\DFF_822.D ),
    .q(\DFF_822.Q )
  );
  al_dffl _11487_ (
    .clk(CK),
    .d(\DFF_823.D ),
    .q(\DFF_823.Q )
  );
  al_dffl _11488_ (
    .clk(CK),
    .d(\DFF_824.D ),
    .q(\DFF_824.Q )
  );
  al_dffl _11489_ (
    .clk(CK),
    .d(\DFF_825.D ),
    .q(\DFF_825.Q )
  );
  al_dffl _11490_ (
    .clk(CK),
    .d(\DFF_826.D ),
    .q(\DFF_826.Q )
  );
  al_dffl _11491_ (
    .clk(CK),
    .d(\DFF_827.D ),
    .q(\DFF_827.Q )
  );
  al_dffl _11492_ (
    .clk(CK),
    .d(\DFF_828.D ),
    .q(\DFF_828.Q )
  );
  al_dffl _11493_ (
    .clk(CK),
    .d(\DFF_829.D ),
    .q(\DFF_829.Q )
  );
  al_dffl _11494_ (
    .clk(CK),
    .d(\DFF_830.D ),
    .q(\DFF_830.Q )
  );
  al_dffl _11495_ (
    .clk(CK),
    .d(\DFF_831.D ),
    .q(\DFF_831.Q )
  );
  al_dffl _11496_ (
    .clk(CK),
    .d(\DFF_832.D ),
    .q(\DFF_832.Q )
  );
  al_dffl _11497_ (
    .clk(CK),
    .d(\DFF_833.D ),
    .q(\DFF_833.Q )
  );
  al_dffl _11498_ (
    .clk(CK),
    .d(\DFF_834.D ),
    .q(\DFF_834.Q )
  );
  al_dffl _11499_ (
    .clk(CK),
    .d(\DFF_835.D ),
    .q(\DFF_835.Q )
  );
  al_dffl _11500_ (
    .clk(CK),
    .d(\DFF_836.D ),
    .q(\DFF_836.Q )
  );
  al_dffl _11501_ (
    .clk(CK),
    .d(\DFF_837.D ),
    .q(\DFF_837.Q )
  );
  al_dffl _11502_ (
    .clk(CK),
    .d(\DFF_838.D ),
    .q(\DFF_838.Q )
  );
  al_dffl _11503_ (
    .clk(CK),
    .d(\DFF_839.D ),
    .q(\DFF_839.Q )
  );
  al_dffl _11504_ (
    .clk(CK),
    .d(\DFF_840.D ),
    .q(\DFF_840.Q )
  );
  al_dffl _11505_ (
    .clk(CK),
    .d(\DFF_841.D ),
    .q(\DFF_841.Q )
  );
  al_dffl _11506_ (
    .clk(CK),
    .d(\DFF_842.D ),
    .q(\DFF_842.Q )
  );
  al_dffl _11507_ (
    .clk(CK),
    .d(\DFF_843.D ),
    .q(\DFF_843.Q )
  );
  al_dffl _11508_ (
    .clk(CK),
    .d(\DFF_844.D ),
    .q(\DFF_844.Q )
  );
  al_dffl _11509_ (
    .clk(CK),
    .d(\DFF_845.D ),
    .q(\DFF_845.Q )
  );
  al_dffl _11510_ (
    .clk(CK),
    .d(\DFF_846.D ),
    .q(\DFF_846.Q )
  );
  al_dffl _11511_ (
    .clk(CK),
    .d(\DFF_847.D ),
    .q(\DFF_847.Q )
  );
  al_dffl _11512_ (
    .clk(CK),
    .d(\DFF_848.D ),
    .q(\DFF_848.Q )
  );
  al_dffl _11513_ (
    .clk(CK),
    .d(\DFF_849.D ),
    .q(\DFF_849.Q )
  );
  al_dffl _11514_ (
    .clk(CK),
    .d(\DFF_850.D ),
    .q(\DFF_850.Q )
  );
  al_dffl _11515_ (
    .clk(CK),
    .d(\DFF_851.D ),
    .q(\DFF_851.Q )
  );
  al_dffl _11516_ (
    .clk(CK),
    .d(\DFF_852.D ),
    .q(\DFF_852.Q )
  );
  al_dffl _11517_ (
    .clk(CK),
    .d(\DFF_853.D ),
    .q(\DFF_853.Q )
  );
  al_dffl _11518_ (
    .clk(CK),
    .d(\DFF_854.D ),
    .q(\DFF_854.Q )
  );
  al_dffl _11519_ (
    .clk(CK),
    .d(\DFF_855.D ),
    .q(\DFF_855.Q )
  );
  al_dffl _11520_ (
    .clk(CK),
    .d(\DFF_856.D ),
    .q(\DFF_856.Q )
  );
  al_dffl _11521_ (
    .clk(CK),
    .d(\DFF_857.D ),
    .q(\DFF_857.Q )
  );
  al_dffl _11522_ (
    .clk(CK),
    .d(\DFF_858.D ),
    .q(\DFF_858.Q )
  );
  al_dffl _11523_ (
    .clk(CK),
    .d(\DFF_859.D ),
    .q(\DFF_859.Q )
  );
  al_dffl _11524_ (
    .clk(CK),
    .d(\DFF_860.D ),
    .q(\DFF_860.Q )
  );
  al_dffl _11525_ (
    .clk(CK),
    .d(\DFF_861.D ),
    .q(\DFF_861.Q )
  );
  al_dffl _11526_ (
    .clk(CK),
    .d(\DFF_862.D ),
    .q(\DFF_862.Q )
  );
  al_dffl _11527_ (
    .clk(CK),
    .d(\DFF_863.D ),
    .q(\DFF_863.Q )
  );
  al_dffl _11528_ (
    .clk(CK),
    .d(\DFF_864.D ),
    .q(\DFF_864.Q )
  );
  al_dffl _11529_ (
    .clk(CK),
    .d(\DFF_865.D ),
    .q(\DFF_865.Q )
  );
  al_dffl _11530_ (
    .clk(CK),
    .d(\DFF_866.D ),
    .q(\DFF_866.Q )
  );
  al_dffl _11531_ (
    .clk(CK),
    .d(\DFF_867.D ),
    .q(\DFF_867.Q )
  );
  al_dffl _11532_ (
    .clk(CK),
    .d(\DFF_868.D ),
    .q(\DFF_868.Q )
  );
  al_dffl _11533_ (
    .clk(CK),
    .d(\DFF_869.D ),
    .q(\DFF_869.Q )
  );
  al_dffl _11534_ (
    .clk(CK),
    .d(\DFF_870.D ),
    .q(\DFF_870.Q )
  );
  al_dffl _11535_ (
    .clk(CK),
    .d(\DFF_871.D ),
    .q(\DFF_871.Q )
  );
  al_dffl _11536_ (
    .clk(CK),
    .d(\DFF_872.D ),
    .q(\DFF_872.Q )
  );
  al_dffl _11537_ (
    .clk(CK),
    .d(\DFF_873.D ),
    .q(\DFF_873.Q )
  );
  al_dffl _11538_ (
    .clk(CK),
    .d(\DFF_874.D ),
    .q(\DFF_874.Q )
  );
  al_dffl _11539_ (
    .clk(CK),
    .d(\DFF_875.D ),
    .q(\DFF_875.Q )
  );
  al_dffl _11540_ (
    .clk(CK),
    .d(\DFF_876.D ),
    .q(\DFF_876.Q )
  );
  al_dffl _11541_ (
    .clk(CK),
    .d(\DFF_877.D ),
    .q(\DFF_877.Q )
  );
  al_dffl _11542_ (
    .clk(CK),
    .d(\DFF_878.D ),
    .q(\DFF_878.Q )
  );
  al_dffl _11543_ (
    .clk(CK),
    .d(\DFF_879.D ),
    .q(\DFF_879.Q )
  );
  al_dffl _11544_ (
    .clk(CK),
    .d(\DFF_880.D ),
    .q(\DFF_880.Q )
  );
  al_dffl _11545_ (
    .clk(CK),
    .d(\DFF_881.D ),
    .q(\DFF_881.Q )
  );
  al_dffl _11546_ (
    .clk(CK),
    .d(\DFF_882.D ),
    .q(\DFF_882.Q )
  );
  al_dffl _11547_ (
    .clk(CK),
    .d(\DFF_883.D ),
    .q(\DFF_883.Q )
  );
  al_dffl _11548_ (
    .clk(CK),
    .d(\DFF_884.D ),
    .q(\DFF_884.Q )
  );
  al_dffl _11549_ (
    .clk(CK),
    .d(\DFF_885.D ),
    .q(\DFF_885.Q )
  );
  al_dffl _11550_ (
    .clk(CK),
    .d(\DFF_886.D ),
    .q(\DFF_886.Q )
  );
  al_dffl _11551_ (
    .clk(CK),
    .d(\DFF_887.D ),
    .q(\DFF_887.Q )
  );
  al_dffl _11552_ (
    .clk(CK),
    .d(\DFF_888.D ),
    .q(\DFF_888.Q )
  );
  al_dffl _11553_ (
    .clk(CK),
    .d(\DFF_889.D ),
    .q(\DFF_889.Q )
  );
  al_dffl _11554_ (
    .clk(CK),
    .d(\DFF_890.D ),
    .q(\DFF_890.Q )
  );
  al_dffl _11555_ (
    .clk(CK),
    .d(\DFF_891.D ),
    .q(\DFF_891.Q )
  );
  al_dffl _11556_ (
    .clk(CK),
    .d(\DFF_892.D ),
    .q(\DFF_892.Q )
  );
  al_dffl _11557_ (
    .clk(CK),
    .d(\DFF_893.D ),
    .q(\DFF_893.Q )
  );
  al_dffl _11558_ (
    .clk(CK),
    .d(\DFF_894.D ),
    .q(\DFF_894.Q )
  );
  al_dffl _11559_ (
    .clk(CK),
    .d(\DFF_895.D ),
    .q(\DFF_895.Q )
  );
  al_dffl _11560_ (
    .clk(CK),
    .d(\DFF_896.D ),
    .q(\DFF_896.Q )
  );
  al_dffl _11561_ (
    .clk(CK),
    .d(\DFF_897.D ),
    .q(\DFF_897.Q )
  );
  al_dffl _11562_ (
    .clk(CK),
    .d(\DFF_898.D ),
    .q(\DFF_898.Q )
  );
  al_dffl _11563_ (
    .clk(CK),
    .d(\DFF_899.D ),
    .q(\DFF_899.Q )
  );
  al_dffl _11564_ (
    .clk(CK),
    .d(\DFF_900.D ),
    .q(\DFF_900.Q )
  );
  al_dffl _11565_ (
    .clk(CK),
    .d(\DFF_901.D ),
    .q(\DFF_901.Q )
  );
  al_dffl _11566_ (
    .clk(CK),
    .d(\DFF_902.D ),
    .q(\DFF_902.Q )
  );
  al_dffl _11567_ (
    .clk(CK),
    .d(\DFF_903.D ),
    .q(\DFF_903.Q )
  );
  al_dffl _11568_ (
    .clk(CK),
    .d(\DFF_904.D ),
    .q(\DFF_904.Q )
  );
  al_dffl _11569_ (
    .clk(CK),
    .d(\DFF_905.D ),
    .q(\DFF_905.Q )
  );
  al_dffl _11570_ (
    .clk(CK),
    .d(\DFF_906.D ),
    .q(\DFF_906.Q )
  );
  al_dffl _11571_ (
    .clk(CK),
    .d(\DFF_907.D ),
    .q(\DFF_907.Q )
  );
  al_dffl _11572_ (
    .clk(CK),
    .d(\DFF_908.D ),
    .q(\DFF_908.Q )
  );
  al_dffl _11573_ (
    .clk(CK),
    .d(\DFF_909.D ),
    .q(\DFF_909.Q )
  );
  al_dffl _11574_ (
    .clk(CK),
    .d(\DFF_910.D ),
    .q(\DFF_910.Q )
  );
  al_dffl _11575_ (
    .clk(CK),
    .d(\DFF_911.D ),
    .q(\DFF_911.Q )
  );
  al_dffl _11576_ (
    .clk(CK),
    .d(\DFF_912.D ),
    .q(\DFF_912.Q )
  );
  al_dffl _11577_ (
    .clk(CK),
    .d(\DFF_913.D ),
    .q(\DFF_913.Q )
  );
  al_dffl _11578_ (
    .clk(CK),
    .d(\DFF_914.D ),
    .q(\DFF_914.Q )
  );
  al_dffl _11579_ (
    .clk(CK),
    .d(\DFF_915.D ),
    .q(\DFF_915.Q )
  );
  al_dffl _11580_ (
    .clk(CK),
    .d(\DFF_916.D ),
    .q(\DFF_916.Q )
  );
  al_dffl _11581_ (
    .clk(CK),
    .d(\DFF_917.D ),
    .q(\DFF_917.Q )
  );
  al_dffl _11582_ (
    .clk(CK),
    .d(\DFF_918.D ),
    .q(\DFF_918.Q )
  );
  al_dffl _11583_ (
    .clk(CK),
    .d(\DFF_919.D ),
    .q(\DFF_919.Q )
  );
  al_dffl _11584_ (
    .clk(CK),
    .d(\DFF_920.D ),
    .q(\DFF_920.Q )
  );
  al_dffl _11585_ (
    .clk(CK),
    .d(\DFF_921.D ),
    .q(\DFF_921.Q )
  );
  al_dffl _11586_ (
    .clk(CK),
    .d(\DFF_922.D ),
    .q(\DFF_922.Q )
  );
  al_dffl _11587_ (
    .clk(CK),
    .d(\DFF_923.D ),
    .q(\DFF_923.Q )
  );
  al_dffl _11588_ (
    .clk(CK),
    .d(\DFF_924.D ),
    .q(\DFF_924.Q )
  );
  al_dffl _11589_ (
    .clk(CK),
    .d(\DFF_925.D ),
    .q(\DFF_925.Q )
  );
  al_dffl _11590_ (
    .clk(CK),
    .d(\DFF_926.D ),
    .q(\DFF_926.Q )
  );
  al_dffl _11591_ (
    .clk(CK),
    .d(\DFF_927.D ),
    .q(\DFF_927.Q )
  );
  al_dffl _11592_ (
    .clk(CK),
    .d(\DFF_928.D ),
    .q(\DFF_928.Q )
  );
  al_dffl _11593_ (
    .clk(CK),
    .d(\DFF_929.D ),
    .q(\DFF_929.Q )
  );
  al_dffl _11594_ (
    .clk(CK),
    .d(\DFF_930.D ),
    .q(\DFF_930.Q )
  );
  al_dffl _11595_ (
    .clk(CK),
    .d(\DFF_931.D ),
    .q(\DFF_931.Q )
  );
  al_dffl _11596_ (
    .clk(CK),
    .d(\DFF_932.D ),
    .q(\DFF_932.Q )
  );
  al_dffl _11597_ (
    .clk(CK),
    .d(\DFF_933.D ),
    .q(\DFF_933.Q )
  );
  al_dffl _11598_ (
    .clk(CK),
    .d(\DFF_934.D ),
    .q(\DFF_934.Q )
  );
  al_dffl _11599_ (
    .clk(CK),
    .d(\DFF_935.D ),
    .q(\DFF_935.Q )
  );
  al_dffl _11600_ (
    .clk(CK),
    .d(\DFF_936.D ),
    .q(\DFF_936.Q )
  );
  al_dffl _11601_ (
    .clk(CK),
    .d(\DFF_937.D ),
    .q(\DFF_937.Q )
  );
  al_dffl _11602_ (
    .clk(CK),
    .d(\DFF_938.D ),
    .q(\DFF_938.Q )
  );
  al_dffl _11603_ (
    .clk(CK),
    .d(\DFF_939.D ),
    .q(\DFF_939.Q )
  );
  al_dffl _11604_ (
    .clk(CK),
    .d(\DFF_940.D ),
    .q(\DFF_940.Q )
  );
  al_dffl _11605_ (
    .clk(CK),
    .d(\DFF_941.D ),
    .q(\DFF_941.Q )
  );
  al_dffl _11606_ (
    .clk(CK),
    .d(\DFF_942.D ),
    .q(\DFF_942.Q )
  );
  al_dffl _11607_ (
    .clk(CK),
    .d(\DFF_943.D ),
    .q(\DFF_943.Q )
  );
  al_dffl _11608_ (
    .clk(CK),
    .d(\DFF_944.D ),
    .q(\DFF_944.Q )
  );
  al_dffl _11609_ (
    .clk(CK),
    .d(\DFF_945.D ),
    .q(\DFF_945.Q )
  );
  al_dffl _11610_ (
    .clk(CK),
    .d(\DFF_946.D ),
    .q(\DFF_946.Q )
  );
  al_dffl _11611_ (
    .clk(CK),
    .d(\DFF_947.D ),
    .q(\DFF_947.Q )
  );
  al_dffl _11612_ (
    .clk(CK),
    .d(\DFF_948.D ),
    .q(\DFF_948.Q )
  );
  al_dffl _11613_ (
    .clk(CK),
    .d(\DFF_949.D ),
    .q(\DFF_949.Q )
  );
  al_dffl _11614_ (
    .clk(CK),
    .d(\DFF_950.D ),
    .q(\DFF_950.Q )
  );
  al_dffl _11615_ (
    .clk(CK),
    .d(\DFF_951.D ),
    .q(\DFF_951.Q )
  );
  al_dffl _11616_ (
    .clk(CK),
    .d(\DFF_952.D ),
    .q(\DFF_952.Q )
  );
  al_dffl _11617_ (
    .clk(CK),
    .d(\DFF_953.D ),
    .q(\DFF_953.Q )
  );
  al_dffl _11618_ (
    .clk(CK),
    .d(\DFF_954.D ),
    .q(\DFF_954.Q )
  );
  al_dffl _11619_ (
    .clk(CK),
    .d(\DFF_955.D ),
    .q(\DFF_955.Q )
  );
  al_dffl _11620_ (
    .clk(CK),
    .d(\DFF_956.D ),
    .q(\DFF_956.Q )
  );
  al_dffl _11621_ (
    .clk(CK),
    .d(\DFF_957.D ),
    .q(\DFF_957.Q )
  );
  al_dffl _11622_ (
    .clk(CK),
    .d(\DFF_958.D ),
    .q(\DFF_958.Q )
  );
  al_dffl _11623_ (
    .clk(CK),
    .d(\DFF_959.D ),
    .q(\DFF_959.Q )
  );
  al_dffl _11624_ (
    .clk(CK),
    .d(\DFF_960.D ),
    .q(\DFF_960.Q )
  );
  al_dffl _11625_ (
    .clk(CK),
    .d(\DFF_961.D ),
    .q(\DFF_961.Q )
  );
  al_dffl _11626_ (
    .clk(CK),
    .d(\DFF_962.D ),
    .q(\DFF_962.Q )
  );
  al_dffl _11627_ (
    .clk(CK),
    .d(\DFF_963.D ),
    .q(\DFF_963.Q )
  );
  al_dffl _11628_ (
    .clk(CK),
    .d(\DFF_964.D ),
    .q(\DFF_964.Q )
  );
  al_dffl _11629_ (
    .clk(CK),
    .d(\DFF_965.D ),
    .q(\DFF_965.Q )
  );
  al_dffl _11630_ (
    .clk(CK),
    .d(\DFF_966.D ),
    .q(\DFF_966.Q )
  );
  al_dffl _11631_ (
    .clk(CK),
    .d(\DFF_967.D ),
    .q(\DFF_967.Q )
  );
  al_dffl _11632_ (
    .clk(CK),
    .d(\DFF_968.D ),
    .q(\DFF_968.Q )
  );
  al_dffl _11633_ (
    .clk(CK),
    .d(\DFF_969.D ),
    .q(\DFF_969.Q )
  );
  al_dffl _11634_ (
    .clk(CK),
    .d(\DFF_970.D ),
    .q(\DFF_970.Q )
  );
  al_dffl _11635_ (
    .clk(CK),
    .d(\DFF_971.D ),
    .q(\DFF_971.Q )
  );
  al_dffl _11636_ (
    .clk(CK),
    .d(\DFF_972.D ),
    .q(\DFF_972.Q )
  );
  al_dffl _11637_ (
    .clk(CK),
    .d(\DFF_973.D ),
    .q(\DFF_973.Q )
  );
  al_dffl _11638_ (
    .clk(CK),
    .d(\DFF_974.D ),
    .q(\DFF_974.Q )
  );
  al_dffl _11639_ (
    .clk(CK),
    .d(\DFF_975.D ),
    .q(\DFF_975.Q )
  );
  al_dffl _11640_ (
    .clk(CK),
    .d(\DFF_976.D ),
    .q(\DFF_976.Q )
  );
  al_dffl _11641_ (
    .clk(CK),
    .d(\DFF_977.D ),
    .q(\DFF_977.Q )
  );
  al_dffl _11642_ (
    .clk(CK),
    .d(\DFF_978.D ),
    .q(\DFF_978.Q )
  );
  al_dffl _11643_ (
    .clk(CK),
    .d(\DFF_979.D ),
    .q(\DFF_979.Q )
  );
  al_dffl _11644_ (
    .clk(CK),
    .d(\DFF_980.D ),
    .q(\DFF_980.Q )
  );
  al_dffl _11645_ (
    .clk(CK),
    .d(\DFF_981.D ),
    .q(\DFF_981.Q )
  );
  al_dffl _11646_ (
    .clk(CK),
    .d(\DFF_982.D ),
    .q(\DFF_982.Q )
  );
  al_dffl _11647_ (
    .clk(CK),
    .d(\DFF_983.D ),
    .q(\DFF_983.Q )
  );
  al_dffl _11648_ (
    .clk(CK),
    .d(\DFF_984.D ),
    .q(\DFF_984.Q )
  );
  al_dffl _11649_ (
    .clk(CK),
    .d(\DFF_985.D ),
    .q(\DFF_985.Q )
  );
  al_dffl _11650_ (
    .clk(CK),
    .d(\DFF_986.D ),
    .q(\DFF_986.Q )
  );
  al_dffl _11651_ (
    .clk(CK),
    .d(\DFF_987.D ),
    .q(\DFF_987.Q )
  );
  al_dffl _11652_ (
    .clk(CK),
    .d(\DFF_988.D ),
    .q(\DFF_988.Q )
  );
  al_dffl _11653_ (
    .clk(CK),
    .d(\DFF_989.D ),
    .q(\DFF_989.Q )
  );
  al_dffl _11654_ (
    .clk(CK),
    .d(\DFF_990.D ),
    .q(\DFF_990.Q )
  );
  al_dffl _11655_ (
    .clk(CK),
    .d(\DFF_991.D ),
    .q(\DFF_991.Q )
  );
  al_dffl _11656_ (
    .clk(CK),
    .d(\DFF_992.D ),
    .q(\DFF_992.Q )
  );
  al_dffl _11657_ (
    .clk(CK),
    .d(\DFF_993.D ),
    .q(\DFF_993.Q )
  );
  al_dffl _11658_ (
    .clk(CK),
    .d(\DFF_994.D ),
    .q(\DFF_994.Q )
  );
  al_dffl _11659_ (
    .clk(CK),
    .d(\DFF_995.D ),
    .q(\DFF_995.Q )
  );
  al_dffl _11660_ (
    .clk(CK),
    .d(\DFF_996.D ),
    .q(\DFF_996.Q )
  );
  al_dffl _11661_ (
    .clk(CK),
    .d(\DFF_997.D ),
    .q(\DFF_997.Q )
  );
  al_dffl _11662_ (
    .clk(CK),
    .d(\DFF_998.D ),
    .q(\DFF_998.Q )
  );
  al_dffl _11663_ (
    .clk(CK),
    .d(\DFF_999.D ),
    .q(\DFF_999.Q )
  );
  al_dffl _11664_ (
    .clk(CK),
    .d(\DFF_1000.D ),
    .q(\DFF_1000.Q )
  );
  al_dffl _11665_ (
    .clk(CK),
    .d(\DFF_1001.D ),
    .q(\DFF_1001.Q )
  );
  al_dffl _11666_ (
    .clk(CK),
    .d(\DFF_1002.D ),
    .q(\DFF_1002.Q )
  );
  al_dffl _11667_ (
    .clk(CK),
    .d(\DFF_1003.D ),
    .q(\DFF_1003.Q )
  );
  al_dffl _11668_ (
    .clk(CK),
    .d(\DFF_1004.D ),
    .q(\DFF_1004.Q )
  );
  al_dffl _11669_ (
    .clk(CK),
    .d(\DFF_1005.D ),
    .q(\DFF_1005.Q )
  );
  al_dffl _11670_ (
    .clk(CK),
    .d(\DFF_1006.D ),
    .q(\DFF_1006.Q )
  );
  al_dffl _11671_ (
    .clk(CK),
    .d(\DFF_1007.D ),
    .q(\DFF_1007.Q )
  );
  al_dffl _11672_ (
    .clk(CK),
    .d(\DFF_1008.D ),
    .q(\DFF_1008.Q )
  );
  al_dffl _11673_ (
    .clk(CK),
    .d(\DFF_1009.D ),
    .q(\DFF_1009.Q )
  );
  al_dffl _11674_ (
    .clk(CK),
    .d(\DFF_1010.D ),
    .q(\DFF_1010.Q )
  );
  al_dffl _11675_ (
    .clk(CK),
    .d(\DFF_1011.D ),
    .q(\DFF_1011.Q )
  );
  al_dffl _11676_ (
    .clk(CK),
    .d(\DFF_1012.D ),
    .q(\DFF_1012.Q )
  );
  al_dffl _11677_ (
    .clk(CK),
    .d(\DFF_1013.D ),
    .q(\DFF_1013.Q )
  );
  al_dffl _11678_ (
    .clk(CK),
    .d(\DFF_1014.D ),
    .q(\DFF_1014.Q )
  );
  al_dffl _11679_ (
    .clk(CK),
    .d(\DFF_1015.D ),
    .q(\DFF_1015.Q )
  );
  al_dffl _11680_ (
    .clk(CK),
    .d(\DFF_1016.D ),
    .q(\DFF_1016.Q )
  );
  al_dffl _11681_ (
    .clk(CK),
    .d(\DFF_1017.D ),
    .q(\DFF_1017.Q )
  );
  al_dffl _11682_ (
    .clk(CK),
    .d(\DFF_1018.D ),
    .q(\DFF_1018.Q )
  );
  al_dffl _11683_ (
    .clk(CK),
    .d(\DFF_1019.D ),
    .q(\DFF_1019.Q )
  );
  al_dffl _11684_ (
    .clk(CK),
    .d(\DFF_1020.D ),
    .q(\DFF_1020.Q )
  );
  al_dffl _11685_ (
    .clk(CK),
    .d(\DFF_1021.D ),
    .q(\DFF_1021.Q )
  );
  al_dffl _11686_ (
    .clk(CK),
    .d(\DFF_1022.D ),
    .q(\DFF_1022.Q )
  );
  al_dffl _11687_ (
    .clk(CK),
    .d(\DFF_1023.D ),
    .q(\DFF_1023.Q )
  );
  al_dffl _11688_ (
    .clk(CK),
    .d(\DFF_1024.D ),
    .q(\DFF_1024.Q )
  );
  al_dffl _11689_ (
    .clk(CK),
    .d(\DFF_1025.D ),
    .q(\DFF_1025.Q )
  );
  al_dffl _11690_ (
    .clk(CK),
    .d(\DFF_1026.D ),
    .q(\DFF_1026.Q )
  );
  al_dffl _11691_ (
    .clk(CK),
    .d(\DFF_1027.D ),
    .q(\DFF_1027.Q )
  );
  al_dffl _11692_ (
    .clk(CK),
    .d(\DFF_1028.D ),
    .q(\DFF_1028.Q )
  );
  al_dffl _11693_ (
    .clk(CK),
    .d(\DFF_1029.D ),
    .q(\DFF_1029.Q )
  );
  al_dffl _11694_ (
    .clk(CK),
    .d(\DFF_1030.D ),
    .q(\DFF_1030.Q )
  );
  al_dffl _11695_ (
    .clk(CK),
    .d(\DFF_1031.D ),
    .q(\DFF_1031.Q )
  );
  al_dffl _11696_ (
    .clk(CK),
    .d(\DFF_1032.D ),
    .q(\DFF_1032.Q )
  );
  al_dffl _11697_ (
    .clk(CK),
    .d(\DFF_1033.D ),
    .q(\DFF_1033.Q )
  );
  al_dffl _11698_ (
    .clk(CK),
    .d(\DFF_1034.D ),
    .q(\DFF_1034.Q )
  );
  al_dffl _11699_ (
    .clk(CK),
    .d(\DFF_1035.D ),
    .q(\DFF_1035.Q )
  );
  al_dffl _11700_ (
    .clk(CK),
    .d(\DFF_1036.D ),
    .q(\DFF_1036.Q )
  );
  al_dffl _11701_ (
    .clk(CK),
    .d(\DFF_1037.D ),
    .q(\DFF_1037.Q )
  );
  al_dffl _11702_ (
    .clk(CK),
    .d(\DFF_1038.D ),
    .q(\DFF_1038.Q )
  );
  al_dffl _11703_ (
    .clk(CK),
    .d(\DFF_1039.D ),
    .q(\DFF_1039.Q )
  );
  al_dffl _11704_ (
    .clk(CK),
    .d(\DFF_1040.D ),
    .q(\DFF_1040.Q )
  );
  al_dffl _11705_ (
    .clk(CK),
    .d(\DFF_1041.D ),
    .q(\DFF_1041.Q )
  );
  al_dffl _11706_ (
    .clk(CK),
    .d(\DFF_1042.D ),
    .q(\DFF_1042.Q )
  );
  al_dffl _11707_ (
    .clk(CK),
    .d(\DFF_1043.D ),
    .q(\DFF_1043.Q )
  );
  al_dffl _11708_ (
    .clk(CK),
    .d(\DFF_1044.D ),
    .q(\DFF_1044.Q )
  );
  al_dffl _11709_ (
    .clk(CK),
    .d(\DFF_1045.D ),
    .q(\DFF_1045.Q )
  );
  al_dffl _11710_ (
    .clk(CK),
    .d(\DFF_1046.D ),
    .q(\DFF_1046.Q )
  );
  al_dffl _11711_ (
    .clk(CK),
    .d(\DFF_1047.D ),
    .q(\DFF_1047.Q )
  );
  al_dffl _11712_ (
    .clk(CK),
    .d(\DFF_1048.D ),
    .q(\DFF_1048.Q )
  );
  al_dffl _11713_ (
    .clk(CK),
    .d(\DFF_1049.D ),
    .q(\DFF_1049.Q )
  );
  al_dffl _11714_ (
    .clk(CK),
    .d(\DFF_1050.D ),
    .q(\DFF_1050.Q )
  );
  al_dffl _11715_ (
    .clk(CK),
    .d(\DFF_1051.D ),
    .q(\DFF_1051.Q )
  );
  al_dffl _11716_ (
    .clk(CK),
    .d(\DFF_1052.D ),
    .q(\DFF_1052.Q )
  );
  al_dffl _11717_ (
    .clk(CK),
    .d(\DFF_1053.D ),
    .q(\DFF_1053.Q )
  );
  al_dffl _11718_ (
    .clk(CK),
    .d(\DFF_1054.D ),
    .q(\DFF_1054.Q )
  );
  al_dffl _11719_ (
    .clk(CK),
    .d(\DFF_1055.D ),
    .q(\DFF_1055.Q )
  );
  al_dffl _11720_ (
    .clk(CK),
    .d(\DFF_1056.D ),
    .q(\DFF_1056.Q )
  );
  al_dffl _11721_ (
    .clk(CK),
    .d(\DFF_1057.D ),
    .q(\DFF_1057.Q )
  );
  al_dffl _11722_ (
    .clk(CK),
    .d(\DFF_1058.D ),
    .q(\DFF_1058.Q )
  );
  al_dffl _11723_ (
    .clk(CK),
    .d(\DFF_1059.D ),
    .q(\DFF_1059.Q )
  );
  al_dffl _11724_ (
    .clk(CK),
    .d(\DFF_1060.D ),
    .q(\DFF_1060.Q )
  );
  al_dffl _11725_ (
    .clk(CK),
    .d(\DFF_1061.D ),
    .q(\DFF_1061.Q )
  );
  al_dffl _11726_ (
    .clk(CK),
    .d(\DFF_1062.D ),
    .q(\DFF_1062.Q )
  );
  al_dffl _11727_ (
    .clk(CK),
    .d(\DFF_1063.D ),
    .q(\DFF_1063.Q )
  );
  al_dffl _11728_ (
    .clk(CK),
    .d(\DFF_1064.D ),
    .q(\DFF_1064.Q )
  );
  al_dffl _11729_ (
    .clk(CK),
    .d(\DFF_1065.D ),
    .q(\DFF_1065.Q )
  );
  al_dffl _11730_ (
    .clk(CK),
    .d(\DFF_1066.D ),
    .q(\DFF_1066.Q )
  );
  al_dffl _11731_ (
    .clk(CK),
    .d(\DFF_1067.D ),
    .q(\DFF_1067.Q )
  );
  al_dffl _11732_ (
    .clk(CK),
    .d(\DFF_1068.D ),
    .q(\DFF_1068.Q )
  );
  al_dffl _11733_ (
    .clk(CK),
    .d(\DFF_1069.D ),
    .q(\DFF_1069.Q )
  );
  al_dffl _11734_ (
    .clk(CK),
    .d(\DFF_1070.D ),
    .q(\DFF_1070.Q )
  );
  al_dffl _11735_ (
    .clk(CK),
    .d(\DFF_1071.D ),
    .q(\DFF_1071.Q )
  );
  al_dffl _11736_ (
    .clk(CK),
    .d(\DFF_1072.D ),
    .q(\DFF_1072.Q )
  );
  al_dffl _11737_ (
    .clk(CK),
    .d(\DFF_1073.D ),
    .q(\DFF_1073.Q )
  );
  al_dffl _11738_ (
    .clk(CK),
    .d(\DFF_1074.D ),
    .q(\DFF_1074.Q )
  );
  al_dffl _11739_ (
    .clk(CK),
    .d(\DFF_1075.D ),
    .q(\DFF_1075.Q )
  );
  al_dffl _11740_ (
    .clk(CK),
    .d(\DFF_1076.D ),
    .q(\DFF_1076.Q )
  );
  al_dffl _11741_ (
    .clk(CK),
    .d(\DFF_1077.D ),
    .q(\DFF_1077.Q )
  );
  al_dffl _11742_ (
    .clk(CK),
    .d(\DFF_1078.D ),
    .q(\DFF_1078.Q )
  );
  al_dffl _11743_ (
    .clk(CK),
    .d(\DFF_1079.D ),
    .q(\DFF_1079.Q )
  );
  al_dffl _11744_ (
    .clk(CK),
    .d(\DFF_1080.D ),
    .q(\DFF_1080.Q )
  );
  al_dffl _11745_ (
    .clk(CK),
    .d(\DFF_1081.D ),
    .q(\DFF_1081.Q )
  );
  al_dffl _11746_ (
    .clk(CK),
    .d(\DFF_1082.D ),
    .q(\DFF_1082.Q )
  );
  al_dffl _11747_ (
    .clk(CK),
    .d(\DFF_1083.D ),
    .q(\DFF_1083.Q )
  );
  al_dffl _11748_ (
    .clk(CK),
    .d(\DFF_1084.D ),
    .q(\DFF_1084.Q )
  );
  al_dffl _11749_ (
    .clk(CK),
    .d(\DFF_1085.D ),
    .q(\DFF_1085.Q )
  );
  al_dffl _11750_ (
    .clk(CK),
    .d(\DFF_1086.D ),
    .q(\DFF_1086.Q )
  );
  al_dffl _11751_ (
    .clk(CK),
    .d(\DFF_1087.D ),
    .q(\DFF_1087.Q )
  );
  al_dffl _11752_ (
    .clk(CK),
    .d(\DFF_1088.D ),
    .q(\DFF_1088.Q )
  );
  al_dffl _11753_ (
    .clk(CK),
    .d(\DFF_1089.D ),
    .q(\DFF_1089.Q )
  );
  al_dffl _11754_ (
    .clk(CK),
    .d(\DFF_1090.D ),
    .q(\DFF_1090.Q )
  );
  al_dffl _11755_ (
    .clk(CK),
    .d(\DFF_1091.D ),
    .q(\DFF_1091.Q )
  );
  al_dffl _11756_ (
    .clk(CK),
    .d(\DFF_1092.D ),
    .q(\DFF_1092.Q )
  );
  al_dffl _11757_ (
    .clk(CK),
    .d(\DFF_1093.D ),
    .q(\DFF_1093.Q )
  );
  al_dffl _11758_ (
    .clk(CK),
    .d(\DFF_1094.D ),
    .q(\DFF_1094.Q )
  );
  al_dffl _11759_ (
    .clk(CK),
    .d(\DFF_1095.D ),
    .q(\DFF_1095.Q )
  );
  al_dffl _11760_ (
    .clk(CK),
    .d(\DFF_1096.D ),
    .q(\DFF_1096.Q )
  );
  al_dffl _11761_ (
    .clk(CK),
    .d(\DFF_1097.D ),
    .q(\DFF_1097.Q )
  );
  al_dffl _11762_ (
    .clk(CK),
    .d(\DFF_1098.D ),
    .q(\DFF_1098.Q )
  );
  al_dffl _11763_ (
    .clk(CK),
    .d(\DFF_1099.D ),
    .q(\DFF_1099.Q )
  );
  al_dffl _11764_ (
    .clk(CK),
    .d(\DFF_1100.D ),
    .q(\DFF_1100.Q )
  );
  al_dffl _11765_ (
    .clk(CK),
    .d(\DFF_1101.D ),
    .q(\DFF_1101.Q )
  );
  al_dffl _11766_ (
    .clk(CK),
    .d(\DFF_1102.D ),
    .q(\DFF_1102.Q )
  );
  al_dffl _11767_ (
    .clk(CK),
    .d(\DFF_1103.D ),
    .q(\DFF_1103.Q )
  );
  al_dffl _11768_ (
    .clk(CK),
    .d(\DFF_1104.D ),
    .q(\DFF_1104.Q )
  );
  al_dffl _11769_ (
    .clk(CK),
    .d(\DFF_1105.D ),
    .q(\DFF_1105.Q )
  );
  al_dffl _11770_ (
    .clk(CK),
    .d(\DFF_1106.D ),
    .q(\DFF_1106.Q )
  );
  al_dffl _11771_ (
    .clk(CK),
    .d(\DFF_1107.D ),
    .q(\DFF_1107.Q )
  );
  al_dffl _11772_ (
    .clk(CK),
    .d(\DFF_1108.D ),
    .q(\DFF_1108.Q )
  );
  al_dffl _11773_ (
    .clk(CK),
    .d(\DFF_1109.D ),
    .q(\DFF_1109.Q )
  );
  al_dffl _11774_ (
    .clk(CK),
    .d(\DFF_1110.D ),
    .q(\DFF_1110.Q )
  );
  al_dffl _11775_ (
    .clk(CK),
    .d(\DFF_1111.D ),
    .q(\DFF_1111.Q )
  );
  al_dffl _11776_ (
    .clk(CK),
    .d(\DFF_1112.D ),
    .q(\DFF_1112.Q )
  );
  al_dffl _11777_ (
    .clk(CK),
    .d(\DFF_1113.D ),
    .q(\DFF_1113.Q )
  );
  al_dffl _11778_ (
    .clk(CK),
    .d(\DFF_1114.D ),
    .q(\DFF_1114.Q )
  );
  al_dffl _11779_ (
    .clk(CK),
    .d(\DFF_1115.D ),
    .q(\DFF_1115.Q )
  );
  al_dffl _11780_ (
    .clk(CK),
    .d(\DFF_1116.D ),
    .q(\DFF_1116.Q )
  );
  al_dffl _11781_ (
    .clk(CK),
    .d(\DFF_1117.D ),
    .q(\DFF_1117.Q )
  );
  al_dffl _11782_ (
    .clk(CK),
    .d(\DFF_1118.D ),
    .q(\DFF_1118.Q )
  );
  al_dffl _11783_ (
    .clk(CK),
    .d(\DFF_1119.D ),
    .q(\DFF_1119.Q )
  );
  al_dffl _11784_ (
    .clk(CK),
    .d(\DFF_1120.D ),
    .q(\DFF_1120.Q )
  );
  al_dffl _11785_ (
    .clk(CK),
    .d(\DFF_1121.D ),
    .q(\DFF_1121.Q )
  );
  al_dffl _11786_ (
    .clk(CK),
    .d(\DFF_1122.D ),
    .q(\DFF_1122.Q )
  );
  al_dffl _11787_ (
    .clk(CK),
    .d(\DFF_1123.D ),
    .q(\DFF_1123.Q )
  );
  al_dffl _11788_ (
    .clk(CK),
    .d(\DFF_1124.D ),
    .q(\DFF_1124.Q )
  );
  al_dffl _11789_ (
    .clk(CK),
    .d(\DFF_1125.D ),
    .q(\DFF_1125.Q )
  );
  al_dffl _11790_ (
    .clk(CK),
    .d(\DFF_1126.D ),
    .q(\DFF_1126.Q )
  );
  al_dffl _11791_ (
    .clk(CK),
    .d(\DFF_1127.D ),
    .q(\DFF_1127.Q )
  );
  al_dffl _11792_ (
    .clk(CK),
    .d(\DFF_1128.D ),
    .q(\DFF_1128.Q )
  );
  al_dffl _11793_ (
    .clk(CK),
    .d(\DFF_1129.D ),
    .q(\DFF_1129.Q )
  );
  al_dffl _11794_ (
    .clk(CK),
    .d(\DFF_1130.D ),
    .q(\DFF_1130.Q )
  );
  al_dffl _11795_ (
    .clk(CK),
    .d(\DFF_1131.D ),
    .q(\DFF_1131.Q )
  );
  al_dffl _11796_ (
    .clk(CK),
    .d(\DFF_1132.D ),
    .q(\DFF_1132.Q )
  );
  al_dffl _11797_ (
    .clk(CK),
    .d(\DFF_1133.D ),
    .q(\DFF_1133.Q )
  );
  al_dffl _11798_ (
    .clk(CK),
    .d(\DFF_1134.D ),
    .q(\DFF_1134.Q )
  );
  al_dffl _11799_ (
    .clk(CK),
    .d(\DFF_1135.D ),
    .q(\DFF_1135.Q )
  );
  al_dffl _11800_ (
    .clk(CK),
    .d(\DFF_1136.D ),
    .q(\DFF_1136.Q )
  );
  al_dffl _11801_ (
    .clk(CK),
    .d(\DFF_1137.D ),
    .q(\DFF_1137.Q )
  );
  al_dffl _11802_ (
    .clk(CK),
    .d(\DFF_1138.D ),
    .q(\DFF_1138.Q )
  );
  al_dffl _11803_ (
    .clk(CK),
    .d(\DFF_1139.D ),
    .q(\DFF_1139.Q )
  );
  al_dffl _11804_ (
    .clk(CK),
    .d(\DFF_1140.D ),
    .q(\DFF_1140.Q )
  );
  al_dffl _11805_ (
    .clk(CK),
    .d(\DFF_1141.D ),
    .q(\DFF_1141.Q )
  );
  al_dffl _11806_ (
    .clk(CK),
    .d(\DFF_1142.D ),
    .q(\DFF_1142.Q )
  );
  al_dffl _11807_ (
    .clk(CK),
    .d(\DFF_1143.D ),
    .q(\DFF_1143.Q )
  );
  al_dffl _11808_ (
    .clk(CK),
    .d(\DFF_1144.D ),
    .q(\DFF_1144.Q )
  );
  al_dffl _11809_ (
    .clk(CK),
    .d(\DFF_1145.D ),
    .q(\DFF_1145.Q )
  );
  al_dffl _11810_ (
    .clk(CK),
    .d(\DFF_1146.D ),
    .q(\DFF_1146.Q )
  );
  al_dffl _11811_ (
    .clk(CK),
    .d(\DFF_1147.D ),
    .q(\DFF_1147.Q )
  );
  al_dffl _11812_ (
    .clk(CK),
    .d(\DFF_1148.D ),
    .q(\DFF_1148.Q )
  );
  al_dffl _11813_ (
    .clk(CK),
    .d(\DFF_1149.D ),
    .q(\DFF_1149.Q )
  );
  al_dffl _11814_ (
    .clk(CK),
    .d(\DFF_1150.D ),
    .q(\DFF_1150.Q )
  );
  al_dffl _11815_ (
    .clk(CK),
    .d(\DFF_1151.D ),
    .q(\DFF_1151.Q )
  );
  al_dffl _11816_ (
    .clk(CK),
    .d(\DFF_1152.D ),
    .q(\DFF_1152.Q )
  );
  al_dffl _11817_ (
    .clk(CK),
    .d(\DFF_1153.D ),
    .q(\DFF_1153.Q )
  );
  al_dffl _11818_ (
    .clk(CK),
    .d(\DFF_1154.D ),
    .q(\DFF_1154.Q )
  );
  al_dffl _11819_ (
    .clk(CK),
    .d(\DFF_1155.D ),
    .q(\DFF_1155.Q )
  );
  al_dffl _11820_ (
    .clk(CK),
    .d(\DFF_1156.D ),
    .q(\DFF_1156.Q )
  );
  al_dffl _11821_ (
    .clk(CK),
    .d(\DFF_1157.D ),
    .q(\DFF_1157.Q )
  );
  al_dffl _11822_ (
    .clk(CK),
    .d(\DFF_1158.D ),
    .q(\DFF_1158.Q )
  );
  al_dffl _11823_ (
    .clk(CK),
    .d(\DFF_1159.D ),
    .q(\DFF_1159.Q )
  );
  al_dffl _11824_ (
    .clk(CK),
    .d(\DFF_1160.D ),
    .q(\DFF_1160.Q )
  );
  al_dffl _11825_ (
    .clk(CK),
    .d(\DFF_1161.D ),
    .q(\DFF_1161.Q )
  );
  al_dffl _11826_ (
    .clk(CK),
    .d(\DFF_1162.D ),
    .q(\DFF_1162.Q )
  );
  al_dffl _11827_ (
    .clk(CK),
    .d(\DFF_1163.D ),
    .q(\DFF_1163.Q )
  );
  al_dffl _11828_ (
    .clk(CK),
    .d(\DFF_1164.D ),
    .q(\DFF_1164.Q )
  );
  al_dffl _11829_ (
    .clk(CK),
    .d(\DFF_1165.D ),
    .q(\DFF_1165.Q )
  );
  al_dffl _11830_ (
    .clk(CK),
    .d(\DFF_1166.D ),
    .q(\DFF_1166.Q )
  );
  al_dffl _11831_ (
    .clk(CK),
    .d(\DFF_1167.D ),
    .q(\DFF_1167.Q )
  );
  al_dffl _11832_ (
    .clk(CK),
    .d(\DFF_1168.D ),
    .q(\DFF_1168.Q )
  );
  al_dffl _11833_ (
    .clk(CK),
    .d(\DFF_1169.D ),
    .q(\DFF_1169.Q )
  );
  al_dffl _11834_ (
    .clk(CK),
    .d(\DFF_1170.D ),
    .q(\DFF_1170.Q )
  );
  al_dffl _11835_ (
    .clk(CK),
    .d(\DFF_1171.D ),
    .q(\DFF_1171.Q )
  );
  al_dffl _11836_ (
    .clk(CK),
    .d(\DFF_1172.D ),
    .q(\DFF_1172.Q )
  );
  al_dffl _11837_ (
    .clk(CK),
    .d(\DFF_1173.D ),
    .q(\DFF_1173.Q )
  );
  al_dffl _11838_ (
    .clk(CK),
    .d(\DFF_1174.D ),
    .q(\DFF_1174.Q )
  );
  al_dffl _11839_ (
    .clk(CK),
    .d(\DFF_1175.D ),
    .q(\DFF_1175.Q )
  );
  al_dffl _11840_ (
    .clk(CK),
    .d(\DFF_1176.D ),
    .q(\DFF_1176.Q )
  );
  al_dffl _11841_ (
    .clk(CK),
    .d(\DFF_1177.D ),
    .q(\DFF_1177.Q )
  );
  al_dffl _11842_ (
    .clk(CK),
    .d(\DFF_1178.D ),
    .q(\DFF_1178.Q )
  );
  al_dffl _11843_ (
    .clk(CK),
    .d(\DFF_1179.D ),
    .q(\DFF_1179.Q )
  );
  al_dffl _11844_ (
    .clk(CK),
    .d(\DFF_1180.D ),
    .q(\DFF_1180.Q )
  );
  al_dffl _11845_ (
    .clk(CK),
    .d(\DFF_1181.D ),
    .q(\DFF_1181.Q )
  );
  al_dffl _11846_ (
    .clk(CK),
    .d(\DFF_1182.D ),
    .q(\DFF_1182.Q )
  );
  al_dffl _11847_ (
    .clk(CK),
    .d(\DFF_1183.D ),
    .q(\DFF_1183.Q )
  );
  al_dffl _11848_ (
    .clk(CK),
    .d(\DFF_1184.D ),
    .q(\DFF_1184.Q )
  );
  al_dffl _11849_ (
    .clk(CK),
    .d(\DFF_1185.D ),
    .q(\DFF_1185.Q )
  );
  al_dffl _11850_ (
    .clk(CK),
    .d(\DFF_1186.D ),
    .q(\DFF_1186.Q )
  );
  al_dffl _11851_ (
    .clk(CK),
    .d(\DFF_1187.D ),
    .q(\DFF_1187.Q )
  );
  al_dffl _11852_ (
    .clk(CK),
    .d(\DFF_1188.D ),
    .q(\DFF_1188.Q )
  );
  al_dffl _11853_ (
    .clk(CK),
    .d(\DFF_1189.D ),
    .q(\DFF_1189.Q )
  );
  al_dffl _11854_ (
    .clk(CK),
    .d(\DFF_1190.D ),
    .q(\DFF_1190.Q )
  );
  al_dffl _11855_ (
    .clk(CK),
    .d(\DFF_1191.D ),
    .q(\DFF_1191.Q )
  );
  al_dffl _11856_ (
    .clk(CK),
    .d(\DFF_1192.D ),
    .q(\DFF_1192.Q )
  );
  al_dffl _11857_ (
    .clk(CK),
    .d(\DFF_1193.D ),
    .q(\DFF_1193.Q )
  );
  al_dffl _11858_ (
    .clk(CK),
    .d(\DFF_1194.D ),
    .q(\DFF_1194.Q )
  );
  al_dffl _11859_ (
    .clk(CK),
    .d(\DFF_1195.D ),
    .q(\DFF_1195.Q )
  );
  al_dffl _11860_ (
    .clk(CK),
    .d(\DFF_1196.D ),
    .q(\DFF_1196.Q )
  );
  al_dffl _11861_ (
    .clk(CK),
    .d(\DFF_1197.D ),
    .q(\DFF_1197.Q )
  );
  al_dffl _11862_ (
    .clk(CK),
    .d(\DFF_1198.D ),
    .q(\DFF_1198.Q )
  );
  al_dffl _11863_ (
    .clk(CK),
    .d(\DFF_1199.D ),
    .q(\DFF_1199.Q )
  );
  al_dffl _11864_ (
    .clk(CK),
    .d(\DFF_1200.D ),
    .q(\DFF_1200.Q )
  );
  al_dffl _11865_ (
    .clk(CK),
    .d(\DFF_1201.D ),
    .q(\DFF_1201.Q )
  );
  al_dffl _11866_ (
    .clk(CK),
    .d(\DFF_1202.D ),
    .q(\DFF_1202.Q )
  );
  al_dffl _11867_ (
    .clk(CK),
    .d(\DFF_1203.D ),
    .q(\DFF_1203.Q )
  );
  al_dffl _11868_ (
    .clk(CK),
    .d(\DFF_1204.D ),
    .q(\DFF_1204.Q )
  );
  al_dffl _11869_ (
    .clk(CK),
    .d(\DFF_1205.D ),
    .q(\DFF_1205.Q )
  );
  al_dffl _11870_ (
    .clk(CK),
    .d(\DFF_1206.D ),
    .q(\DFF_1206.Q )
  );
  al_dffl _11871_ (
    .clk(CK),
    .d(\DFF_1207.D ),
    .q(\DFF_1207.Q )
  );
  al_dffl _11872_ (
    .clk(CK),
    .d(\DFF_1208.D ),
    .q(\DFF_1208.Q )
  );
  al_dffl _11873_ (
    .clk(CK),
    .d(\DFF_1209.D ),
    .q(\DFF_1209.Q )
  );
  al_dffl _11874_ (
    .clk(CK),
    .d(\DFF_1210.D ),
    .q(\DFF_1210.Q )
  );
  al_dffl _11875_ (
    .clk(CK),
    .d(\DFF_1211.D ),
    .q(\DFF_1211.Q )
  );
  al_dffl _11876_ (
    .clk(CK),
    .d(\DFF_1212.D ),
    .q(\DFF_1212.Q )
  );
  al_dffl _11877_ (
    .clk(CK),
    .d(\DFF_1213.D ),
    .q(\DFF_1213.Q )
  );
  al_dffl _11878_ (
    .clk(CK),
    .d(\DFF_1214.D ),
    .q(\DFF_1214.Q )
  );
  al_dffl _11879_ (
    .clk(CK),
    .d(\DFF_1215.D ),
    .q(\DFF_1215.Q )
  );
  al_dffl _11880_ (
    .clk(CK),
    .d(\DFF_1216.D ),
    .q(\DFF_1216.Q )
  );
  al_dffl _11881_ (
    .clk(CK),
    .d(\DFF_1217.D ),
    .q(\DFF_1217.Q )
  );
  al_dffl _11882_ (
    .clk(CK),
    .d(\DFF_1218.D ),
    .q(\DFF_1218.Q )
  );
  al_dffl _11883_ (
    .clk(CK),
    .d(\DFF_1219.D ),
    .q(\DFF_1219.Q )
  );
  al_dffl _11884_ (
    .clk(CK),
    .d(\DFF_1220.D ),
    .q(\DFF_1220.Q )
  );
  al_dffl _11885_ (
    .clk(CK),
    .d(\DFF_1221.D ),
    .q(\DFF_1221.Q )
  );
  al_dffl _11886_ (
    .clk(CK),
    .d(\DFF_1222.D ),
    .q(\DFF_1222.Q )
  );
  al_dffl _11887_ (
    .clk(CK),
    .d(\DFF_1223.D ),
    .q(\DFF_1223.Q )
  );
  al_dffl _11888_ (
    .clk(CK),
    .d(\DFF_1224.D ),
    .q(\DFF_1224.Q )
  );
  al_dffl _11889_ (
    .clk(CK),
    .d(\DFF_1225.D ),
    .q(\DFF_1225.Q )
  );
  al_dffl _11890_ (
    .clk(CK),
    .d(\DFF_1226.D ),
    .q(\DFF_1226.Q )
  );
  al_dffl _11891_ (
    .clk(CK),
    .d(\DFF_1227.D ),
    .q(\DFF_1227.Q )
  );
  al_dffl _11892_ (
    .clk(CK),
    .d(\DFF_1228.D ),
    .q(\DFF_1228.Q )
  );
  al_dffl _11893_ (
    .clk(CK),
    .d(\DFF_1229.D ),
    .q(\DFF_1229.Q )
  );
  al_dffl _11894_ (
    .clk(CK),
    .d(\DFF_1230.D ),
    .q(\DFF_1230.Q )
  );
  al_dffl _11895_ (
    .clk(CK),
    .d(\DFF_1231.D ),
    .q(\DFF_1231.Q )
  );
  al_dffl _11896_ (
    .clk(CK),
    .d(\DFF_1232.D ),
    .q(\DFF_1232.Q )
  );
  al_dffl _11897_ (
    .clk(CK),
    .d(\DFF_1233.D ),
    .q(\DFF_1233.Q )
  );
  al_dffl _11898_ (
    .clk(CK),
    .d(\DFF_1234.D ),
    .q(\DFF_1234.Q )
  );
  al_dffl _11899_ (
    .clk(CK),
    .d(\DFF_1235.D ),
    .q(\DFF_1235.Q )
  );
  al_dffl _11900_ (
    .clk(CK),
    .d(\DFF_1236.D ),
    .q(\DFF_1236.Q )
  );
  al_dffl _11901_ (
    .clk(CK),
    .d(\DFF_1237.D ),
    .q(\DFF_1237.Q )
  );
  al_dffl _11902_ (
    .clk(CK),
    .d(\DFF_1238.D ),
    .q(\DFF_1238.Q )
  );
  al_dffl _11903_ (
    .clk(CK),
    .d(\DFF_1239.D ),
    .q(\DFF_1239.Q )
  );
  al_dffl _11904_ (
    .clk(CK),
    .d(\DFF_1240.D ),
    .q(\DFF_1240.Q )
  );
  al_dffl _11905_ (
    .clk(CK),
    .d(\DFF_1241.D ),
    .q(\DFF_1241.Q )
  );
  al_dffl _11906_ (
    .clk(CK),
    .d(\DFF_1242.D ),
    .q(\DFF_1242.Q )
  );
  al_dffl _11907_ (
    .clk(CK),
    .d(\DFF_1243.D ),
    .q(\DFF_1243.Q )
  );
  al_dffl _11908_ (
    .clk(CK),
    .d(\DFF_1244.D ),
    .q(\DFF_1244.Q )
  );
  al_dffl _11909_ (
    .clk(CK),
    .d(\DFF_1245.D ),
    .q(\DFF_1245.Q )
  );
  al_dffl _11910_ (
    .clk(CK),
    .d(\DFF_1246.D ),
    .q(\DFF_1246.Q )
  );
  al_dffl _11911_ (
    .clk(CK),
    .d(\DFF_1247.D ),
    .q(\DFF_1247.Q )
  );
  al_dffl _11912_ (
    .clk(CK),
    .d(\DFF_1248.D ),
    .q(\DFF_1248.Q )
  );
  al_dffl _11913_ (
    .clk(CK),
    .d(\DFF_1249.D ),
    .q(\DFF_1249.Q )
  );
  al_dffl _11914_ (
    .clk(CK),
    .d(\DFF_1250.D ),
    .q(\DFF_1250.Q )
  );
  al_dffl _11915_ (
    .clk(CK),
    .d(\DFF_1251.D ),
    .q(\DFF_1251.Q )
  );
  al_dffl _11916_ (
    .clk(CK),
    .d(\DFF_1252.D ),
    .q(\DFF_1252.Q )
  );
  al_dffl _11917_ (
    .clk(CK),
    .d(\DFF_1253.D ),
    .q(\DFF_1253.Q )
  );
  al_dffl _11918_ (
    .clk(CK),
    .d(\DFF_1254.D ),
    .q(\DFF_1254.Q )
  );
  al_dffl _11919_ (
    .clk(CK),
    .d(\DFF_1255.D ),
    .q(\DFF_1255.Q )
  );
  al_dffl _11920_ (
    .clk(CK),
    .d(\DFF_1256.D ),
    .q(\DFF_1256.Q )
  );
  al_dffl _11921_ (
    .clk(CK),
    .d(\DFF_1257.D ),
    .q(\DFF_1257.Q )
  );
  al_dffl _11922_ (
    .clk(CK),
    .d(\DFF_1258.D ),
    .q(\DFF_1258.Q )
  );
  al_dffl _11923_ (
    .clk(CK),
    .d(\DFF_1259.D ),
    .q(\DFF_1259.Q )
  );
  al_dffl _11924_ (
    .clk(CK),
    .d(\DFF_1260.D ),
    .q(\DFF_1260.Q )
  );
  al_dffl _11925_ (
    .clk(CK),
    .d(\DFF_1261.D ),
    .q(\DFF_1261.Q )
  );
  al_dffl _11926_ (
    .clk(CK),
    .d(\DFF_1262.D ),
    .q(\DFF_1262.Q )
  );
  al_dffl _11927_ (
    .clk(CK),
    .d(\DFF_1263.D ),
    .q(\DFF_1263.Q )
  );
  al_dffl _11928_ (
    .clk(CK),
    .d(\DFF_1264.D ),
    .q(\DFF_1264.Q )
  );
  al_dffl _11929_ (
    .clk(CK),
    .d(\DFF_1265.D ),
    .q(\DFF_1265.Q )
  );
  al_dffl _11930_ (
    .clk(CK),
    .d(\DFF_1266.D ),
    .q(\DFF_1266.Q )
  );
  al_dffl _11931_ (
    .clk(CK),
    .d(\DFF_1267.D ),
    .q(\DFF_1267.Q )
  );
  al_dffl _11932_ (
    .clk(CK),
    .d(\DFF_1268.D ),
    .q(\DFF_1268.Q )
  );
  al_dffl _11933_ (
    .clk(CK),
    .d(\DFF_1269.D ),
    .q(\DFF_1269.Q )
  );
  al_dffl _11934_ (
    .clk(CK),
    .d(\DFF_1270.D ),
    .q(\DFF_1270.Q )
  );
  al_dffl _11935_ (
    .clk(CK),
    .d(\DFF_1271.D ),
    .q(\DFF_1271.Q )
  );
  al_dffl _11936_ (
    .clk(CK),
    .d(\DFF_1272.D ),
    .q(\DFF_1272.Q )
  );
  al_dffl _11937_ (
    .clk(CK),
    .d(\DFF_1273.D ),
    .q(\DFF_1273.Q )
  );
  al_dffl _11938_ (
    .clk(CK),
    .d(\DFF_1274.D ),
    .q(\DFF_1274.Q )
  );
  al_dffl _11939_ (
    .clk(CK),
    .d(\DFF_1275.D ),
    .q(\DFF_1275.Q )
  );
  al_dffl _11940_ (
    .clk(CK),
    .d(\DFF_1276.D ),
    .q(\DFF_1276.Q )
  );
  al_dffl _11941_ (
    .clk(CK),
    .d(\DFF_1277.D ),
    .q(\DFF_1277.Q )
  );
  al_dffl _11942_ (
    .clk(CK),
    .d(\DFF_1278.D ),
    .q(\DFF_1278.Q )
  );
  al_dffl _11943_ (
    .clk(CK),
    .d(\DFF_1279.D ),
    .q(\DFF_1279.Q )
  );
  al_dffl _11944_ (
    .clk(CK),
    .d(\DFF_1280.D ),
    .q(\DFF_1280.Q )
  );
  al_dffl _11945_ (
    .clk(CK),
    .d(\DFF_1281.D ),
    .q(\DFF_1281.Q )
  );
  al_dffl _11946_ (
    .clk(CK),
    .d(\DFF_1282.D ),
    .q(\DFF_1282.Q )
  );
  al_dffl _11947_ (
    .clk(CK),
    .d(\DFF_1283.D ),
    .q(\DFF_1283.Q )
  );
  al_dffl _11948_ (
    .clk(CK),
    .d(\DFF_1284.D ),
    .q(\DFF_1284.Q )
  );
  al_dffl _11949_ (
    .clk(CK),
    .d(\DFF_1285.D ),
    .q(\DFF_1285.Q )
  );
  al_dffl _11950_ (
    .clk(CK),
    .d(\DFF_1286.D ),
    .q(\DFF_1286.Q )
  );
  al_dffl _11951_ (
    .clk(CK),
    .d(\DFF_1287.D ),
    .q(\DFF_1287.Q )
  );
  al_dffl _11952_ (
    .clk(CK),
    .d(\DFF_1288.D ),
    .q(\DFF_1288.Q )
  );
  al_dffl _11953_ (
    .clk(CK),
    .d(\DFF_1289.D ),
    .q(\DFF_1289.Q )
  );
  al_dffl _11954_ (
    .clk(CK),
    .d(\DFF_1290.D ),
    .q(\DFF_1290.Q )
  );
  al_dffl _11955_ (
    .clk(CK),
    .d(\DFF_1291.D ),
    .q(\DFF_1291.Q )
  );
  al_dffl _11956_ (
    .clk(CK),
    .d(\DFF_1292.D ),
    .q(\DFF_1292.Q )
  );
  al_dffl _11957_ (
    .clk(CK),
    .d(\DFF_1293.D ),
    .q(\DFF_1293.Q )
  );
  al_dffl _11958_ (
    .clk(CK),
    .d(\DFF_1294.D ),
    .q(\DFF_1294.Q )
  );
  al_dffl _11959_ (
    .clk(CK),
    .d(\DFF_1295.D ),
    .q(\DFF_1295.Q )
  );
  al_dffl _11960_ (
    .clk(CK),
    .d(\DFF_1296.D ),
    .q(\DFF_1296.Q )
  );
  al_dffl _11961_ (
    .clk(CK),
    .d(\DFF_1297.D ),
    .q(\DFF_1297.Q )
  );
  al_dffl _11962_ (
    .clk(CK),
    .d(\DFF_1298.D ),
    .q(\DFF_1298.Q )
  );
  al_dffl _11963_ (
    .clk(CK),
    .d(\DFF_1299.D ),
    .q(\DFF_1299.Q )
  );
  al_dffl _11964_ (
    .clk(CK),
    .d(\DFF_1300.D ),
    .q(\DFF_1300.Q )
  );
  al_dffl _11965_ (
    .clk(CK),
    .d(\DFF_1301.D ),
    .q(\DFF_1301.Q )
  );
  al_dffl _11966_ (
    .clk(CK),
    .d(\DFF_1302.D ),
    .q(\DFF_1302.Q )
  );
  al_dffl _11967_ (
    .clk(CK),
    .d(\DFF_1303.D ),
    .q(\DFF_1303.Q )
  );
  al_dffl _11968_ (
    .clk(CK),
    .d(\DFF_1304.D ),
    .q(\DFF_1304.Q )
  );
  al_dffl _11969_ (
    .clk(CK),
    .d(\DFF_1305.D ),
    .q(\DFF_1305.Q )
  );
  al_dffl _11970_ (
    .clk(CK),
    .d(\DFF_1306.D ),
    .q(\DFF_1306.Q )
  );
  al_dffl _11971_ (
    .clk(CK),
    .d(\DFF_1307.D ),
    .q(\DFF_1307.Q )
  );
  al_dffl _11972_ (
    .clk(CK),
    .d(\DFF_1308.D ),
    .q(\DFF_1308.Q )
  );
  al_dffl _11973_ (
    .clk(CK),
    .d(\DFF_1309.D ),
    .q(\DFF_1309.Q )
  );
  al_dffl _11974_ (
    .clk(CK),
    .d(\DFF_1310.D ),
    .q(\DFF_1310.Q )
  );
  al_dffl _11975_ (
    .clk(CK),
    .d(\DFF_1311.D ),
    .q(\DFF_1311.Q )
  );
  al_dffl _11976_ (
    .clk(CK),
    .d(\DFF_1312.D ),
    .q(\DFF_1312.Q )
  );
  al_dffl _11977_ (
    .clk(CK),
    .d(\DFF_1313.D ),
    .q(\DFF_1313.Q )
  );
  al_dffl _11978_ (
    .clk(CK),
    .d(\DFF_1314.D ),
    .q(\DFF_1314.Q )
  );
  al_dffl _11979_ (
    .clk(CK),
    .d(\DFF_1315.D ),
    .q(\DFF_1315.Q )
  );
  al_dffl _11980_ (
    .clk(CK),
    .d(\DFF_1316.D ),
    .q(\DFF_1316.Q )
  );
  al_dffl _11981_ (
    .clk(CK),
    .d(\DFF_1317.D ),
    .q(\DFF_1317.Q )
  );
  al_dffl _11982_ (
    .clk(CK),
    .d(\DFF_1318.D ),
    .q(\DFF_1318.Q )
  );
  al_dffl _11983_ (
    .clk(CK),
    .d(\DFF_1319.D ),
    .q(\DFF_1319.Q )
  );
  al_dffl _11984_ (
    .clk(CK),
    .d(\DFF_1320.D ),
    .q(\DFF_1320.Q )
  );
  al_dffl _11985_ (
    .clk(CK),
    .d(\DFF_1321.D ),
    .q(\DFF_1321.Q )
  );
  al_dffl _11986_ (
    .clk(CK),
    .d(\DFF_1322.D ),
    .q(\DFF_1322.Q )
  );
  al_dffl _11987_ (
    .clk(CK),
    .d(\DFF_1323.D ),
    .q(\DFF_1323.Q )
  );
  al_dffl _11988_ (
    .clk(CK),
    .d(\DFF_1324.D ),
    .q(\DFF_1324.Q )
  );
  al_dffl _11989_ (
    .clk(CK),
    .d(\DFF_1325.D ),
    .q(\DFF_1325.Q )
  );
  al_dffl _11990_ (
    .clk(CK),
    .d(\DFF_1326.D ),
    .q(\DFF_1326.Q )
  );
  al_dffl _11991_ (
    .clk(CK),
    .d(\DFF_1327.D ),
    .q(\DFF_1327.Q )
  );
  al_dffl _11992_ (
    .clk(CK),
    .d(\DFF_1328.D ),
    .q(\DFF_1328.Q )
  );
  al_dffl _11993_ (
    .clk(CK),
    .d(\DFF_1329.D ),
    .q(\DFF_1329.Q )
  );
  al_dffl _11994_ (
    .clk(CK),
    .d(\DFF_1330.D ),
    .q(\DFF_1330.Q )
  );
  al_dffl _11995_ (
    .clk(CK),
    .d(\DFF_1331.D ),
    .q(\DFF_1331.Q )
  );
  al_dffl _11996_ (
    .clk(CK),
    .d(\DFF_1332.D ),
    .q(\DFF_1332.Q )
  );
  al_dffl _11997_ (
    .clk(CK),
    .d(\DFF_1333.D ),
    .q(\DFF_1333.Q )
  );
  al_dffl _11998_ (
    .clk(CK),
    .d(\DFF_1334.D ),
    .q(\DFF_1334.Q )
  );
  al_dffl _11999_ (
    .clk(CK),
    .d(\DFF_1335.D ),
    .q(\DFF_1335.Q )
  );
  al_dffl _12000_ (
    .clk(CK),
    .d(\DFF_1336.D ),
    .q(\DFF_1336.Q )
  );
  al_dffl _12001_ (
    .clk(CK),
    .d(\DFF_1337.D ),
    .q(\DFF_1337.Q )
  );
  al_dffl _12002_ (
    .clk(CK),
    .d(\DFF_1338.D ),
    .q(\DFF_1338.Q )
  );
  al_dffl _12003_ (
    .clk(CK),
    .d(\DFF_1339.D ),
    .q(\DFF_1339.Q )
  );
  al_dffl _12004_ (
    .clk(CK),
    .d(\DFF_1340.D ),
    .q(\DFF_1340.Q )
  );
  al_dffl _12005_ (
    .clk(CK),
    .d(\DFF_1341.D ),
    .q(\DFF_1341.Q )
  );
  al_dffl _12006_ (
    .clk(CK),
    .d(\DFF_1342.D ),
    .q(\DFF_1342.Q )
  );
  al_dffl _12007_ (
    .clk(CK),
    .d(\DFF_1343.D ),
    .q(\DFF_1343.Q )
  );
  al_dffl _12008_ (
    .clk(CK),
    .d(\DFF_1344.D ),
    .q(\DFF_1344.Q )
  );
  al_dffl _12009_ (
    .clk(CK),
    .d(\DFF_1345.D ),
    .q(\DFF_1345.Q )
  );
  al_dffl _12010_ (
    .clk(CK),
    .d(\DFF_1346.D ),
    .q(\DFF_1346.Q )
  );
  al_dffl _12011_ (
    .clk(CK),
    .d(\DFF_1347.D ),
    .q(\DFF_1347.Q )
  );
  al_dffl _12012_ (
    .clk(CK),
    .d(\DFF_1348.D ),
    .q(\DFF_1348.Q )
  );
  al_dffl _12013_ (
    .clk(CK),
    .d(\DFF_1349.D ),
    .q(\DFF_1349.Q )
  );
  al_dffl _12014_ (
    .clk(CK),
    .d(\DFF_1350.D ),
    .q(\DFF_1350.Q )
  );
  al_dffl _12015_ (
    .clk(CK),
    .d(\DFF_1351.D ),
    .q(\DFF_1351.Q )
  );
  al_dffl _12016_ (
    .clk(CK),
    .d(\DFF_1352.D ),
    .q(\DFF_1352.Q )
  );
  al_dffl _12017_ (
    .clk(CK),
    .d(\DFF_1353.D ),
    .q(\DFF_1353.Q )
  );
  al_dffl _12018_ (
    .clk(CK),
    .d(\DFF_1354.D ),
    .q(\DFF_1354.Q )
  );
  al_dffl _12019_ (
    .clk(CK),
    .d(\DFF_1355.D ),
    .q(\DFF_1355.Q )
  );
  al_dffl _12020_ (
    .clk(CK),
    .d(\DFF_1356.D ),
    .q(\DFF_1356.Q )
  );
  al_dffl _12021_ (
    .clk(CK),
    .d(\DFF_1357.D ),
    .q(\DFF_1357.Q )
  );
  al_dffl _12022_ (
    .clk(CK),
    .d(\DFF_1358.D ),
    .q(\DFF_1358.Q )
  );
  al_dffl _12023_ (
    .clk(CK),
    .d(\DFF_1359.D ),
    .q(\DFF_1359.Q )
  );
  al_dffl _12024_ (
    .clk(CK),
    .d(\DFF_1360.D ),
    .q(\DFF_1360.Q )
  );
  al_dffl _12025_ (
    .clk(CK),
    .d(\DFF_1361.D ),
    .q(\DFF_1361.Q )
  );
  al_dffl _12026_ (
    .clk(CK),
    .d(\DFF_1362.D ),
    .q(\DFF_1362.Q )
  );
  al_dffl _12027_ (
    .clk(CK),
    .d(\DFF_1363.D ),
    .q(\DFF_1363.Q )
  );
  al_dffl _12028_ (
    .clk(CK),
    .d(\DFF_1364.D ),
    .q(\DFF_1364.Q )
  );
  al_dffl _12029_ (
    .clk(CK),
    .d(\DFF_1365.D ),
    .q(\DFF_1365.Q )
  );
  al_dffl _12030_ (
    .clk(CK),
    .d(\DFF_1366.D ),
    .q(\DFF_1366.Q )
  );
  al_dffl _12031_ (
    .clk(CK),
    .d(\DFF_1367.D ),
    .q(\DFF_1367.Q )
  );
  al_dffl _12032_ (
    .clk(CK),
    .d(\DFF_1368.D ),
    .q(\DFF_1368.Q )
  );
  al_dffl _12033_ (
    .clk(CK),
    .d(\DFF_1369.D ),
    .q(\DFF_1369.Q )
  );
  al_dffl _12034_ (
    .clk(CK),
    .d(\DFF_1370.D ),
    .q(\DFF_1370.Q )
  );
  al_dffl _12035_ (
    .clk(CK),
    .d(\DFF_1371.D ),
    .q(\DFF_1371.Q )
  );
  al_dffl _12036_ (
    .clk(CK),
    .d(\DFF_1372.D ),
    .q(\DFF_1372.Q )
  );
  al_dffl _12037_ (
    .clk(CK),
    .d(\DFF_1373.D ),
    .q(\DFF_1373.Q )
  );
  al_dffl _12038_ (
    .clk(CK),
    .d(\DFF_1374.D ),
    .q(\DFF_1374.Q )
  );
  al_dffl _12039_ (
    .clk(CK),
    .d(\DFF_1375.D ),
    .q(\DFF_1375.Q )
  );
  al_dffl _12040_ (
    .clk(CK),
    .d(\DFF_1376.D ),
    .q(\DFF_1376.Q )
  );
  al_dffl _12041_ (
    .clk(CK),
    .d(\DFF_1377.D ),
    .q(\DFF_1377.Q )
  );
  al_dffl _12042_ (
    .clk(CK),
    .d(\DFF_1378.D ),
    .q(\DFF_1378.Q )
  );
  al_dffl _12043_ (
    .clk(CK),
    .d(\DFF_1379.D ),
    .q(\DFF_1379.Q )
  );
  al_dffl _12044_ (
    .clk(CK),
    .d(\DFF_1380.D ),
    .q(\DFF_1380.Q )
  );
  al_dffl _12045_ (
    .clk(CK),
    .d(\DFF_1381.D ),
    .q(\DFF_1381.Q )
  );
  al_dffl _12046_ (
    .clk(CK),
    .d(\DFF_1382.D ),
    .q(\DFF_1382.Q )
  );
  al_dffl _12047_ (
    .clk(CK),
    .d(\DFF_1383.D ),
    .q(\DFF_1383.Q )
  );
  al_dffl _12048_ (
    .clk(CK),
    .d(\DFF_1384.D ),
    .q(\DFF_1384.Q )
  );
  al_dffl _12049_ (
    .clk(CK),
    .d(\DFF_1385.D ),
    .q(\DFF_1385.Q )
  );
  al_dffl _12050_ (
    .clk(CK),
    .d(\DFF_1386.D ),
    .q(\DFF_1386.Q )
  );
  al_dffl _12051_ (
    .clk(CK),
    .d(\DFF_1387.D ),
    .q(\DFF_1387.Q )
  );
  al_dffl _12052_ (
    .clk(CK),
    .d(\DFF_1388.D ),
    .q(\DFF_1388.Q )
  );
  al_dffl _12053_ (
    .clk(CK),
    .d(\DFF_1389.D ),
    .q(\DFF_1389.Q )
  );
  al_dffl _12054_ (
    .clk(CK),
    .d(\DFF_1390.D ),
    .q(\DFF_1390.Q )
  );
  al_dffl _12055_ (
    .clk(CK),
    .d(\DFF_1391.D ),
    .q(\DFF_1391.Q )
  );
  al_dffl _12056_ (
    .clk(CK),
    .d(\DFF_1392.D ),
    .q(\DFF_1392.Q )
  );
  al_dffl _12057_ (
    .clk(CK),
    .d(\DFF_1393.D ),
    .q(\DFF_1393.Q )
  );
  al_dffl _12058_ (
    .clk(CK),
    .d(\DFF_1394.D ),
    .q(\DFF_1394.Q )
  );
  al_dffl _12059_ (
    .clk(CK),
    .d(\DFF_1395.D ),
    .q(\DFF_1395.Q )
  );
  al_dffl _12060_ (
    .clk(CK),
    .d(\DFF_1396.D ),
    .q(\DFF_1396.Q )
  );
  al_dffl _12061_ (
    .clk(CK),
    .d(\DFF_1397.D ),
    .q(\DFF_1397.Q )
  );
  al_dffl _12062_ (
    .clk(CK),
    .d(\DFF_1398.D ),
    .q(\DFF_1398.Q )
  );
  al_dffl _12063_ (
    .clk(CK),
    .d(\DFF_1399.D ),
    .q(\DFF_1399.Q )
  );
  al_dffl _12064_ (
    .clk(CK),
    .d(\DFF_1400.D ),
    .q(\DFF_1400.Q )
  );
  al_dffl _12065_ (
    .clk(CK),
    .d(\DFF_1401.D ),
    .q(\DFF_1401.Q )
  );
  al_dffl _12066_ (
    .clk(CK),
    .d(\DFF_1402.D ),
    .q(\DFF_1402.Q )
  );
  al_dffl _12067_ (
    .clk(CK),
    .d(\DFF_1403.D ),
    .q(\DFF_1403.Q )
  );
  al_dffl _12068_ (
    .clk(CK),
    .d(\DFF_1404.D ),
    .q(\DFF_1404.Q )
  );
  al_dffl _12069_ (
    .clk(CK),
    .d(\DFF_1405.D ),
    .q(\DFF_1405.Q )
  );
  al_dffl _12070_ (
    .clk(CK),
    .d(\DFF_1406.D ),
    .q(\DFF_1406.Q )
  );
  al_dffl _12071_ (
    .clk(CK),
    .d(\DFF_1407.D ),
    .q(\DFF_1407.Q )
  );
  al_dffl _12072_ (
    .clk(CK),
    .d(\DFF_1408.D ),
    .q(\DFF_1408.Q )
  );
  al_dffl _12073_ (
    .clk(CK),
    .d(\DFF_1409.D ),
    .q(\DFF_1409.Q )
  );
  al_dffl _12074_ (
    .clk(CK),
    .d(\DFF_1410.D ),
    .q(\DFF_1410.Q )
  );
  al_dffl _12075_ (
    .clk(CK),
    .d(\DFF_1411.D ),
    .q(\DFF_1411.Q )
  );
  al_dffl _12076_ (
    .clk(CK),
    .d(\DFF_1412.D ),
    .q(\DFF_1412.Q )
  );
  al_dffl _12077_ (
    .clk(CK),
    .d(\DFF_1413.D ),
    .q(\DFF_1413.Q )
  );
  al_dffl _12078_ (
    .clk(CK),
    .d(\DFF_1414.D ),
    .q(\DFF_1414.Q )
  );
  al_dffl _12079_ (
    .clk(CK),
    .d(\DFF_1415.D ),
    .q(\DFF_1415.Q )
  );
  al_dffl _12080_ (
    .clk(CK),
    .d(\DFF_1416.D ),
    .q(\DFF_1416.Q )
  );
  al_dffl _12081_ (
    .clk(CK),
    .d(\DFF_1417.D ),
    .q(\DFF_1417.Q )
  );
  al_dffl _12082_ (
    .clk(CK),
    .d(\DFF_1418.D ),
    .q(\DFF_1418.Q )
  );
  al_dffl _12083_ (
    .clk(CK),
    .d(\DFF_1419.D ),
    .q(\DFF_1419.Q )
  );
  al_dffl _12084_ (
    .clk(CK),
    .d(\DFF_1420.D ),
    .q(\DFF_1420.Q )
  );
  al_dffl _12085_ (
    .clk(CK),
    .d(\DFF_1421.D ),
    .q(\DFF_1421.Q )
  );
  al_dffl _12086_ (
    .clk(CK),
    .d(\DFF_1422.D ),
    .q(\DFF_1422.Q )
  );
  al_dffl _12087_ (
    .clk(CK),
    .d(\DFF_1423.D ),
    .q(\DFF_1423.Q )
  );
  al_dffl _12088_ (
    .clk(CK),
    .d(\DFF_1424.D ),
    .q(\DFF_1424.Q )
  );
  al_dffl _12089_ (
    .clk(CK),
    .d(\DFF_1425.D ),
    .q(\DFF_1425.Q )
  );
  al_dffl _12090_ (
    .clk(CK),
    .d(\DFF_1426.D ),
    .q(\DFF_1426.Q )
  );
  al_dffl _12091_ (
    .clk(CK),
    .d(\DFF_1427.D ),
    .q(\DFF_1427.Q )
  );
  al_dffl _12092_ (
    .clk(CK),
    .d(\DFF_1428.D ),
    .q(\DFF_1428.Q )
  );
  al_dffl _12093_ (
    .clk(CK),
    .d(\DFF_1429.D ),
    .q(\DFF_1429.Q )
  );
  al_dffl _12094_ (
    .clk(CK),
    .d(\DFF_1430.D ),
    .q(\DFF_1430.Q )
  );
  al_dffl _12095_ (
    .clk(CK),
    .d(\DFF_1431.D ),
    .q(\DFF_1431.Q )
  );
  al_dffl _12096_ (
    .clk(CK),
    .d(\DFF_1432.D ),
    .q(\DFF_1432.Q )
  );
  al_dffl _12097_ (
    .clk(CK),
    .d(\DFF_1433.D ),
    .q(\DFF_1433.Q )
  );
  al_dffl _12098_ (
    .clk(CK),
    .d(\DFF_1434.D ),
    .q(\DFF_1434.Q )
  );
  al_dffl _12099_ (
    .clk(CK),
    .d(\DFF_1435.D ),
    .q(\DFF_1435.Q )
  );
  al_dffl _12100_ (
    .clk(CK),
    .d(\DFF_1436.D ),
    .q(\DFF_1436.Q )
  );
  al_dffl _12101_ (
    .clk(CK),
    .d(\DFF_1437.D ),
    .q(\DFF_1437.Q )
  );
  al_dffl _12102_ (
    .clk(CK),
    .d(\DFF_1438.D ),
    .q(\DFF_1438.Q )
  );
  al_dffl _12103_ (
    .clk(CK),
    .d(\DFF_1439.D ),
    .q(\DFF_1439.Q )
  );
  al_dffl _12104_ (
    .clk(CK),
    .d(\DFF_1440.D ),
    .q(\DFF_1440.Q )
  );
  al_dffl _12105_ (
    .clk(CK),
    .d(\DFF_1441.D ),
    .q(\DFF_1441.Q )
  );
  al_dffl _12106_ (
    .clk(CK),
    .d(\DFF_1442.D ),
    .q(\DFF_1442.Q )
  );
  al_dffl _12107_ (
    .clk(CK),
    .d(\DFF_1443.D ),
    .q(\DFF_1443.Q )
  );
  al_dffl _12108_ (
    .clk(CK),
    .d(\DFF_1444.D ),
    .q(\DFF_1444.Q )
  );
  al_dffl _12109_ (
    .clk(CK),
    .d(\DFF_1445.D ),
    .q(\DFF_1445.Q )
  );
  al_dffl _12110_ (
    .clk(CK),
    .d(\DFF_1446.D ),
    .q(\DFF_1446.Q )
  );
  al_dffl _12111_ (
    .clk(CK),
    .d(\DFF_1447.D ),
    .q(\DFF_1447.Q )
  );
  al_dffl _12112_ (
    .clk(CK),
    .d(\DFF_1448.D ),
    .q(\DFF_1448.Q )
  );
  al_dffl _12113_ (
    .clk(CK),
    .d(\DFF_1449.D ),
    .q(\DFF_1449.Q )
  );
  al_dffl _12114_ (
    .clk(CK),
    .d(\DFF_1450.D ),
    .q(\DFF_1450.Q )
  );
  al_dffl _12115_ (
    .clk(CK),
    .d(\DFF_1451.D ),
    .q(\DFF_1451.Q )
  );
  al_dffl _12116_ (
    .clk(CK),
    .d(\DFF_1452.D ),
    .q(\DFF_1452.Q )
  );
  al_dffl _12117_ (
    .clk(CK),
    .d(\DFF_1453.D ),
    .q(\DFF_1453.Q )
  );
  al_dffl _12118_ (
    .clk(CK),
    .d(\DFF_1454.D ),
    .q(\DFF_1454.Q )
  );
  al_dffl _12119_ (
    .clk(CK),
    .d(\DFF_1455.D ),
    .q(\DFF_1455.Q )
  );
  al_dffl _12120_ (
    .clk(CK),
    .d(\DFF_1456.D ),
    .q(\DFF_1456.Q )
  );
  al_dffl _12121_ (
    .clk(CK),
    .d(\DFF_1457.D ),
    .q(\DFF_1457.Q )
  );
  al_dffl _12122_ (
    .clk(CK),
    .d(\DFF_1458.D ),
    .q(\DFF_1458.Q )
  );
  al_dffl _12123_ (
    .clk(CK),
    .d(\DFF_1459.D ),
    .q(\DFF_1459.Q )
  );
  al_dffl _12124_ (
    .clk(CK),
    .d(\DFF_1460.D ),
    .q(\DFF_1460.Q )
  );
  al_dffl _12125_ (
    .clk(CK),
    .d(\DFF_1461.D ),
    .q(\DFF_1461.Q )
  );
  al_dffl _12126_ (
    .clk(CK),
    .d(\DFF_1462.D ),
    .q(\DFF_1462.Q )
  );
  al_dffl _12127_ (
    .clk(CK),
    .d(\DFF_1463.D ),
    .q(\DFF_1463.Q )
  );
  al_dffl _12128_ (
    .clk(CK),
    .d(\DFF_1464.D ),
    .q(\DFF_1464.Q )
  );
  al_dffl _12129_ (
    .clk(CK),
    .d(\DFF_1465.D ),
    .q(\DFF_1465.Q )
  );
  al_dffl _12130_ (
    .clk(CK),
    .d(\DFF_1466.D ),
    .q(\DFF_1466.Q )
  );
  al_dffl _12131_ (
    .clk(CK),
    .d(\DFF_1467.D ),
    .q(\DFF_1467.Q )
  );
  al_dffl _12132_ (
    .clk(CK),
    .d(\DFF_1468.D ),
    .q(\DFF_1468.Q )
  );
  al_dffl _12133_ (
    .clk(CK),
    .d(\DFF_1469.D ),
    .q(\DFF_1469.Q )
  );
  al_dffl _12134_ (
    .clk(CK),
    .d(\DFF_1470.D ),
    .q(\DFF_1470.Q )
  );
  al_dffl _12135_ (
    .clk(CK),
    .d(\DFF_1471.D ),
    .q(\DFF_1471.Q )
  );
  al_dffl _12136_ (
    .clk(CK),
    .d(\DFF_1472.D ),
    .q(\DFF_1472.Q )
  );
  al_dffl _12137_ (
    .clk(CK),
    .d(\DFF_1473.D ),
    .q(\DFF_1473.Q )
  );
  al_dffl _12138_ (
    .clk(CK),
    .d(\DFF_1474.D ),
    .q(\DFF_1474.Q )
  );
  al_dffl _12139_ (
    .clk(CK),
    .d(\DFF_1475.D ),
    .q(\DFF_1475.Q )
  );
  al_dffl _12140_ (
    .clk(CK),
    .d(\DFF_1476.D ),
    .q(\DFF_1476.Q )
  );
  al_dffl _12141_ (
    .clk(CK),
    .d(\DFF_1477.D ),
    .q(\DFF_1477.Q )
  );
  al_dffl _12142_ (
    .clk(CK),
    .d(\DFF_1478.D ),
    .q(\DFF_1478.Q )
  );
  al_dffl _12143_ (
    .clk(CK),
    .d(\DFF_1479.D ),
    .q(\DFF_1479.Q )
  );
  al_dffl _12144_ (
    .clk(CK),
    .d(\DFF_1480.D ),
    .q(\DFF_1480.Q )
  );
  al_dffl _12145_ (
    .clk(CK),
    .d(\DFF_1481.D ),
    .q(\DFF_1481.Q )
  );
  al_dffl _12146_ (
    .clk(CK),
    .d(\DFF_1482.D ),
    .q(\DFF_1482.Q )
  );
  al_dffl _12147_ (
    .clk(CK),
    .d(\DFF_1483.D ),
    .q(\DFF_1483.Q )
  );
  al_dffl _12148_ (
    .clk(CK),
    .d(\DFF_1484.D ),
    .q(\DFF_1484.Q )
  );
  al_dffl _12149_ (
    .clk(CK),
    .d(\DFF_1485.D ),
    .q(\DFF_1485.Q )
  );
  al_dffl _12150_ (
    .clk(CK),
    .d(\DFF_1486.D ),
    .q(\DFF_1486.Q )
  );
  al_dffl _12151_ (
    .clk(CK),
    .d(\DFF_1487.D ),
    .q(\DFF_1487.Q )
  );
  al_dffl _12152_ (
    .clk(CK),
    .d(\DFF_1488.D ),
    .q(\DFF_1488.Q )
  );
  al_dffl _12153_ (
    .clk(CK),
    .d(\DFF_1489.D ),
    .q(\DFF_1489.Q )
  );
  al_dffl _12154_ (
    .clk(CK),
    .d(\DFF_1490.D ),
    .q(\DFF_1490.Q )
  );
  al_dffl _12155_ (
    .clk(CK),
    .d(\DFF_1491.D ),
    .q(\DFF_1491.Q )
  );
  al_dffl _12156_ (
    .clk(CK),
    .d(\DFF_1492.D ),
    .q(\DFF_1492.Q )
  );
  al_dffl _12157_ (
    .clk(CK),
    .d(\DFF_1493.D ),
    .q(\DFF_1493.Q )
  );
  al_dffl _12158_ (
    .clk(CK),
    .d(\DFF_1494.D ),
    .q(\DFF_1494.Q )
  );
  al_dffl _12159_ (
    .clk(CK),
    .d(\DFF_1495.D ),
    .q(\DFF_1495.Q )
  );
  al_dffl _12160_ (
    .clk(CK),
    .d(\DFF_1496.D ),
    .q(\DFF_1496.Q )
  );
  al_dffl _12161_ (
    .clk(CK),
    .d(\DFF_1497.D ),
    .q(\DFF_1497.Q )
  );
  al_dffl _12162_ (
    .clk(CK),
    .d(\DFF_1498.D ),
    .q(\DFF_1498.Q )
  );
  al_dffl _12163_ (
    .clk(CK),
    .d(\DFF_1499.D ),
    .q(\DFF_1499.Q )
  );
  al_dffl _12164_ (
    .clk(CK),
    .d(\DFF_1500.D ),
    .q(\DFF_1500.Q )
  );
  al_dffl _12165_ (
    .clk(CK),
    .d(\DFF_1501.D ),
    .q(\DFF_1501.Q )
  );
  al_dffl _12166_ (
    .clk(CK),
    .d(\DFF_1502.D ),
    .q(\DFF_1502.Q )
  );
  al_dffl _12167_ (
    .clk(CK),
    .d(\DFF_1503.D ),
    .q(\DFF_1503.Q )
  );
  al_dffl _12168_ (
    .clk(CK),
    .d(\DFF_1504.D ),
    .q(\DFF_1504.Q )
  );
  al_dffl _12169_ (
    .clk(CK),
    .d(\DFF_1505.D ),
    .q(\DFF_1505.Q )
  );
  al_dffl _12170_ (
    .clk(CK),
    .d(\DFF_1506.D ),
    .q(\DFF_1506.Q )
  );
  al_dffl _12171_ (
    .clk(CK),
    .d(\DFF_1507.D ),
    .q(\DFF_1507.Q )
  );
  al_dffl _12172_ (
    .clk(CK),
    .d(\DFF_1508.D ),
    .q(\DFF_1508.Q )
  );
  al_dffl _12173_ (
    .clk(CK),
    .d(\DFF_1509.D ),
    .q(\DFF_1509.Q )
  );
  al_dffl _12174_ (
    .clk(CK),
    .d(\DFF_1510.D ),
    .q(\DFF_1510.Q )
  );
  al_dffl _12175_ (
    .clk(CK),
    .d(\DFF_1511.D ),
    .q(\DFF_1511.Q )
  );
  al_dffl _12176_ (
    .clk(CK),
    .d(\DFF_1512.D ),
    .q(\DFF_1512.Q )
  );
  al_dffl _12177_ (
    .clk(CK),
    .d(\DFF_1513.D ),
    .q(\DFF_1513.Q )
  );
  al_dffl _12178_ (
    .clk(CK),
    .d(\DFF_1514.D ),
    .q(\DFF_1514.Q )
  );
  al_dffl _12179_ (
    .clk(CK),
    .d(\DFF_1515.D ),
    .q(\DFF_1515.Q )
  );
  al_dffl _12180_ (
    .clk(CK),
    .d(\DFF_1516.D ),
    .q(\DFF_1516.Q )
  );
  al_dffl _12181_ (
    .clk(CK),
    .d(\DFF_1517.D ),
    .q(\DFF_1517.Q )
  );
  al_dffl _12182_ (
    .clk(CK),
    .d(\DFF_1518.D ),
    .q(\DFF_1518.Q )
  );
  al_dffl _12183_ (
    .clk(CK),
    .d(\DFF_1519.D ),
    .q(\DFF_1519.Q )
  );
  al_dffl _12184_ (
    .clk(CK),
    .d(\DFF_1520.D ),
    .q(\DFF_1520.Q )
  );
  al_dffl _12185_ (
    .clk(CK),
    .d(\DFF_1521.D ),
    .q(\DFF_1521.Q )
  );
  al_dffl _12186_ (
    .clk(CK),
    .d(\DFF_1522.D ),
    .q(\DFF_1522.Q )
  );
  al_dffl _12187_ (
    .clk(CK),
    .d(\DFF_1523.D ),
    .q(\DFF_1523.Q )
  );
  al_dffl _12188_ (
    .clk(CK),
    .d(\DFF_1524.D ),
    .q(\DFF_1524.Q )
  );
  al_dffl _12189_ (
    .clk(CK),
    .d(\DFF_1525.D ),
    .q(\DFF_1525.Q )
  );
  al_dffl _12190_ (
    .clk(CK),
    .d(\DFF_1526.D ),
    .q(\DFF_1526.Q )
  );
  al_dffl _12191_ (
    .clk(CK),
    .d(\DFF_1527.D ),
    .q(\DFF_1527.Q )
  );
  al_dffl _12192_ (
    .clk(CK),
    .d(\DFF_1528.D ),
    .q(\DFF_1528.Q )
  );
  al_dffl _12193_ (
    .clk(CK),
    .d(\DFF_1529.D ),
    .q(\DFF_1529.Q )
  );
  al_dffl _12194_ (
    .clk(CK),
    .d(\DFF_1530.D ),
    .q(\DFF_1530.Q )
  );
  al_dffl _12195_ (
    .clk(CK),
    .d(\DFF_1531.D ),
    .q(\DFF_1531.Q )
  );
  al_dffl _12196_ (
    .clk(CK),
    .d(\DFF_1532.D ),
    .q(\DFF_1532.Q )
  );
  al_dffl _12197_ (
    .clk(CK),
    .d(\DFF_1533.D ),
    .q(\DFF_1533.Q )
  );
  al_dffl _12198_ (
    .clk(CK),
    .d(\DFF_1534.D ),
    .q(\DFF_1534.Q )
  );
  al_dffl _12199_ (
    .clk(CK),
    .d(\DFF_1535.D ),
    .q(\DFF_1535.Q )
  );
  al_dffl _12200_ (
    .clk(CK),
    .d(\DFF_1536.D ),
    .q(\DFF_1536.Q )
  );
  al_dffl _12201_ (
    .clk(CK),
    .d(\DFF_1537.D ),
    .q(\DFF_1537.Q )
  );
  al_dffl _12202_ (
    .clk(CK),
    .d(\DFF_1538.D ),
    .q(\DFF_1538.Q )
  );
  al_dffl _12203_ (
    .clk(CK),
    .d(\DFF_1539.D ),
    .q(\DFF_1539.Q )
  );
  al_dffl _12204_ (
    .clk(CK),
    .d(\DFF_1540.D ),
    .q(\DFF_1540.Q )
  );
  al_dffl _12205_ (
    .clk(CK),
    .d(\DFF_1541.D ),
    .q(\DFF_1541.Q )
  );
  al_dffl _12206_ (
    .clk(CK),
    .d(\DFF_1542.D ),
    .q(\DFF_1542.Q )
  );
  al_dffl _12207_ (
    .clk(CK),
    .d(\DFF_1543.D ),
    .q(\DFF_1543.Q )
  );
  al_dffl _12208_ (
    .clk(CK),
    .d(\DFF_1544.D ),
    .q(\DFF_1544.Q )
  );
  al_dffl _12209_ (
    .clk(CK),
    .d(\DFF_1545.D ),
    .q(\DFF_1545.Q )
  );
  al_dffl _12210_ (
    .clk(CK),
    .d(\DFF_1546.D ),
    .q(\DFF_1546.Q )
  );
  al_dffl _12211_ (
    .clk(CK),
    .d(\DFF_1547.D ),
    .q(\DFF_1547.Q )
  );
  al_dffl _12212_ (
    .clk(CK),
    .d(\DFF_1548.D ),
    .q(\DFF_1548.Q )
  );
  al_dffl _12213_ (
    .clk(CK),
    .d(\DFF_1549.D ),
    .q(\DFF_1549.Q )
  );
  al_dffl _12214_ (
    .clk(CK),
    .d(\DFF_1550.D ),
    .q(\DFF_1550.Q )
  );
  al_dffl _12215_ (
    .clk(CK),
    .d(\DFF_1551.D ),
    .q(\DFF_1551.Q )
  );
  al_dffl _12216_ (
    .clk(CK),
    .d(\DFF_1552.D ),
    .q(\DFF_1552.Q )
  );
  al_dffl _12217_ (
    .clk(CK),
    .d(\DFF_1553.D ),
    .q(\DFF_1553.Q )
  );
  al_dffl _12218_ (
    .clk(CK),
    .d(\DFF_1554.D ),
    .q(\DFF_1554.Q )
  );
  al_dffl _12219_ (
    .clk(CK),
    .d(\DFF_1555.D ),
    .q(\DFF_1555.Q )
  );
  al_dffl _12220_ (
    .clk(CK),
    .d(\DFF_1556.D ),
    .q(\DFF_1556.Q )
  );
  al_dffl _12221_ (
    .clk(CK),
    .d(\DFF_1557.D ),
    .q(\DFF_1557.Q )
  );
  al_dffl _12222_ (
    .clk(CK),
    .d(\DFF_1558.D ),
    .q(\DFF_1558.Q )
  );
  al_dffl _12223_ (
    .clk(CK),
    .d(\DFF_1559.D ),
    .q(\DFF_1559.Q )
  );
  al_dffl _12224_ (
    .clk(CK),
    .d(\DFF_1560.D ),
    .q(\DFF_1560.Q )
  );
  al_dffl _12225_ (
    .clk(CK),
    .d(\DFF_1561.D ),
    .q(\DFF_1561.Q )
  );
  al_dffl _12226_ (
    .clk(CK),
    .d(\DFF_1562.D ),
    .q(\DFF_1562.Q )
  );
  al_dffl _12227_ (
    .clk(CK),
    .d(\DFF_1563.D ),
    .q(\DFF_1563.Q )
  );
  al_dffl _12228_ (
    .clk(CK),
    .d(\DFF_1564.D ),
    .q(\DFF_1564.Q )
  );
  al_dffl _12229_ (
    .clk(CK),
    .d(\DFF_1565.D ),
    .q(\DFF_1565.Q )
  );
  al_dffl _12230_ (
    .clk(CK),
    .d(\DFF_1566.D ),
    .q(\DFF_1566.Q )
  );
  al_dffl _12231_ (
    .clk(CK),
    .d(\DFF_1567.D ),
    .q(\DFF_1567.Q )
  );
  al_dffl _12232_ (
    .clk(CK),
    .d(\DFF_1568.D ),
    .q(\DFF_1568.Q )
  );
  al_dffl _12233_ (
    .clk(CK),
    .d(\DFF_1569.D ),
    .q(\DFF_1569.Q )
  );
  al_dffl _12234_ (
    .clk(CK),
    .d(\DFF_1570.D ),
    .q(\DFF_1570.Q )
  );
  al_dffl _12235_ (
    .clk(CK),
    .d(\DFF_1571.D ),
    .q(\DFF_1571.Q )
  );
  al_dffl _12236_ (
    .clk(CK),
    .d(\DFF_1572.D ),
    .q(\DFF_1572.Q )
  );
  al_dffl _12237_ (
    .clk(CK),
    .d(\DFF_1573.D ),
    .q(\DFF_1573.Q )
  );
  al_dffl _12238_ (
    .clk(CK),
    .d(\DFF_1574.D ),
    .q(\DFF_1574.Q )
  );
  al_dffl _12239_ (
    .clk(CK),
    .d(\DFF_1575.D ),
    .q(\DFF_1575.Q )
  );
  al_dffl _12240_ (
    .clk(CK),
    .d(\DFF_1576.D ),
    .q(\DFF_1576.Q )
  );
  al_dffl _12241_ (
    .clk(CK),
    .d(\DFF_1577.D ),
    .q(\DFF_1577.Q )
  );
  al_dffl _12242_ (
    .clk(CK),
    .d(\DFF_1578.D ),
    .q(\DFF_1578.Q )
  );
  al_dffl _12243_ (
    .clk(CK),
    .d(\DFF_1579.D ),
    .q(\DFF_1579.Q )
  );
  al_dffl _12244_ (
    .clk(CK),
    .d(\DFF_1580.D ),
    .q(\DFF_1580.Q )
  );
  al_dffl _12245_ (
    .clk(CK),
    .d(\DFF_1581.D ),
    .q(\DFF_1581.Q )
  );
  al_dffl _12246_ (
    .clk(CK),
    .d(\DFF_1582.D ),
    .q(\DFF_1582.Q )
  );
  al_dffl _12247_ (
    .clk(CK),
    .d(\DFF_1583.D ),
    .q(\DFF_1583.Q )
  );
  al_dffl _12248_ (
    .clk(CK),
    .d(\DFF_1584.D ),
    .q(\DFF_1584.Q )
  );
  al_dffl _12249_ (
    .clk(CK),
    .d(\DFF_1585.D ),
    .q(\DFF_1585.Q )
  );
  al_dffl _12250_ (
    .clk(CK),
    .d(\DFF_1586.D ),
    .q(\DFF_1586.Q )
  );
  al_dffl _12251_ (
    .clk(CK),
    .d(\DFF_1587.D ),
    .q(\DFF_1587.Q )
  );
  al_dffl _12252_ (
    .clk(CK),
    .d(\DFF_1588.D ),
    .q(\DFF_1588.Q )
  );
  al_dffl _12253_ (
    .clk(CK),
    .d(\DFF_1589.D ),
    .q(\DFF_1589.Q )
  );
  al_dffl _12254_ (
    .clk(CK),
    .d(\DFF_1590.D ),
    .q(\DFF_1590.Q )
  );
  al_dffl _12255_ (
    .clk(CK),
    .d(\DFF_1591.D ),
    .q(\DFF_1591.Q )
  );
  al_dffl _12256_ (
    .clk(CK),
    .d(\DFF_1592.D ),
    .q(\DFF_1592.Q )
  );
  al_dffl _12257_ (
    .clk(CK),
    .d(\DFF_1593.D ),
    .q(\DFF_1593.Q )
  );
  al_dffl _12258_ (
    .clk(CK),
    .d(\DFF_1594.D ),
    .q(\DFF_1594.Q )
  );
  al_dffl _12259_ (
    .clk(CK),
    .d(\DFF_1595.D ),
    .q(\DFF_1595.Q )
  );
  al_dffl _12260_ (
    .clk(CK),
    .d(\DFF_1596.D ),
    .q(\DFF_1596.Q )
  );
  al_dffl _12261_ (
    .clk(CK),
    .d(\DFF_1597.D ),
    .q(\DFF_1597.Q )
  );
  al_dffl _12262_ (
    .clk(CK),
    .d(\DFF_1598.D ),
    .q(\DFF_1598.Q )
  );
  al_dffl _12263_ (
    .clk(CK),
    .d(\DFF_1599.D ),
    .q(\DFF_1599.Q )
  );
  al_dffl _12264_ (
    .clk(CK),
    .d(\DFF_1600.D ),
    .q(\DFF_1600.Q )
  );
  al_dffl _12265_ (
    .clk(CK),
    .d(\DFF_1601.D ),
    .q(\DFF_1601.Q )
  );
  al_dffl _12266_ (
    .clk(CK),
    .d(\DFF_1602.D ),
    .q(\DFF_1602.Q )
  );
  al_dffl _12267_ (
    .clk(CK),
    .d(\DFF_1603.D ),
    .q(\DFF_1603.Q )
  );
  al_dffl _12268_ (
    .clk(CK),
    .d(\DFF_1604.D ),
    .q(\DFF_1604.Q )
  );
  al_dffl _12269_ (
    .clk(CK),
    .d(\DFF_1605.D ),
    .q(\DFF_1605.Q )
  );
  al_dffl _12270_ (
    .clk(CK),
    .d(\DFF_1606.D ),
    .q(\DFF_1606.Q )
  );
  al_dffl _12271_ (
    .clk(CK),
    .d(\DFF_1607.D ),
    .q(\DFF_1607.Q )
  );
  al_dffl _12272_ (
    .clk(CK),
    .d(\DFF_1608.D ),
    .q(\DFF_1608.Q )
  );
  al_dffl _12273_ (
    .clk(CK),
    .d(\DFF_1609.D ),
    .q(\DFF_1609.Q )
  );
  al_dffl _12274_ (
    .clk(CK),
    .d(\DFF_1610.D ),
    .q(\DFF_1610.Q )
  );
  al_dffl _12275_ (
    .clk(CK),
    .d(\DFF_1611.D ),
    .q(\DFF_1611.Q )
  );
  al_dffl _12276_ (
    .clk(CK),
    .d(\DFF_1612.D ),
    .q(\DFF_1612.Q )
  );
  al_dffl _12277_ (
    .clk(CK),
    .d(\DFF_1613.D ),
    .q(\DFF_1613.Q )
  );
  al_dffl _12278_ (
    .clk(CK),
    .d(\DFF_1614.D ),
    .q(\DFF_1614.Q )
  );
  al_dffl _12279_ (
    .clk(CK),
    .d(\DFF_1615.D ),
    .q(\DFF_1615.Q )
  );
  al_dffl _12280_ (
    .clk(CK),
    .d(\DFF_1616.D ),
    .q(\DFF_1616.Q )
  );
  al_dffl _12281_ (
    .clk(CK),
    .d(\DFF_1617.D ),
    .q(\DFF_1617.Q )
  );
  al_dffl _12282_ (
    .clk(CK),
    .d(\DFF_1618.D ),
    .q(\DFF_1618.Q )
  );
  al_dffl _12283_ (
    .clk(CK),
    .d(\DFF_1619.D ),
    .q(\DFF_1619.Q )
  );
  al_dffl _12284_ (
    .clk(CK),
    .d(\DFF_1620.D ),
    .q(\DFF_1620.Q )
  );
  al_dffl _12285_ (
    .clk(CK),
    .d(\DFF_1621.D ),
    .q(\DFF_1621.Q )
  );
  al_dffl _12286_ (
    .clk(CK),
    .d(\DFF_1622.D ),
    .q(\DFF_1622.Q )
  );
  al_dffl _12287_ (
    .clk(CK),
    .d(\DFF_1623.D ),
    .q(\DFF_1623.Q )
  );
  al_dffl _12288_ (
    .clk(CK),
    .d(\DFF_1624.D ),
    .q(\DFF_1624.Q )
  );
  al_dffl _12289_ (
    .clk(CK),
    .d(\DFF_1625.D ),
    .q(\DFF_1625.Q )
  );
  al_dffl _12290_ (
    .clk(CK),
    .d(\DFF_1626.D ),
    .q(\DFF_1626.Q )
  );
  al_dffl _12291_ (
    .clk(CK),
    .d(\DFF_1627.D ),
    .q(\DFF_1627.Q )
  );
  al_dffl _12292_ (
    .clk(CK),
    .d(\DFF_1628.D ),
    .q(\DFF_1628.Q )
  );
  al_dffl _12293_ (
    .clk(CK),
    .d(\DFF_1629.D ),
    .q(\DFF_1629.Q )
  );
  al_dffl _12294_ (
    .clk(CK),
    .d(\DFF_1630.D ),
    .q(\DFF_1630.Q )
  );
  al_dffl _12295_ (
    .clk(CK),
    .d(\DFF_1631.D ),
    .q(\DFF_1631.Q )
  );
  al_dffl _12296_ (
    .clk(CK),
    .d(\DFF_1632.D ),
    .q(\DFF_1632.Q )
  );
  al_dffl _12297_ (
    .clk(CK),
    .d(\DFF_1633.D ),
    .q(\DFF_1633.Q )
  );
  al_dffl _12298_ (
    .clk(CK),
    .d(\DFF_1634.D ),
    .q(\DFF_1634.Q )
  );
  al_dffl _12299_ (
    .clk(CK),
    .d(\DFF_1635.D ),
    .q(\DFF_1635.Q )
  );
  al_dffl _12300_ (
    .clk(CK),
    .d(\DFF_1636.D ),
    .q(\DFF_1636.Q )
  );
  al_dffl _12301_ (
    .clk(CK),
    .d(\DFF_1637.D ),
    .q(\DFF_1637.Q )
  );
  al_dffl _12302_ (
    .clk(CK),
    .d(\DFF_1638.D ),
    .q(\DFF_1638.Q )
  );
  al_dffl _12303_ (
    .clk(CK),
    .d(\DFF_1639.D ),
    .q(\DFF_1639.Q )
  );
  al_dffl _12304_ (
    .clk(CK),
    .d(\DFF_1640.D ),
    .q(\DFF_1640.Q )
  );
  al_dffl _12305_ (
    .clk(CK),
    .d(\DFF_1641.D ),
    .q(\DFF_1641.Q )
  );
  al_dffl _12306_ (
    .clk(CK),
    .d(\DFF_1642.D ),
    .q(\DFF_1642.Q )
  );
  al_dffl _12307_ (
    .clk(CK),
    .d(\DFF_1643.D ),
    .q(\DFF_1643.Q )
  );
  al_dffl _12308_ (
    .clk(CK),
    .d(\DFF_1644.D ),
    .q(\DFF_1644.Q )
  );
  al_dffl _12309_ (
    .clk(CK),
    .d(\DFF_1645.D ),
    .q(\DFF_1645.Q )
  );
  al_dffl _12310_ (
    .clk(CK),
    .d(\DFF_1646.D ),
    .q(\DFF_1646.Q )
  );
  al_dffl _12311_ (
    .clk(CK),
    .d(\DFF_1647.D ),
    .q(\DFF_1647.Q )
  );
  al_dffl _12312_ (
    .clk(CK),
    .d(\DFF_1648.D ),
    .q(\DFF_1648.Q )
  );
  al_dffl _12313_ (
    .clk(CK),
    .d(\DFF_1649.D ),
    .q(\DFF_1649.Q )
  );
  al_dffl _12314_ (
    .clk(CK),
    .d(\DFF_1650.D ),
    .q(\DFF_1650.Q )
  );
  al_dffl _12315_ (
    .clk(CK),
    .d(\DFF_1651.D ),
    .q(\DFF_1651.Q )
  );
  al_dffl _12316_ (
    .clk(CK),
    .d(\DFF_1652.D ),
    .q(\DFF_1652.Q )
  );
  al_dffl _12317_ (
    .clk(CK),
    .d(\DFF_1653.D ),
    .q(\DFF_1653.Q )
  );
  al_dffl _12318_ (
    .clk(CK),
    .d(\DFF_1654.D ),
    .q(\DFF_1654.Q )
  );
  al_dffl _12319_ (
    .clk(CK),
    .d(\DFF_1655.D ),
    .q(\DFF_1655.Q )
  );
  al_dffl _12320_ (
    .clk(CK),
    .d(\DFF_1656.D ),
    .q(\DFF_1656.Q )
  );
  al_dffl _12321_ (
    .clk(CK),
    .d(\DFF_1657.D ),
    .q(\DFF_1657.Q )
  );
  al_dffl _12322_ (
    .clk(CK),
    .d(\DFF_1658.D ),
    .q(\DFF_1658.Q )
  );
  al_dffl _12323_ (
    .clk(CK),
    .d(\DFF_1659.D ),
    .q(\DFF_1659.Q )
  );
  al_dffl _12324_ (
    .clk(CK),
    .d(\DFF_1660.D ),
    .q(\DFF_1660.Q )
  );
  al_dffl _12325_ (
    .clk(CK),
    .d(\DFF_1661.D ),
    .q(\DFF_1661.Q )
  );
  al_dffl _12326_ (
    .clk(CK),
    .d(\DFF_1662.D ),
    .q(\DFF_1662.Q )
  );
  al_dffl _12327_ (
    .clk(CK),
    .d(\DFF_1663.D ),
    .q(\DFF_1663.Q )
  );
  al_dffl _12328_ (
    .clk(CK),
    .d(\DFF_1664.D ),
    .q(\DFF_1664.Q )
  );
  al_dffl _12329_ (
    .clk(CK),
    .d(\DFF_1665.D ),
    .q(\DFF_1665.Q )
  );
  al_dffl _12330_ (
    .clk(CK),
    .d(\DFF_1666.D ),
    .q(\DFF_1666.Q )
  );
  al_dffl _12331_ (
    .clk(CK),
    .d(\DFF_1667.D ),
    .q(\DFF_1667.Q )
  );
  al_dffl _12332_ (
    .clk(CK),
    .d(\DFF_1668.D ),
    .q(\DFF_1668.Q )
  );
  al_dffl _12333_ (
    .clk(CK),
    .d(\DFF_1669.D ),
    .q(\DFF_1669.Q )
  );
  al_dffl _12334_ (
    .clk(CK),
    .d(\DFF_1670.D ),
    .q(\DFF_1670.Q )
  );
  al_dffl _12335_ (
    .clk(CK),
    .d(\DFF_1671.D ),
    .q(\DFF_1671.Q )
  );
  al_dffl _12336_ (
    .clk(CK),
    .d(\DFF_1672.D ),
    .q(\DFF_1672.Q )
  );
  al_dffl _12337_ (
    .clk(CK),
    .d(\DFF_1673.D ),
    .q(\DFF_1673.Q )
  );
  al_dffl _12338_ (
    .clk(CK),
    .d(\DFF_1674.D ),
    .q(\DFF_1674.Q )
  );
  al_dffl _12339_ (
    .clk(CK),
    .d(\DFF_1675.D ),
    .q(\DFF_1675.Q )
  );
  al_dffl _12340_ (
    .clk(CK),
    .d(\DFF_1676.D ),
    .q(\DFF_1676.Q )
  );
  al_dffl _12341_ (
    .clk(CK),
    .d(\DFF_1677.D ),
    .q(\DFF_1677.Q )
  );
  al_dffl _12342_ (
    .clk(CK),
    .d(\DFF_1678.D ),
    .q(\DFF_1678.Q )
  );
  al_dffl _12343_ (
    .clk(CK),
    .d(\DFF_1679.D ),
    .q(\DFF_1679.Q )
  );
  al_dffl _12344_ (
    .clk(CK),
    .d(\DFF_1680.D ),
    .q(\DFF_1680.Q )
  );
  al_dffl _12345_ (
    .clk(CK),
    .d(\DFF_1681.D ),
    .q(\DFF_1681.Q )
  );
  al_dffl _12346_ (
    .clk(CK),
    .d(\DFF_1682.D ),
    .q(\DFF_1682.Q )
  );
  al_dffl _12347_ (
    .clk(CK),
    .d(\DFF_1683.D ),
    .q(\DFF_1683.Q )
  );
  al_dffl _12348_ (
    .clk(CK),
    .d(\DFF_1684.D ),
    .q(\DFF_1684.Q )
  );
  al_dffl _12349_ (
    .clk(CK),
    .d(\DFF_1685.D ),
    .q(\DFF_1685.Q )
  );
  al_dffl _12350_ (
    .clk(CK),
    .d(\DFF_1686.D ),
    .q(\DFF_1686.Q )
  );
  al_dffl _12351_ (
    .clk(CK),
    .d(\DFF_1687.D ),
    .q(\DFF_1687.Q )
  );
  al_dffl _12352_ (
    .clk(CK),
    .d(\DFF_1688.D ),
    .q(\DFF_1688.Q )
  );
  al_dffl _12353_ (
    .clk(CK),
    .d(\DFF_1689.D ),
    .q(\DFF_1689.Q )
  );
  al_dffl _12354_ (
    .clk(CK),
    .d(\DFF_1690.D ),
    .q(\DFF_1690.Q )
  );
  al_dffl _12355_ (
    .clk(CK),
    .d(\DFF_1691.D ),
    .q(\DFF_1691.Q )
  );
  al_dffl _12356_ (
    .clk(CK),
    .d(\DFF_1692.D ),
    .q(\DFF_1692.Q )
  );
  al_dffl _12357_ (
    .clk(CK),
    .d(\DFF_1693.D ),
    .q(\DFF_1693.Q )
  );
  al_dffl _12358_ (
    .clk(CK),
    .d(\DFF_1694.D ),
    .q(\DFF_1694.Q )
  );
  al_dffl _12359_ (
    .clk(CK),
    .d(\DFF_1695.D ),
    .q(\DFF_1695.Q )
  );
  al_dffl _12360_ (
    .clk(CK),
    .d(\DFF_1696.D ),
    .q(\DFF_1696.Q )
  );
  al_dffl _12361_ (
    .clk(CK),
    .d(\DFF_1697.D ),
    .q(\DFF_1697.Q )
  );
  al_dffl _12362_ (
    .clk(CK),
    .d(\DFF_1698.D ),
    .q(\DFF_1698.Q )
  );
  al_dffl _12363_ (
    .clk(CK),
    .d(\DFF_1699.D ),
    .q(\DFF_1699.Q )
  );
  al_dffl _12364_ (
    .clk(CK),
    .d(\DFF_1700.D ),
    .q(\DFF_1700.Q )
  );
  al_dffl _12365_ (
    .clk(CK),
    .d(\DFF_1701.D ),
    .q(\DFF_1701.Q )
  );
  al_dffl _12366_ (
    .clk(CK),
    .d(\DFF_1702.D ),
    .q(\DFF_1702.Q )
  );
  al_dffl _12367_ (
    .clk(CK),
    .d(\DFF_1703.D ),
    .q(\DFF_1703.Q )
  );
  al_dffl _12368_ (
    .clk(CK),
    .d(\DFF_1704.D ),
    .q(\DFF_1704.Q )
  );
  al_dffl _12369_ (
    .clk(CK),
    .d(\DFF_1705.D ),
    .q(\DFF_1705.Q )
  );
  al_dffl _12370_ (
    .clk(CK),
    .d(\DFF_1706.D ),
    .q(\DFF_1706.Q )
  );
  al_dffl _12371_ (
    .clk(CK),
    .d(\DFF_1707.D ),
    .q(\DFF_1707.Q )
  );
  al_dffl _12372_ (
    .clk(CK),
    .d(\DFF_1708.D ),
    .q(\DFF_1708.Q )
  );
  al_dffl _12373_ (
    .clk(CK),
    .d(\DFF_1709.D ),
    .q(\DFF_1709.Q )
  );
  al_dffl _12374_ (
    .clk(CK),
    .d(\DFF_1710.D ),
    .q(\DFF_1710.Q )
  );
  al_dffl _12375_ (
    .clk(CK),
    .d(\DFF_1711.D ),
    .q(\DFF_1711.Q )
  );
  al_dffl _12376_ (
    .clk(CK),
    .d(\DFF_1712.D ),
    .q(\DFF_1712.Q )
  );
  al_dffl _12377_ (
    .clk(CK),
    .d(\DFF_1713.D ),
    .q(\DFF_1713.Q )
  );
  al_dffl _12378_ (
    .clk(CK),
    .d(\DFF_1714.D ),
    .q(\DFF_1714.Q )
  );
  al_dffl _12379_ (
    .clk(CK),
    .d(\DFF_1715.D ),
    .q(\DFF_1715.Q )
  );
  al_dffl _12380_ (
    .clk(CK),
    .d(\DFF_1716.D ),
    .q(\DFF_1716.Q )
  );
  al_dffl _12381_ (
    .clk(CK),
    .d(\DFF_1717.D ),
    .q(\DFF_1717.Q )
  );
  al_dffl _12382_ (
    .clk(CK),
    .d(\DFF_1718.D ),
    .q(\DFF_1718.Q )
  );
  al_dffl _12383_ (
    .clk(CK),
    .d(\DFF_1719.D ),
    .q(\DFF_1719.Q )
  );
  al_dffl _12384_ (
    .clk(CK),
    .d(\DFF_1720.D ),
    .q(\DFF_1720.Q )
  );
  al_dffl _12385_ (
    .clk(CK),
    .d(\DFF_1721.D ),
    .q(\DFF_1721.Q )
  );
  al_dffl _12386_ (
    .clk(CK),
    .d(\DFF_1722.D ),
    .q(\DFF_1722.Q )
  );
  al_dffl _12387_ (
    .clk(CK),
    .d(\DFF_1723.D ),
    .q(\DFF_1723.Q )
  );
  al_dffl _12388_ (
    .clk(CK),
    .d(\DFF_1724.D ),
    .q(\DFF_1724.Q )
  );
  al_dffl _12389_ (
    .clk(CK),
    .d(\DFF_1725.D ),
    .q(\DFF_1725.Q )
  );
  al_dffl _12390_ (
    .clk(CK),
    .d(\DFF_1726.D ),
    .q(\DFF_1726.Q )
  );
  al_dffl _12391_ (
    .clk(CK),
    .d(\DFF_1727.D ),
    .q(\DFF_1727.Q )
  );
  assign CRC_OUT_1_0 = \DFF_1696.Q ;
  assign CRC_OUT_1_1 = \DFF_1697.Q ;
  assign CRC_OUT_1_10 = \DFF_1706.Q ;
  assign CRC_OUT_1_11 = \DFF_1707.Q ;
  assign CRC_OUT_1_12 = \DFF_1708.Q ;
  assign CRC_OUT_1_13 = \DFF_1709.Q ;
  assign CRC_OUT_1_14 = \DFF_1710.Q ;
  assign CRC_OUT_1_15 = \DFF_1711.Q ;
  assign CRC_OUT_1_16 = \DFF_1712.Q ;
  assign CRC_OUT_1_17 = \DFF_1713.Q ;
  assign CRC_OUT_1_18 = \DFF_1714.Q ;
  assign CRC_OUT_1_19 = \DFF_1715.Q ;
  assign CRC_OUT_1_2 = \DFF_1698.Q ;
  assign CRC_OUT_1_20 = \DFF_1716.Q ;
  assign CRC_OUT_1_21 = \DFF_1717.Q ;
  assign CRC_OUT_1_22 = \DFF_1718.Q ;
  assign CRC_OUT_1_23 = \DFF_1719.Q ;
  assign CRC_OUT_1_24 = \DFF_1720.Q ;
  assign CRC_OUT_1_25 = \DFF_1721.Q ;
  assign CRC_OUT_1_26 = \DFF_1722.Q ;
  assign CRC_OUT_1_27 = \DFF_1723.Q ;
  assign CRC_OUT_1_28 = \DFF_1724.Q ;
  assign CRC_OUT_1_29 = \DFF_1725.Q ;
  assign CRC_OUT_1_3 = \DFF_1699.Q ;
  assign CRC_OUT_1_30 = \DFF_1726.Q ;
  assign CRC_OUT_1_31 = \DFF_1727.Q ;
  assign CRC_OUT_1_4 = \DFF_1700.Q ;
  assign CRC_OUT_1_5 = \DFF_1701.Q ;
  assign CRC_OUT_1_6 = \DFF_1702.Q ;
  assign CRC_OUT_1_7 = \DFF_1703.Q ;
  assign CRC_OUT_1_8 = \DFF_1704.Q ;
  assign CRC_OUT_1_9 = \DFF_1705.Q ;
  assign CRC_OUT_2_0 = \DFF_1504.Q ;
  assign CRC_OUT_2_1 = \DFF_1505.Q ;
  assign CRC_OUT_2_10 = \DFF_1514.Q ;
  assign CRC_OUT_2_11 = \DFF_1515.Q ;
  assign CRC_OUT_2_12 = \DFF_1516.Q ;
  assign CRC_OUT_2_13 = \DFF_1517.Q ;
  assign CRC_OUT_2_14 = \DFF_1518.Q ;
  assign CRC_OUT_2_15 = \DFF_1519.Q ;
  assign CRC_OUT_2_16 = \DFF_1520.Q ;
  assign CRC_OUT_2_17 = \DFF_1521.Q ;
  assign CRC_OUT_2_18 = \DFF_1522.Q ;
  assign CRC_OUT_2_19 = \DFF_1523.Q ;
  assign CRC_OUT_2_2 = \DFF_1506.Q ;
  assign CRC_OUT_2_20 = \DFF_1524.Q ;
  assign CRC_OUT_2_21 = \DFF_1525.Q ;
  assign CRC_OUT_2_22 = \DFF_1526.Q ;
  assign CRC_OUT_2_23 = \DFF_1527.Q ;
  assign CRC_OUT_2_24 = \DFF_1528.Q ;
  assign CRC_OUT_2_25 = \DFF_1529.Q ;
  assign CRC_OUT_2_26 = \DFF_1530.Q ;
  assign CRC_OUT_2_27 = \DFF_1531.Q ;
  assign CRC_OUT_2_28 = \DFF_1532.Q ;
  assign CRC_OUT_2_29 = \DFF_1533.Q ;
  assign CRC_OUT_2_3 = \DFF_1507.Q ;
  assign CRC_OUT_2_30 = \DFF_1534.Q ;
  assign CRC_OUT_2_31 = \DFF_1535.Q ;
  assign CRC_OUT_2_4 = \DFF_1508.Q ;
  assign CRC_OUT_2_5 = \DFF_1509.Q ;
  assign CRC_OUT_2_6 = \DFF_1510.Q ;
  assign CRC_OUT_2_7 = \DFF_1511.Q ;
  assign CRC_OUT_2_8 = \DFF_1512.Q ;
  assign CRC_OUT_2_9 = \DFF_1513.Q ;
  assign CRC_OUT_3_0 = \DFF_1312.Q ;
  assign CRC_OUT_3_1 = \DFF_1313.Q ;
  assign CRC_OUT_3_10 = \DFF_1322.Q ;
  assign CRC_OUT_3_11 = \DFF_1323.Q ;
  assign CRC_OUT_3_12 = \DFF_1324.Q ;
  assign CRC_OUT_3_13 = \DFF_1325.Q ;
  assign CRC_OUT_3_14 = \DFF_1326.Q ;
  assign CRC_OUT_3_15 = \DFF_1327.Q ;
  assign CRC_OUT_3_16 = \DFF_1328.Q ;
  assign CRC_OUT_3_17 = \DFF_1329.Q ;
  assign CRC_OUT_3_18 = \DFF_1330.Q ;
  assign CRC_OUT_3_19 = \DFF_1331.Q ;
  assign CRC_OUT_3_2 = \DFF_1314.Q ;
  assign CRC_OUT_3_20 = \DFF_1332.Q ;
  assign CRC_OUT_3_21 = \DFF_1333.Q ;
  assign CRC_OUT_3_22 = \DFF_1334.Q ;
  assign CRC_OUT_3_23 = \DFF_1335.Q ;
  assign CRC_OUT_3_24 = \DFF_1336.Q ;
  assign CRC_OUT_3_25 = \DFF_1337.Q ;
  assign CRC_OUT_3_26 = \DFF_1338.Q ;
  assign CRC_OUT_3_27 = \DFF_1339.Q ;
  assign CRC_OUT_3_28 = \DFF_1340.Q ;
  assign CRC_OUT_3_29 = \DFF_1341.Q ;
  assign CRC_OUT_3_3 = \DFF_1315.Q ;
  assign CRC_OUT_3_30 = \DFF_1342.Q ;
  assign CRC_OUT_3_31 = \DFF_1343.Q ;
  assign CRC_OUT_3_4 = \DFF_1316.Q ;
  assign CRC_OUT_3_5 = \DFF_1317.Q ;
  assign CRC_OUT_3_6 = \DFF_1318.Q ;
  assign CRC_OUT_3_7 = \DFF_1319.Q ;
  assign CRC_OUT_3_8 = \DFF_1320.Q ;
  assign CRC_OUT_3_9 = \DFF_1321.Q ;
  assign CRC_OUT_4_0 = \DFF_1120.Q ;
  assign CRC_OUT_4_1 = \DFF_1121.Q ;
  assign CRC_OUT_4_10 = \DFF_1130.Q ;
  assign CRC_OUT_4_11 = \DFF_1131.Q ;
  assign CRC_OUT_4_12 = \DFF_1132.Q ;
  assign CRC_OUT_4_13 = \DFF_1133.Q ;
  assign CRC_OUT_4_14 = \DFF_1134.Q ;
  assign CRC_OUT_4_15 = \DFF_1135.Q ;
  assign CRC_OUT_4_16 = \DFF_1136.Q ;
  assign CRC_OUT_4_17 = \DFF_1137.Q ;
  assign CRC_OUT_4_18 = \DFF_1138.Q ;
  assign CRC_OUT_4_19 = \DFF_1139.Q ;
  assign CRC_OUT_4_2 = \DFF_1122.Q ;
  assign CRC_OUT_4_20 = \DFF_1140.Q ;
  assign CRC_OUT_4_21 = \DFF_1141.Q ;
  assign CRC_OUT_4_22 = \DFF_1142.Q ;
  assign CRC_OUT_4_23 = \DFF_1143.Q ;
  assign CRC_OUT_4_24 = \DFF_1144.Q ;
  assign CRC_OUT_4_25 = \DFF_1145.Q ;
  assign CRC_OUT_4_26 = \DFF_1146.Q ;
  assign CRC_OUT_4_27 = \DFF_1147.Q ;
  assign CRC_OUT_4_28 = \DFF_1148.Q ;
  assign CRC_OUT_4_29 = \DFF_1149.Q ;
  assign CRC_OUT_4_3 = \DFF_1123.Q ;
  assign CRC_OUT_4_30 = \DFF_1150.Q ;
  assign CRC_OUT_4_31 = \DFF_1151.Q ;
  assign CRC_OUT_4_4 = \DFF_1124.Q ;
  assign CRC_OUT_4_5 = \DFF_1125.Q ;
  assign CRC_OUT_4_6 = \DFF_1126.Q ;
  assign CRC_OUT_4_7 = \DFF_1127.Q ;
  assign CRC_OUT_4_8 = \DFF_1128.Q ;
  assign CRC_OUT_4_9 = \DFF_1129.Q ;
  assign CRC_OUT_5_0 = \DFF_928.Q ;
  assign CRC_OUT_5_1 = \DFF_929.Q ;
  assign CRC_OUT_5_10 = \DFF_938.Q ;
  assign CRC_OUT_5_11 = \DFF_939.Q ;
  assign CRC_OUT_5_12 = \DFF_940.Q ;
  assign CRC_OUT_5_13 = \DFF_941.Q ;
  assign CRC_OUT_5_14 = \DFF_942.Q ;
  assign CRC_OUT_5_15 = \DFF_943.Q ;
  assign CRC_OUT_5_16 = \DFF_944.Q ;
  assign CRC_OUT_5_17 = \DFF_945.Q ;
  assign CRC_OUT_5_18 = \DFF_946.Q ;
  assign CRC_OUT_5_19 = \DFF_947.Q ;
  assign CRC_OUT_5_2 = \DFF_930.Q ;
  assign CRC_OUT_5_20 = \DFF_948.Q ;
  assign CRC_OUT_5_21 = \DFF_949.Q ;
  assign CRC_OUT_5_22 = \DFF_950.Q ;
  assign CRC_OUT_5_23 = \DFF_951.Q ;
  assign CRC_OUT_5_24 = \DFF_952.Q ;
  assign CRC_OUT_5_25 = \DFF_953.Q ;
  assign CRC_OUT_5_26 = \DFF_954.Q ;
  assign CRC_OUT_5_27 = \DFF_955.Q ;
  assign CRC_OUT_5_28 = \DFF_956.Q ;
  assign CRC_OUT_5_29 = \DFF_957.Q ;
  assign CRC_OUT_5_3 = \DFF_931.Q ;
  assign CRC_OUT_5_30 = \DFF_958.Q ;
  assign CRC_OUT_5_31 = \DFF_959.Q ;
  assign CRC_OUT_5_4 = \DFF_932.Q ;
  assign CRC_OUT_5_5 = \DFF_933.Q ;
  assign CRC_OUT_5_6 = \DFF_934.Q ;
  assign CRC_OUT_5_7 = \DFF_935.Q ;
  assign CRC_OUT_5_8 = \DFF_936.Q ;
  assign CRC_OUT_5_9 = \DFF_937.Q ;
  assign CRC_OUT_6_0 = \DFF_736.Q ;
  assign CRC_OUT_6_1 = \DFF_737.Q ;
  assign CRC_OUT_6_10 = \DFF_746.Q ;
  assign CRC_OUT_6_11 = \DFF_747.Q ;
  assign CRC_OUT_6_12 = \DFF_748.Q ;
  assign CRC_OUT_6_13 = \DFF_749.Q ;
  assign CRC_OUT_6_14 = \DFF_750.Q ;
  assign CRC_OUT_6_15 = \DFF_751.Q ;
  assign CRC_OUT_6_16 = \DFF_752.Q ;
  assign CRC_OUT_6_17 = \DFF_753.Q ;
  assign CRC_OUT_6_18 = \DFF_754.Q ;
  assign CRC_OUT_6_19 = \DFF_755.Q ;
  assign CRC_OUT_6_2 = \DFF_738.Q ;
  assign CRC_OUT_6_20 = \DFF_756.Q ;
  assign CRC_OUT_6_21 = \DFF_757.Q ;
  assign CRC_OUT_6_22 = \DFF_758.Q ;
  assign CRC_OUT_6_23 = \DFF_759.Q ;
  assign CRC_OUT_6_24 = \DFF_760.Q ;
  assign CRC_OUT_6_25 = \DFF_761.Q ;
  assign CRC_OUT_6_26 = \DFF_762.Q ;
  assign CRC_OUT_6_27 = \DFF_763.Q ;
  assign CRC_OUT_6_28 = \DFF_764.Q ;
  assign CRC_OUT_6_29 = \DFF_765.Q ;
  assign CRC_OUT_6_3 = \DFF_739.Q ;
  assign CRC_OUT_6_30 = \DFF_766.Q ;
  assign CRC_OUT_6_31 = \DFF_767.Q ;
  assign CRC_OUT_6_4 = \DFF_740.Q ;
  assign CRC_OUT_6_5 = \DFF_741.Q ;
  assign CRC_OUT_6_6 = \DFF_742.Q ;
  assign CRC_OUT_6_7 = \DFF_743.Q ;
  assign CRC_OUT_6_8 = \DFF_744.Q ;
  assign CRC_OUT_6_9 = \DFF_745.Q ;
  assign CRC_OUT_7_0 = \DFF_544.Q ;
  assign CRC_OUT_7_1 = \DFF_545.Q ;
  assign CRC_OUT_7_10 = \DFF_554.Q ;
  assign CRC_OUT_7_11 = \DFF_555.Q ;
  assign CRC_OUT_7_12 = \DFF_556.Q ;
  assign CRC_OUT_7_13 = \DFF_557.Q ;
  assign CRC_OUT_7_14 = \DFF_558.Q ;
  assign CRC_OUT_7_15 = \DFF_559.Q ;
  assign CRC_OUT_7_16 = \DFF_560.Q ;
  assign CRC_OUT_7_17 = \DFF_561.Q ;
  assign CRC_OUT_7_18 = \DFF_562.Q ;
  assign CRC_OUT_7_19 = \DFF_563.Q ;
  assign CRC_OUT_7_2 = \DFF_546.Q ;
  assign CRC_OUT_7_20 = \DFF_564.Q ;
  assign CRC_OUT_7_21 = \DFF_565.Q ;
  assign CRC_OUT_7_22 = \DFF_566.Q ;
  assign CRC_OUT_7_23 = \DFF_567.Q ;
  assign CRC_OUT_7_24 = \DFF_568.Q ;
  assign CRC_OUT_7_25 = \DFF_569.Q ;
  assign CRC_OUT_7_26 = \DFF_570.Q ;
  assign CRC_OUT_7_27 = \DFF_571.Q ;
  assign CRC_OUT_7_28 = \DFF_572.Q ;
  assign CRC_OUT_7_29 = \DFF_573.Q ;
  assign CRC_OUT_7_3 = \DFF_547.Q ;
  assign CRC_OUT_7_30 = \DFF_574.Q ;
  assign CRC_OUT_7_31 = \DFF_575.Q ;
  assign CRC_OUT_7_4 = \DFF_548.Q ;
  assign CRC_OUT_7_5 = \DFF_549.Q ;
  assign CRC_OUT_7_6 = \DFF_550.Q ;
  assign CRC_OUT_7_7 = \DFF_551.Q ;
  assign CRC_OUT_7_8 = \DFF_552.Q ;
  assign CRC_OUT_7_9 = \DFF_553.Q ;
  assign CRC_OUT_8_0 = \DFF_352.Q ;
  assign CRC_OUT_8_1 = \DFF_353.Q ;
  assign CRC_OUT_8_10 = \DFF_362.Q ;
  assign CRC_OUT_8_11 = \DFF_363.Q ;
  assign CRC_OUT_8_12 = \DFF_364.Q ;
  assign CRC_OUT_8_13 = \DFF_365.Q ;
  assign CRC_OUT_8_14 = \DFF_366.Q ;
  assign CRC_OUT_8_15 = \DFF_367.Q ;
  assign CRC_OUT_8_16 = \DFF_368.Q ;
  assign CRC_OUT_8_17 = \DFF_369.Q ;
  assign CRC_OUT_8_18 = \DFF_370.Q ;
  assign CRC_OUT_8_19 = \DFF_371.Q ;
  assign CRC_OUT_8_2 = \DFF_354.Q ;
  assign CRC_OUT_8_20 = \DFF_372.Q ;
  assign CRC_OUT_8_21 = \DFF_373.Q ;
  assign CRC_OUT_8_22 = \DFF_374.Q ;
  assign CRC_OUT_8_23 = \DFF_375.Q ;
  assign CRC_OUT_8_24 = \DFF_376.Q ;
  assign CRC_OUT_8_25 = \DFF_377.Q ;
  assign CRC_OUT_8_26 = \DFF_378.Q ;
  assign CRC_OUT_8_27 = \DFF_379.Q ;
  assign CRC_OUT_8_28 = \DFF_380.Q ;
  assign CRC_OUT_8_29 = \DFF_381.Q ;
  assign CRC_OUT_8_3 = \DFF_355.Q ;
  assign CRC_OUT_8_30 = \DFF_382.Q ;
  assign CRC_OUT_8_31 = \DFF_383.Q ;
  assign CRC_OUT_8_4 = \DFF_356.Q ;
  assign CRC_OUT_8_5 = \DFF_357.Q ;
  assign CRC_OUT_8_6 = \DFF_358.Q ;
  assign CRC_OUT_8_7 = \DFF_359.Q ;
  assign CRC_OUT_8_8 = \DFF_360.Q ;
  assign CRC_OUT_8_9 = \DFF_361.Q ;
  assign CRC_OUT_9_0 = \DFF_160.Q ;
  assign CRC_OUT_9_1 = \DFF_161.Q ;
  assign CRC_OUT_9_10 = \DFF_170.Q ;
  assign CRC_OUT_9_11 = \DFF_171.Q ;
  assign CRC_OUT_9_12 = \DFF_172.Q ;
  assign CRC_OUT_9_13 = \DFF_173.Q ;
  assign CRC_OUT_9_14 = \DFF_174.Q ;
  assign CRC_OUT_9_15 = \DFF_175.Q ;
  assign CRC_OUT_9_16 = \DFF_176.Q ;
  assign CRC_OUT_9_17 = \DFF_177.Q ;
  assign CRC_OUT_9_18 = \DFF_178.Q ;
  assign CRC_OUT_9_19 = \DFF_179.Q ;
  assign CRC_OUT_9_2 = \DFF_162.Q ;
  assign CRC_OUT_9_20 = \DFF_180.Q ;
  assign CRC_OUT_9_21 = \DFF_181.Q ;
  assign CRC_OUT_9_22 = \DFF_182.Q ;
  assign CRC_OUT_9_23 = \DFF_183.Q ;
  assign CRC_OUT_9_24 = \DFF_184.Q ;
  assign CRC_OUT_9_25 = \DFF_185.Q ;
  assign CRC_OUT_9_26 = \DFF_186.Q ;
  assign CRC_OUT_9_27 = \DFF_187.Q ;
  assign CRC_OUT_9_28 = \DFF_188.Q ;
  assign CRC_OUT_9_29 = \DFF_189.Q ;
  assign CRC_OUT_9_3 = \DFF_163.Q ;
  assign CRC_OUT_9_30 = \DFF_190.Q ;
  assign CRC_OUT_9_31 = \DFF_191.Q ;
  assign CRC_OUT_9_4 = \DFF_164.Q ;
  assign CRC_OUT_9_5 = \DFF_165.Q ;
  assign CRC_OUT_9_6 = \DFF_166.Q ;
  assign CRC_OUT_9_7 = \DFF_167.Q ;
  assign CRC_OUT_9_8 = \DFF_168.Q ;
  assign CRC_OUT_9_9 = \DFF_169.Q ;
  assign \DFF_0.CK  = CK;
  assign \DFF_1.CK  = CK;
  assign \DFF_10.CK  = CK;
  assign \DFF_100.CK  = CK;
  assign \DFF_1000.CK  = CK;
  assign \DFF_1001.CK  = CK;
  assign \DFF_1002.CK  = CK;
  assign \DFF_1003.CK  = CK;
  assign \DFF_1004.CK  = CK;
  assign \DFF_1005.CK  = CK;
  assign \DFF_1006.CK  = CK;
  assign \DFF_1007.CK  = CK;
  assign \DFF_1008.CK  = CK;
  assign \DFF_1009.CK  = CK;
  assign \DFF_101.CK  = CK;
  assign \DFF_1010.CK  = CK;
  assign \DFF_1011.CK  = CK;
  assign \DFF_1012.CK  = CK;
  assign \DFF_1013.CK  = CK;
  assign \DFF_1014.CK  = CK;
  assign \DFF_1015.CK  = CK;
  assign \DFF_1016.CK  = CK;
  assign \DFF_1017.CK  = CK;
  assign \DFF_1018.CK  = CK;
  assign \DFF_1019.CK  = CK;
  assign \DFF_102.CK  = CK;
  assign \DFF_1020.CK  = CK;
  assign \DFF_1021.CK  = CK;
  assign \DFF_1022.CK  = CK;
  assign \DFF_1023.CK  = CK;
  assign \DFF_1024.CK  = CK;
  assign \DFF_1025.CK  = CK;
  assign \DFF_1026.CK  = CK;
  assign \DFF_1027.CK  = CK;
  assign \DFF_1028.CK  = CK;
  assign \DFF_1029.CK  = CK;
  assign \DFF_103.CK  = CK;
  assign \DFF_1030.CK  = CK;
  assign \DFF_1031.CK  = CK;
  assign \DFF_1032.CK  = CK;
  assign \DFF_1033.CK  = CK;
  assign \DFF_1034.CK  = CK;
  assign \DFF_1035.CK  = CK;
  assign \DFF_1036.CK  = CK;
  assign \DFF_1037.CK  = CK;
  assign \DFF_1038.CK  = CK;
  assign \DFF_1039.CK  = CK;
  assign \DFF_104.CK  = CK;
  assign \DFF_1040.CK  = CK;
  assign \DFF_1041.CK  = CK;
  assign \DFF_1042.CK  = CK;
  assign \DFF_1043.CK  = CK;
  assign \DFF_1044.CK  = CK;
  assign \DFF_1045.CK  = CK;
  assign \DFF_1046.CK  = CK;
  assign \DFF_1047.CK  = CK;
  assign \DFF_1048.CK  = CK;
  assign \DFF_1049.CK  = CK;
  assign \DFF_105.CK  = CK;
  assign \DFF_1050.CK  = CK;
  assign \DFF_1051.CK  = CK;
  assign \DFF_1052.CK  = CK;
  assign \DFF_1053.CK  = CK;
  assign \DFF_1054.CK  = CK;
  assign \DFF_1055.CK  = CK;
  assign \DFF_1056.CK  = CK;
  assign \DFF_1057.CK  = CK;
  assign \DFF_1058.CK  = CK;
  assign \DFF_1059.CK  = CK;
  assign \DFF_106.CK  = CK;
  assign \DFF_1060.CK  = CK;
  assign \DFF_1061.CK  = CK;
  assign \DFF_1062.CK  = CK;
  assign \DFF_1063.CK  = CK;
  assign \DFF_1064.CK  = CK;
  assign \DFF_1065.CK  = CK;
  assign \DFF_1066.CK  = CK;
  assign \DFF_1067.CK  = CK;
  assign \DFF_1068.CK  = CK;
  assign \DFF_1069.CK  = CK;
  assign \DFF_107.CK  = CK;
  assign \DFF_1070.CK  = CK;
  assign \DFF_1071.CK  = CK;
  assign \DFF_1072.CK  = CK;
  assign \DFF_1073.CK  = CK;
  assign \DFF_1074.CK  = CK;
  assign \DFF_1075.CK  = CK;
  assign \DFF_1076.CK  = CK;
  assign \DFF_1077.CK  = CK;
  assign \DFF_1078.CK  = CK;
  assign \DFF_1079.CK  = CK;
  assign \DFF_108.CK  = CK;
  assign \DFF_1080.CK  = CK;
  assign \DFF_1081.CK  = CK;
  assign \DFF_1082.CK  = CK;
  assign \DFF_1083.CK  = CK;
  assign \DFF_1084.CK  = CK;
  assign \DFF_1085.CK  = CK;
  assign \DFF_1086.CK  = CK;
  assign \DFF_1087.CK  = CK;
  assign \DFF_1088.CK  = CK;
  assign \DFF_1089.CK  = CK;
  assign \DFF_109.CK  = CK;
  assign \DFF_1090.CK  = CK;
  assign \DFF_1091.CK  = CK;
  assign \DFF_1092.CK  = CK;
  assign \DFF_1093.CK  = CK;
  assign \DFF_1094.CK  = CK;
  assign \DFF_1095.CK  = CK;
  assign \DFF_1096.CK  = CK;
  assign \DFF_1097.CK  = CK;
  assign \DFF_1098.CK  = CK;
  assign \DFF_1099.CK  = CK;
  assign \DFF_11.CK  = CK;
  assign \DFF_110.CK  = CK;
  assign \DFF_1100.CK  = CK;
  assign \DFF_1101.CK  = CK;
  assign \DFF_1102.CK  = CK;
  assign \DFF_1103.CK  = CK;
  assign \DFF_1104.CK  = CK;
  assign \DFF_1105.CK  = CK;
  assign \DFF_1106.CK  = CK;
  assign \DFF_1107.CK  = CK;
  assign \DFF_1108.CK  = CK;
  assign \DFF_1109.CK  = CK;
  assign \DFF_111.CK  = CK;
  assign \DFF_1110.CK  = CK;
  assign \DFF_1111.CK  = CK;
  assign \DFF_1112.CK  = CK;
  assign \DFF_1113.CK  = CK;
  assign \DFF_1114.CK  = CK;
  assign \DFF_1115.CK  = CK;
  assign \DFF_1116.CK  = CK;
  assign \DFF_1117.CK  = CK;
  assign \DFF_1118.CK  = CK;
  assign \DFF_1119.CK  = CK;
  assign \DFF_112.CK  = CK;
  assign \DFF_1120.CK  = CK;
  assign \DFF_1121.CK  = CK;
  assign \DFF_1122.CK  = CK;
  assign \DFF_1123.CK  = CK;
  assign \DFF_1124.CK  = CK;
  assign \DFF_1125.CK  = CK;
  assign \DFF_1126.CK  = CK;
  assign \DFF_1127.CK  = CK;
  assign \DFF_1128.CK  = CK;
  assign \DFF_1129.CK  = CK;
  assign \DFF_113.CK  = CK;
  assign \DFF_1130.CK  = CK;
  assign \DFF_1131.CK  = CK;
  assign \DFF_1132.CK  = CK;
  assign \DFF_1133.CK  = CK;
  assign \DFF_1134.CK  = CK;
  assign \DFF_1135.CK  = CK;
  assign \DFF_1136.CK  = CK;
  assign \DFF_1137.CK  = CK;
  assign \DFF_1138.CK  = CK;
  assign \DFF_1139.CK  = CK;
  assign \DFF_114.CK  = CK;
  assign \DFF_1140.CK  = CK;
  assign \DFF_1141.CK  = CK;
  assign \DFF_1142.CK  = CK;
  assign \DFF_1143.CK  = CK;
  assign \DFF_1144.CK  = CK;
  assign \DFF_1145.CK  = CK;
  assign \DFF_1146.CK  = CK;
  assign \DFF_1147.CK  = CK;
  assign \DFF_1148.CK  = CK;
  assign \DFF_1149.CK  = CK;
  assign \DFF_115.CK  = CK;
  assign \DFF_1150.CK  = CK;
  assign \DFF_1151.CK  = CK;
  assign \DFF_1152.CK  = CK;
  assign \DFF_1153.CK  = CK;
  assign \DFF_1154.CK  = CK;
  assign \DFF_1155.CK  = CK;
  assign \DFF_1156.CK  = CK;
  assign \DFF_1157.CK  = CK;
  assign \DFF_1158.CK  = CK;
  assign \DFF_1159.CK  = CK;
  assign \DFF_116.CK  = CK;
  assign \DFF_1160.CK  = CK;
  assign \DFF_1161.CK  = CK;
  assign \DFF_1162.CK  = CK;
  assign \DFF_1163.CK  = CK;
  assign \DFF_1164.CK  = CK;
  assign \DFF_1165.CK  = CK;
  assign \DFF_1166.CK  = CK;
  assign \DFF_1167.CK  = CK;
  assign \DFF_1168.CK  = CK;
  assign \DFF_1169.CK  = CK;
  assign \DFF_117.CK  = CK;
  assign \DFF_1170.CK  = CK;
  assign \DFF_1171.CK  = CK;
  assign \DFF_1172.CK  = CK;
  assign \DFF_1173.CK  = CK;
  assign \DFF_1174.CK  = CK;
  assign \DFF_1175.CK  = CK;
  assign \DFF_1176.CK  = CK;
  assign \DFF_1177.CK  = CK;
  assign \DFF_1178.CK  = CK;
  assign \DFF_1179.CK  = CK;
  assign \DFF_118.CK  = CK;
  assign \DFF_1180.CK  = CK;
  assign \DFF_1181.CK  = CK;
  assign \DFF_1182.CK  = CK;
  assign \DFF_1183.CK  = CK;
  assign \DFF_1184.CK  = CK;
  assign \DFF_1185.CK  = CK;
  assign \DFF_1186.CK  = CK;
  assign \DFF_1187.CK  = CK;
  assign \DFF_1188.CK  = CK;
  assign \DFF_1189.CK  = CK;
  assign \DFF_119.CK  = CK;
  assign \DFF_1190.CK  = CK;
  assign \DFF_1191.CK  = CK;
  assign \DFF_1192.CK  = CK;
  assign \DFF_1193.CK  = CK;
  assign \DFF_1194.CK  = CK;
  assign \DFF_1195.CK  = CK;
  assign \DFF_1196.CK  = CK;
  assign \DFF_1197.CK  = CK;
  assign \DFF_1198.CK  = CK;
  assign \DFF_1199.CK  = CK;
  assign \DFF_12.CK  = CK;
  assign \DFF_120.CK  = CK;
  assign \DFF_1200.CK  = CK;
  assign \DFF_1201.CK  = CK;
  assign \DFF_1202.CK  = CK;
  assign \DFF_1203.CK  = CK;
  assign \DFF_1204.CK  = CK;
  assign \DFF_1205.CK  = CK;
  assign \DFF_1206.CK  = CK;
  assign \DFF_1207.CK  = CK;
  assign \DFF_1208.CK  = CK;
  assign \DFF_1209.CK  = CK;
  assign \DFF_121.CK  = CK;
  assign \DFF_1210.CK  = CK;
  assign \DFF_1211.CK  = CK;
  assign \DFF_1212.CK  = CK;
  assign \DFF_1213.CK  = CK;
  assign \DFF_1214.CK  = CK;
  assign \DFF_1215.CK  = CK;
  assign \DFF_1216.CK  = CK;
  assign \DFF_1217.CK  = CK;
  assign \DFF_1218.CK  = CK;
  assign \DFF_1219.CK  = CK;
  assign \DFF_122.CK  = CK;
  assign \DFF_1220.CK  = CK;
  assign \DFF_1221.CK  = CK;
  assign \DFF_1222.CK  = CK;
  assign \DFF_1223.CK  = CK;
  assign \DFF_1224.CK  = CK;
  assign \DFF_1225.CK  = CK;
  assign \DFF_1226.CK  = CK;
  assign \DFF_1227.CK  = CK;
  assign \DFF_1228.CK  = CK;
  assign \DFF_1229.CK  = CK;
  assign \DFF_123.CK  = CK;
  assign \DFF_1230.CK  = CK;
  assign \DFF_1231.CK  = CK;
  assign \DFF_1232.CK  = CK;
  assign \DFF_1233.CK  = CK;
  assign \DFF_1234.CK  = CK;
  assign \DFF_1235.CK  = CK;
  assign \DFF_1236.CK  = CK;
  assign \DFF_1237.CK  = CK;
  assign \DFF_1238.CK  = CK;
  assign \DFF_1239.CK  = CK;
  assign \DFF_124.CK  = CK;
  assign \DFF_1240.CK  = CK;
  assign \DFF_1241.CK  = CK;
  assign \DFF_1242.CK  = CK;
  assign \DFF_1243.CK  = CK;
  assign \DFF_1244.CK  = CK;
  assign \DFF_1245.CK  = CK;
  assign \DFF_1246.CK  = CK;
  assign \DFF_1247.CK  = CK;
  assign \DFF_1248.CK  = CK;
  assign \DFF_1249.CK  = CK;
  assign \DFF_125.CK  = CK;
  assign \DFF_1250.CK  = CK;
  assign \DFF_1251.CK  = CK;
  assign \DFF_1252.CK  = CK;
  assign \DFF_1253.CK  = CK;
  assign \DFF_1254.CK  = CK;
  assign \DFF_1255.CK  = CK;
  assign \DFF_1256.CK  = CK;
  assign \DFF_1257.CK  = CK;
  assign \DFF_1258.CK  = CK;
  assign \DFF_1259.CK  = CK;
  assign \DFF_126.CK  = CK;
  assign \DFF_1260.CK  = CK;
  assign \DFF_1261.CK  = CK;
  assign \DFF_1262.CK  = CK;
  assign \DFF_1263.CK  = CK;
  assign \DFF_1264.CK  = CK;
  assign \DFF_1265.CK  = CK;
  assign \DFF_1266.CK  = CK;
  assign \DFF_1267.CK  = CK;
  assign \DFF_1268.CK  = CK;
  assign \DFF_1269.CK  = CK;
  assign \DFF_127.CK  = CK;
  assign \DFF_1270.CK  = CK;
  assign \DFF_1271.CK  = CK;
  assign \DFF_1272.CK  = CK;
  assign \DFF_1273.CK  = CK;
  assign \DFF_1274.CK  = CK;
  assign \DFF_1275.CK  = CK;
  assign \DFF_1276.CK  = CK;
  assign \DFF_1277.CK  = CK;
  assign \DFF_1278.CK  = CK;
  assign \DFF_1279.CK  = CK;
  assign \DFF_128.CK  = CK;
  assign \DFF_1280.CK  = CK;
  assign \DFF_1281.CK  = CK;
  assign \DFF_1282.CK  = CK;
  assign \DFF_1283.CK  = CK;
  assign \DFF_1284.CK  = CK;
  assign \DFF_1285.CK  = CK;
  assign \DFF_1286.CK  = CK;
  assign \DFF_1287.CK  = CK;
  assign \DFF_1288.CK  = CK;
  assign \DFF_1289.CK  = CK;
  assign \DFF_129.CK  = CK;
  assign \DFF_1290.CK  = CK;
  assign \DFF_1291.CK  = CK;
  assign \DFF_1292.CK  = CK;
  assign \DFF_1293.CK  = CK;
  assign \DFF_1294.CK  = CK;
  assign \DFF_1295.CK  = CK;
  assign \DFF_1296.CK  = CK;
  assign \DFF_1297.CK  = CK;
  assign \DFF_1298.CK  = CK;
  assign \DFF_1299.CK  = CK;
  assign \DFF_13.CK  = CK;
  assign \DFF_130.CK  = CK;
  assign \DFF_1300.CK  = CK;
  assign \DFF_1301.CK  = CK;
  assign \DFF_1302.CK  = CK;
  assign \DFF_1303.CK  = CK;
  assign \DFF_1304.CK  = CK;
  assign \DFF_1305.CK  = CK;
  assign \DFF_1306.CK  = CK;
  assign \DFF_1307.CK  = CK;
  assign \DFF_1308.CK  = CK;
  assign \DFF_1309.CK  = CK;
  assign \DFF_131.CK  = CK;
  assign \DFF_1310.CK  = CK;
  assign \DFF_1311.CK  = CK;
  assign \DFF_1312.CK  = CK;
  assign \DFF_1313.CK  = CK;
  assign \DFF_1314.CK  = CK;
  assign \DFF_1315.CK  = CK;
  assign \DFF_1316.CK  = CK;
  assign \DFF_1317.CK  = CK;
  assign \DFF_1318.CK  = CK;
  assign \DFF_1319.CK  = CK;
  assign \DFF_132.CK  = CK;
  assign \DFF_1320.CK  = CK;
  assign \DFF_1321.CK  = CK;
  assign \DFF_1322.CK  = CK;
  assign \DFF_1323.CK  = CK;
  assign \DFF_1324.CK  = CK;
  assign \DFF_1325.CK  = CK;
  assign \DFF_1326.CK  = CK;
  assign \DFF_1327.CK  = CK;
  assign \DFF_1328.CK  = CK;
  assign \DFF_1329.CK  = CK;
  assign \DFF_133.CK  = CK;
  assign \DFF_1330.CK  = CK;
  assign \DFF_1331.CK  = CK;
  assign \DFF_1332.CK  = CK;
  assign \DFF_1333.CK  = CK;
  assign \DFF_1334.CK  = CK;
  assign \DFF_1335.CK  = CK;
  assign \DFF_1336.CK  = CK;
  assign \DFF_1337.CK  = CK;
  assign \DFF_1338.CK  = CK;
  assign \DFF_1339.CK  = CK;
  assign \DFF_134.CK  = CK;
  assign \DFF_1340.CK  = CK;
  assign \DFF_1341.CK  = CK;
  assign \DFF_1342.CK  = CK;
  assign \DFF_1343.CK  = CK;
  assign \DFF_1344.CK  = CK;
  assign \DFF_1345.CK  = CK;
  assign \DFF_1346.CK  = CK;
  assign \DFF_1347.CK  = CK;
  assign \DFF_1348.CK  = CK;
  assign \DFF_1349.CK  = CK;
  assign \DFF_135.CK  = CK;
  assign \DFF_1350.CK  = CK;
  assign \DFF_1351.CK  = CK;
  assign \DFF_1352.CK  = CK;
  assign \DFF_1353.CK  = CK;
  assign \DFF_1354.CK  = CK;
  assign \DFF_1355.CK  = CK;
  assign \DFF_1356.CK  = CK;
  assign \DFF_1357.CK  = CK;
  assign \DFF_1358.CK  = CK;
  assign \DFF_1359.CK  = CK;
  assign \DFF_136.CK  = CK;
  assign \DFF_1360.CK  = CK;
  assign \DFF_1361.CK  = CK;
  assign \DFF_1362.CK  = CK;
  assign \DFF_1363.CK  = CK;
  assign \DFF_1364.CK  = CK;
  assign \DFF_1365.CK  = CK;
  assign \DFF_1366.CK  = CK;
  assign \DFF_1367.CK  = CK;
  assign \DFF_1368.CK  = CK;
  assign \DFF_1369.CK  = CK;
  assign \DFF_137.CK  = CK;
  assign \DFF_1370.CK  = CK;
  assign \DFF_1371.CK  = CK;
  assign \DFF_1372.CK  = CK;
  assign \DFF_1373.CK  = CK;
  assign \DFF_1374.CK  = CK;
  assign \DFF_1375.CK  = CK;
  assign \DFF_1376.CK  = CK;
  assign \DFF_1377.CK  = CK;
  assign \DFF_1378.CK  = CK;
  assign \DFF_1379.CK  = CK;
  assign \DFF_138.CK  = CK;
  assign \DFF_1380.CK  = CK;
  assign \DFF_1381.CK  = CK;
  assign \DFF_1382.CK  = CK;
  assign \DFF_1383.CK  = CK;
  assign \DFF_1384.CK  = CK;
  assign \DFF_1385.CK  = CK;
  assign \DFF_1386.CK  = CK;
  assign \DFF_1387.CK  = CK;
  assign \DFF_1388.CK  = CK;
  assign \DFF_1389.CK  = CK;
  assign \DFF_139.CK  = CK;
  assign \DFF_1390.CK  = CK;
  assign \DFF_1391.CK  = CK;
  assign \DFF_1392.CK  = CK;
  assign \DFF_1393.CK  = CK;
  assign \DFF_1394.CK  = CK;
  assign \DFF_1395.CK  = CK;
  assign \DFF_1396.CK  = CK;
  assign \DFF_1397.CK  = CK;
  assign \DFF_1398.CK  = CK;
  assign \DFF_1399.CK  = CK;
  assign \DFF_14.CK  = CK;
  assign \DFF_140.CK  = CK;
  assign \DFF_1400.CK  = CK;
  assign \DFF_1401.CK  = CK;
  assign \DFF_1402.CK  = CK;
  assign \DFF_1403.CK  = CK;
  assign \DFF_1404.CK  = CK;
  assign \DFF_1405.CK  = CK;
  assign \DFF_1406.CK  = CK;
  assign \DFF_1407.CK  = CK;
  assign \DFF_1408.CK  = CK;
  assign \DFF_1409.CK  = CK;
  assign \DFF_141.CK  = CK;
  assign \DFF_1410.CK  = CK;
  assign \DFF_1411.CK  = CK;
  assign \DFF_1412.CK  = CK;
  assign \DFF_1413.CK  = CK;
  assign \DFF_1414.CK  = CK;
  assign \DFF_1415.CK  = CK;
  assign \DFF_1416.CK  = CK;
  assign \DFF_1417.CK  = CK;
  assign \DFF_1418.CK  = CK;
  assign \DFF_1419.CK  = CK;
  assign \DFF_142.CK  = CK;
  assign \DFF_1420.CK  = CK;
  assign \DFF_1421.CK  = CK;
  assign \DFF_1422.CK  = CK;
  assign \DFF_1423.CK  = CK;
  assign \DFF_1424.CK  = CK;
  assign \DFF_1425.CK  = CK;
  assign \DFF_1426.CK  = CK;
  assign \DFF_1427.CK  = CK;
  assign \DFF_1428.CK  = CK;
  assign \DFF_1429.CK  = CK;
  assign \DFF_143.CK  = CK;
  assign \DFF_1430.CK  = CK;
  assign \DFF_1431.CK  = CK;
  assign \DFF_1432.CK  = CK;
  assign \DFF_1433.CK  = CK;
  assign \DFF_1434.CK  = CK;
  assign \DFF_1435.CK  = CK;
  assign \DFF_1436.CK  = CK;
  assign \DFF_1437.CK  = CK;
  assign \DFF_1438.CK  = CK;
  assign \DFF_1439.CK  = CK;
  assign \DFF_144.CK  = CK;
  assign \DFF_1440.CK  = CK;
  assign \DFF_1441.CK  = CK;
  assign \DFF_1442.CK  = CK;
  assign \DFF_1443.CK  = CK;
  assign \DFF_1444.CK  = CK;
  assign \DFF_1445.CK  = CK;
  assign \DFF_1446.CK  = CK;
  assign \DFF_1447.CK  = CK;
  assign \DFF_1448.CK  = CK;
  assign \DFF_1449.CK  = CK;
  assign \DFF_145.CK  = CK;
  assign \DFF_1450.CK  = CK;
  assign \DFF_1451.CK  = CK;
  assign \DFF_1452.CK  = CK;
  assign \DFF_1453.CK  = CK;
  assign \DFF_1454.CK  = CK;
  assign \DFF_1455.CK  = CK;
  assign \DFF_1456.CK  = CK;
  assign \DFF_1457.CK  = CK;
  assign \DFF_1458.CK  = CK;
  assign \DFF_1459.CK  = CK;
  assign \DFF_146.CK  = CK;
  assign \DFF_1460.CK  = CK;
  assign \DFF_1461.CK  = CK;
  assign \DFF_1462.CK  = CK;
  assign \DFF_1463.CK  = CK;
  assign \DFF_1464.CK  = CK;
  assign \DFF_1465.CK  = CK;
  assign \DFF_1466.CK  = CK;
  assign \DFF_1467.CK  = CK;
  assign \DFF_1468.CK  = CK;
  assign \DFF_1469.CK  = CK;
  assign \DFF_147.CK  = CK;
  assign \DFF_1470.CK  = CK;
  assign \DFF_1471.CK  = CK;
  assign \DFF_1472.CK  = CK;
  assign \DFF_1473.CK  = CK;
  assign \DFF_1474.CK  = CK;
  assign \DFF_1475.CK  = CK;
  assign \DFF_1476.CK  = CK;
  assign \DFF_1477.CK  = CK;
  assign \DFF_1478.CK  = CK;
  assign \DFF_1479.CK  = CK;
  assign \DFF_148.CK  = CK;
  assign \DFF_1480.CK  = CK;
  assign \DFF_1481.CK  = CK;
  assign \DFF_1482.CK  = CK;
  assign \DFF_1483.CK  = CK;
  assign \DFF_1484.CK  = CK;
  assign \DFF_1485.CK  = CK;
  assign \DFF_1486.CK  = CK;
  assign \DFF_1487.CK  = CK;
  assign \DFF_1488.CK  = CK;
  assign \DFF_1489.CK  = CK;
  assign \DFF_149.CK  = CK;
  assign \DFF_1490.CK  = CK;
  assign \DFF_1491.CK  = CK;
  assign \DFF_1492.CK  = CK;
  assign \DFF_1493.CK  = CK;
  assign \DFF_1494.CK  = CK;
  assign \DFF_1495.CK  = CK;
  assign \DFF_1496.CK  = CK;
  assign \DFF_1497.CK  = CK;
  assign \DFF_1498.CK  = CK;
  assign \DFF_1499.CK  = CK;
  assign \DFF_15.CK  = CK;
  assign \DFF_150.CK  = CK;
  assign \DFF_1500.CK  = CK;
  assign \DFF_1501.CK  = CK;
  assign \DFF_1502.CK  = CK;
  assign \DFF_1503.CK  = CK;
  assign \DFF_1504.CK  = CK;
  assign \DFF_1505.CK  = CK;
  assign \DFF_1506.CK  = CK;
  assign \DFF_1507.CK  = CK;
  assign \DFF_1508.CK  = CK;
  assign \DFF_1509.CK  = CK;
  assign \DFF_151.CK  = CK;
  assign \DFF_1510.CK  = CK;
  assign \DFF_1511.CK  = CK;
  assign \DFF_1512.CK  = CK;
  assign \DFF_1513.CK  = CK;
  assign \DFF_1514.CK  = CK;
  assign \DFF_1515.CK  = CK;
  assign \DFF_1516.CK  = CK;
  assign \DFF_1517.CK  = CK;
  assign \DFF_1518.CK  = CK;
  assign \DFF_1519.CK  = CK;
  assign \DFF_152.CK  = CK;
  assign \DFF_1520.CK  = CK;
  assign \DFF_1521.CK  = CK;
  assign \DFF_1522.CK  = CK;
  assign \DFF_1523.CK  = CK;
  assign \DFF_1524.CK  = CK;
  assign \DFF_1525.CK  = CK;
  assign \DFF_1526.CK  = CK;
  assign \DFF_1527.CK  = CK;
  assign \DFF_1528.CK  = CK;
  assign \DFF_1529.CK  = CK;
  assign \DFF_153.CK  = CK;
  assign \DFF_1530.CK  = CK;
  assign \DFF_1531.CK  = CK;
  assign \DFF_1532.CK  = CK;
  assign \DFF_1533.CK  = CK;
  assign \DFF_1534.CK  = CK;
  assign \DFF_1535.CK  = CK;
  assign \DFF_1536.CK  = CK;
  assign \DFF_1537.CK  = CK;
  assign \DFF_1538.CK  = CK;
  assign \DFF_1539.CK  = CK;
  assign \DFF_154.CK  = CK;
  assign \DFF_1540.CK  = CK;
  assign \DFF_1541.CK  = CK;
  assign \DFF_1542.CK  = CK;
  assign \DFF_1543.CK  = CK;
  assign \DFF_1544.CK  = CK;
  assign \DFF_1545.CK  = CK;
  assign \DFF_1546.CK  = CK;
  assign \DFF_1547.CK  = CK;
  assign \DFF_1548.CK  = CK;
  assign \DFF_1549.CK  = CK;
  assign \DFF_155.CK  = CK;
  assign \DFF_1550.CK  = CK;
  assign \DFF_1551.CK  = CK;
  assign \DFF_1552.CK  = CK;
  assign \DFF_1553.CK  = CK;
  assign \DFF_1554.CK  = CK;
  assign \DFF_1555.CK  = CK;
  assign \DFF_1556.CK  = CK;
  assign \DFF_1557.CK  = CK;
  assign \DFF_1558.CK  = CK;
  assign \DFF_1559.CK  = CK;
  assign \DFF_156.CK  = CK;
  assign \DFF_1560.CK  = CK;
  assign \DFF_1561.CK  = CK;
  assign \DFF_1562.CK  = CK;
  assign \DFF_1563.CK  = CK;
  assign \DFF_1564.CK  = CK;
  assign \DFF_1565.CK  = CK;
  assign \DFF_1566.CK  = CK;
  assign \DFF_1567.CK  = CK;
  assign \DFF_1568.CK  = CK;
  assign \DFF_1569.CK  = CK;
  assign \DFF_157.CK  = CK;
  assign \DFF_1570.CK  = CK;
  assign \DFF_1571.CK  = CK;
  assign \DFF_1572.CK  = CK;
  assign \DFF_1573.CK  = CK;
  assign \DFF_1574.CK  = CK;
  assign \DFF_1575.CK  = CK;
  assign \DFF_1576.CK  = CK;
  assign \DFF_1577.CK  = CK;
  assign \DFF_1578.CK  = CK;
  assign \DFF_1579.CK  = CK;
  assign \DFF_158.CK  = CK;
  assign \DFF_1580.CK  = CK;
  assign \DFF_1581.CK  = CK;
  assign \DFF_1582.CK  = CK;
  assign \DFF_1583.CK  = CK;
  assign \DFF_1584.CK  = CK;
  assign \DFF_1585.CK  = CK;
  assign \DFF_1586.CK  = CK;
  assign \DFF_1587.CK  = CK;
  assign \DFF_1588.CK  = CK;
  assign \DFF_1589.CK  = CK;
  assign \DFF_159.CK  = CK;
  assign \DFF_1590.CK  = CK;
  assign \DFF_1591.CK  = CK;
  assign \DFF_1592.CK  = CK;
  assign \DFF_1593.CK  = CK;
  assign \DFF_1594.CK  = CK;
  assign \DFF_1595.CK  = CK;
  assign \DFF_1596.CK  = CK;
  assign \DFF_1597.CK  = CK;
  assign \DFF_1598.CK  = CK;
  assign \DFF_1599.CK  = CK;
  assign \DFF_16.CK  = CK;
  assign \DFF_160.CK  = CK;
  assign \DFF_1600.CK  = CK;
  assign \DFF_1601.CK  = CK;
  assign \DFF_1602.CK  = CK;
  assign \DFF_1603.CK  = CK;
  assign \DFF_1604.CK  = CK;
  assign \DFF_1605.CK  = CK;
  assign \DFF_1606.CK  = CK;
  assign \DFF_1607.CK  = CK;
  assign \DFF_1608.CK  = CK;
  assign \DFF_1609.CK  = CK;
  assign \DFF_161.CK  = CK;
  assign \DFF_1610.CK  = CK;
  assign \DFF_1611.CK  = CK;
  assign \DFF_1612.CK  = CK;
  assign \DFF_1613.CK  = CK;
  assign \DFF_1614.CK  = CK;
  assign \DFF_1615.CK  = CK;
  assign \DFF_1616.CK  = CK;
  assign \DFF_1617.CK  = CK;
  assign \DFF_1618.CK  = CK;
  assign \DFF_1619.CK  = CK;
  assign \DFF_162.CK  = CK;
  assign \DFF_1620.CK  = CK;
  assign \DFF_1621.CK  = CK;
  assign \DFF_1622.CK  = CK;
  assign \DFF_1623.CK  = CK;
  assign \DFF_1624.CK  = CK;
  assign \DFF_1625.CK  = CK;
  assign \DFF_1626.CK  = CK;
  assign \DFF_1627.CK  = CK;
  assign \DFF_1628.CK  = CK;
  assign \DFF_1629.CK  = CK;
  assign \DFF_163.CK  = CK;
  assign \DFF_1630.CK  = CK;
  assign \DFF_1631.CK  = CK;
  assign \DFF_1632.CK  = CK;
  assign \DFF_1633.CK  = CK;
  assign \DFF_1634.CK  = CK;
  assign \DFF_1635.CK  = CK;
  assign \DFF_1636.CK  = CK;
  assign \DFF_1637.CK  = CK;
  assign \DFF_1638.CK  = CK;
  assign \DFF_1639.CK  = CK;
  assign \DFF_164.CK  = CK;
  assign \DFF_1640.CK  = CK;
  assign \DFF_1641.CK  = CK;
  assign \DFF_1642.CK  = CK;
  assign \DFF_1643.CK  = CK;
  assign \DFF_1644.CK  = CK;
  assign \DFF_1645.CK  = CK;
  assign \DFF_1646.CK  = CK;
  assign \DFF_1647.CK  = CK;
  assign \DFF_1648.CK  = CK;
  assign \DFF_1649.CK  = CK;
  assign \DFF_165.CK  = CK;
  assign \DFF_1650.CK  = CK;
  assign \DFF_1651.CK  = CK;
  assign \DFF_1652.CK  = CK;
  assign \DFF_1653.CK  = CK;
  assign \DFF_1654.CK  = CK;
  assign \DFF_1655.CK  = CK;
  assign \DFF_1656.CK  = CK;
  assign \DFF_1657.CK  = CK;
  assign \DFF_1658.CK  = CK;
  assign \DFF_1659.CK  = CK;
  assign \DFF_166.CK  = CK;
  assign \DFF_1660.CK  = CK;
  assign \DFF_1661.CK  = CK;
  assign \DFF_1662.CK  = CK;
  assign \DFF_1663.CK  = CK;
  assign \DFF_1664.CK  = CK;
  assign \DFF_1665.CK  = CK;
  assign \DFF_1666.CK  = CK;
  assign \DFF_1667.CK  = CK;
  assign \DFF_1668.CK  = CK;
  assign \DFF_1669.CK  = CK;
  assign \DFF_167.CK  = CK;
  assign \DFF_1670.CK  = CK;
  assign \DFF_1671.CK  = CK;
  assign \DFF_1672.CK  = CK;
  assign \DFF_1673.CK  = CK;
  assign \DFF_1674.CK  = CK;
  assign \DFF_1675.CK  = CK;
  assign \DFF_1676.CK  = CK;
  assign \DFF_1677.CK  = CK;
  assign \DFF_1678.CK  = CK;
  assign \DFF_1679.CK  = CK;
  assign \DFF_168.CK  = CK;
  assign \DFF_1680.CK  = CK;
  assign \DFF_1681.CK  = CK;
  assign \DFF_1682.CK  = CK;
  assign \DFF_1683.CK  = CK;
  assign \DFF_1684.CK  = CK;
  assign \DFF_1685.CK  = CK;
  assign \DFF_1686.CK  = CK;
  assign \DFF_1687.CK  = CK;
  assign \DFF_1688.CK  = CK;
  assign \DFF_1689.CK  = CK;
  assign \DFF_169.CK  = CK;
  assign \DFF_1690.CK  = CK;
  assign \DFF_1691.CK  = CK;
  assign \DFF_1692.CK  = CK;
  assign \DFF_1693.CK  = CK;
  assign \DFF_1694.CK  = CK;
  assign \DFF_1695.CK  = CK;
  assign \DFF_1696.CK  = CK;
  assign \DFF_1697.CK  = CK;
  assign \DFF_1698.CK  = CK;
  assign \DFF_1699.CK  = CK;
  assign \DFF_17.CK  = CK;
  assign \DFF_170.CK  = CK;
  assign \DFF_1700.CK  = CK;
  assign \DFF_1701.CK  = CK;
  assign \DFF_1702.CK  = CK;
  assign \DFF_1703.CK  = CK;
  assign \DFF_1704.CK  = CK;
  assign \DFF_1705.CK  = CK;
  assign \DFF_1706.CK  = CK;
  assign \DFF_1707.CK  = CK;
  assign \DFF_1708.CK  = CK;
  assign \DFF_1709.CK  = CK;
  assign \DFF_171.CK  = CK;
  assign \DFF_1710.CK  = CK;
  assign \DFF_1711.CK  = CK;
  assign \DFF_1712.CK  = CK;
  assign \DFF_1713.CK  = CK;
  assign \DFF_1714.CK  = CK;
  assign \DFF_1715.CK  = CK;
  assign \DFF_1716.CK  = CK;
  assign \DFF_1717.CK  = CK;
  assign \DFF_1718.CK  = CK;
  assign \DFF_1719.CK  = CK;
  assign \DFF_172.CK  = CK;
  assign \DFF_1720.CK  = CK;
  assign \DFF_1721.CK  = CK;
  assign \DFF_1722.CK  = CK;
  assign \DFF_1723.CK  = CK;
  assign \DFF_1724.CK  = CK;
  assign \DFF_1725.CK  = CK;
  assign \DFF_1726.CK  = CK;
  assign \DFF_1727.CK  = CK;
  assign \DFF_173.CK  = CK;
  assign \DFF_174.CK  = CK;
  assign \DFF_175.CK  = CK;
  assign \DFF_176.CK  = CK;
  assign \DFF_177.CK  = CK;
  assign \DFF_178.CK  = CK;
  assign \DFF_179.CK  = CK;
  assign \DFF_18.CK  = CK;
  assign \DFF_180.CK  = CK;
  assign \DFF_181.CK  = CK;
  assign \DFF_182.CK  = CK;
  assign \DFF_183.CK  = CK;
  assign \DFF_184.CK  = CK;
  assign \DFF_185.CK  = CK;
  assign \DFF_186.CK  = CK;
  assign \DFF_187.CK  = CK;
  assign \DFF_188.CK  = CK;
  assign \DFF_189.CK  = CK;
  assign \DFF_19.CK  = CK;
  assign \DFF_190.CK  = CK;
  assign \DFF_191.CK  = CK;
  assign \DFF_192.CK  = CK;
  assign \DFF_193.CK  = CK;
  assign \DFF_194.CK  = CK;
  assign \DFF_195.CK  = CK;
  assign \DFF_196.CK  = CK;
  assign \DFF_197.CK  = CK;
  assign \DFF_198.CK  = CK;
  assign \DFF_199.CK  = CK;
  assign \DFF_2.CK  = CK;
  assign \DFF_20.CK  = CK;
  assign \DFF_200.CK  = CK;
  assign \DFF_201.CK  = CK;
  assign \DFF_202.CK  = CK;
  assign \DFF_203.CK  = CK;
  assign \DFF_204.CK  = CK;
  assign \DFF_205.CK  = CK;
  assign \DFF_206.CK  = CK;
  assign \DFF_207.CK  = CK;
  assign \DFF_208.CK  = CK;
  assign \DFF_209.CK  = CK;
  assign \DFF_21.CK  = CK;
  assign \DFF_210.CK  = CK;
  assign \DFF_211.CK  = CK;
  assign \DFF_212.CK  = CK;
  assign \DFF_213.CK  = CK;
  assign \DFF_214.CK  = CK;
  assign \DFF_215.CK  = CK;
  assign \DFF_216.CK  = CK;
  assign \DFF_217.CK  = CK;
  assign \DFF_218.CK  = CK;
  assign \DFF_219.CK  = CK;
  assign \DFF_22.CK  = CK;
  assign \DFF_220.CK  = CK;
  assign \DFF_221.CK  = CK;
  assign \DFF_222.CK  = CK;
  assign \DFF_223.CK  = CK;
  assign \DFF_224.CK  = CK;
  assign \DFF_225.CK  = CK;
  assign \DFF_226.CK  = CK;
  assign \DFF_227.CK  = CK;
  assign \DFF_228.CK  = CK;
  assign \DFF_229.CK  = CK;
  assign \DFF_23.CK  = CK;
  assign \DFF_230.CK  = CK;
  assign \DFF_231.CK  = CK;
  assign \DFF_232.CK  = CK;
  assign \DFF_233.CK  = CK;
  assign \DFF_234.CK  = CK;
  assign \DFF_235.CK  = CK;
  assign \DFF_236.CK  = CK;
  assign \DFF_237.CK  = CK;
  assign \DFF_238.CK  = CK;
  assign \DFF_239.CK  = CK;
  assign \DFF_24.CK  = CK;
  assign \DFF_240.CK  = CK;
  assign \DFF_241.CK  = CK;
  assign \DFF_242.CK  = CK;
  assign \DFF_243.CK  = CK;
  assign \DFF_244.CK  = CK;
  assign \DFF_245.CK  = CK;
  assign \DFF_246.CK  = CK;
  assign \DFF_247.CK  = CK;
  assign \DFF_248.CK  = CK;
  assign \DFF_249.CK  = CK;
  assign \DFF_25.CK  = CK;
  assign \DFF_250.CK  = CK;
  assign \DFF_251.CK  = CK;
  assign \DFF_252.CK  = CK;
  assign \DFF_253.CK  = CK;
  assign \DFF_254.CK  = CK;
  assign \DFF_255.CK  = CK;
  assign \DFF_256.CK  = CK;
  assign \DFF_257.CK  = CK;
  assign \DFF_258.CK  = CK;
  assign \DFF_259.CK  = CK;
  assign \DFF_26.CK  = CK;
  assign \DFF_260.CK  = CK;
  assign \DFF_261.CK  = CK;
  assign \DFF_262.CK  = CK;
  assign \DFF_263.CK  = CK;
  assign \DFF_264.CK  = CK;
  assign \DFF_265.CK  = CK;
  assign \DFF_266.CK  = CK;
  assign \DFF_267.CK  = CK;
  assign \DFF_268.CK  = CK;
  assign \DFF_269.CK  = CK;
  assign \DFF_27.CK  = CK;
  assign \DFF_270.CK  = CK;
  assign \DFF_271.CK  = CK;
  assign \DFF_272.CK  = CK;
  assign \DFF_273.CK  = CK;
  assign \DFF_274.CK  = CK;
  assign \DFF_275.CK  = CK;
  assign \DFF_276.CK  = CK;
  assign \DFF_277.CK  = CK;
  assign \DFF_278.CK  = CK;
  assign \DFF_279.CK  = CK;
  assign \DFF_28.CK  = CK;
  assign \DFF_280.CK  = CK;
  assign \DFF_281.CK  = CK;
  assign \DFF_282.CK  = CK;
  assign \DFF_283.CK  = CK;
  assign \DFF_284.CK  = CK;
  assign \DFF_285.CK  = CK;
  assign \DFF_286.CK  = CK;
  assign \DFF_287.CK  = CK;
  assign \DFF_288.CK  = CK;
  assign \DFF_289.CK  = CK;
  assign \DFF_29.CK  = CK;
  assign \DFF_290.CK  = CK;
  assign \DFF_291.CK  = CK;
  assign \DFF_292.CK  = CK;
  assign \DFF_293.CK  = CK;
  assign \DFF_294.CK  = CK;
  assign \DFF_295.CK  = CK;
  assign \DFF_296.CK  = CK;
  assign \DFF_297.CK  = CK;
  assign \DFF_298.CK  = CK;
  assign \DFF_299.CK  = CK;
  assign \DFF_3.CK  = CK;
  assign \DFF_30.CK  = CK;
  assign \DFF_300.CK  = CK;
  assign \DFF_301.CK  = CK;
  assign \DFF_302.CK  = CK;
  assign \DFF_303.CK  = CK;
  assign \DFF_304.CK  = CK;
  assign \DFF_305.CK  = CK;
  assign \DFF_306.CK  = CK;
  assign \DFF_307.CK  = CK;
  assign \DFF_308.CK  = CK;
  assign \DFF_309.CK  = CK;
  assign \DFF_31.CK  = CK;
  assign \DFF_310.CK  = CK;
  assign \DFF_311.CK  = CK;
  assign \DFF_312.CK  = CK;
  assign \DFF_313.CK  = CK;
  assign \DFF_314.CK  = CK;
  assign \DFF_315.CK  = CK;
  assign \DFF_316.CK  = CK;
  assign \DFF_317.CK  = CK;
  assign \DFF_318.CK  = CK;
  assign \DFF_319.CK  = CK;
  assign \DFF_32.CK  = CK;
  assign \DFF_320.CK  = CK;
  assign \DFF_321.CK  = CK;
  assign \DFF_322.CK  = CK;
  assign \DFF_323.CK  = CK;
  assign \DFF_324.CK  = CK;
  assign \DFF_325.CK  = CK;
  assign \DFF_326.CK  = CK;
  assign \DFF_327.CK  = CK;
  assign \DFF_328.CK  = CK;
  assign \DFF_329.CK  = CK;
  assign \DFF_33.CK  = CK;
  assign \DFF_330.CK  = CK;
  assign \DFF_331.CK  = CK;
  assign \DFF_332.CK  = CK;
  assign \DFF_333.CK  = CK;
  assign \DFF_334.CK  = CK;
  assign \DFF_335.CK  = CK;
  assign \DFF_336.CK  = CK;
  assign \DFF_337.CK  = CK;
  assign \DFF_338.CK  = CK;
  assign \DFF_339.CK  = CK;
  assign \DFF_34.CK  = CK;
  assign \DFF_340.CK  = CK;
  assign \DFF_341.CK  = CK;
  assign \DFF_342.CK  = CK;
  assign \DFF_343.CK  = CK;
  assign \DFF_344.CK  = CK;
  assign \DFF_345.CK  = CK;
  assign \DFF_346.CK  = CK;
  assign \DFF_347.CK  = CK;
  assign \DFF_348.CK  = CK;
  assign \DFF_349.CK  = CK;
  assign \DFF_35.CK  = CK;
  assign \DFF_350.CK  = CK;
  assign \DFF_351.CK  = CK;
  assign \DFF_352.CK  = CK;
  assign \DFF_353.CK  = CK;
  assign \DFF_354.CK  = CK;
  assign \DFF_355.CK  = CK;
  assign \DFF_356.CK  = CK;
  assign \DFF_357.CK  = CK;
  assign \DFF_358.CK  = CK;
  assign \DFF_359.CK  = CK;
  assign \DFF_36.CK  = CK;
  assign \DFF_360.CK  = CK;
  assign \DFF_361.CK  = CK;
  assign \DFF_362.CK  = CK;
  assign \DFF_363.CK  = CK;
  assign \DFF_364.CK  = CK;
  assign \DFF_365.CK  = CK;
  assign \DFF_366.CK  = CK;
  assign \DFF_367.CK  = CK;
  assign \DFF_368.CK  = CK;
  assign \DFF_369.CK  = CK;
  assign \DFF_37.CK  = CK;
  assign \DFF_370.CK  = CK;
  assign \DFF_371.CK  = CK;
  assign \DFF_372.CK  = CK;
  assign \DFF_373.CK  = CK;
  assign \DFF_374.CK  = CK;
  assign \DFF_375.CK  = CK;
  assign \DFF_376.CK  = CK;
  assign \DFF_377.CK  = CK;
  assign \DFF_378.CK  = CK;
  assign \DFF_379.CK  = CK;
  assign \DFF_38.CK  = CK;
  assign \DFF_380.CK  = CK;
  assign \DFF_381.CK  = CK;
  assign \DFF_382.CK  = CK;
  assign \DFF_383.CK  = CK;
  assign \DFF_384.CK  = CK;
  assign \DFF_385.CK  = CK;
  assign \DFF_386.CK  = CK;
  assign \DFF_387.CK  = CK;
  assign \DFF_388.CK  = CK;
  assign \DFF_389.CK  = CK;
  assign \DFF_39.CK  = CK;
  assign \DFF_390.CK  = CK;
  assign \DFF_391.CK  = CK;
  assign \DFF_392.CK  = CK;
  assign \DFF_393.CK  = CK;
  assign \DFF_394.CK  = CK;
  assign \DFF_395.CK  = CK;
  assign \DFF_396.CK  = CK;
  assign \DFF_397.CK  = CK;
  assign \DFF_398.CK  = CK;
  assign \DFF_399.CK  = CK;
  assign \DFF_4.CK  = CK;
  assign \DFF_40.CK  = CK;
  assign \DFF_400.CK  = CK;
  assign \DFF_401.CK  = CK;
  assign \DFF_402.CK  = CK;
  assign \DFF_403.CK  = CK;
  assign \DFF_404.CK  = CK;
  assign \DFF_405.CK  = CK;
  assign \DFF_406.CK  = CK;
  assign \DFF_407.CK  = CK;
  assign \DFF_408.CK  = CK;
  assign \DFF_409.CK  = CK;
  assign \DFF_41.CK  = CK;
  assign \DFF_410.CK  = CK;
  assign \DFF_411.CK  = CK;
  assign \DFF_412.CK  = CK;
  assign \DFF_413.CK  = CK;
  assign \DFF_414.CK  = CK;
  assign \DFF_415.CK  = CK;
  assign \DFF_416.CK  = CK;
  assign \DFF_417.CK  = CK;
  assign \DFF_418.CK  = CK;
  assign \DFF_419.CK  = CK;
  assign \DFF_42.CK  = CK;
  assign \DFF_420.CK  = CK;
  assign \DFF_421.CK  = CK;
  assign \DFF_422.CK  = CK;
  assign \DFF_423.CK  = CK;
  assign \DFF_424.CK  = CK;
  assign \DFF_425.CK  = CK;
  assign \DFF_426.CK  = CK;
  assign \DFF_427.CK  = CK;
  assign \DFF_428.CK  = CK;
  assign \DFF_429.CK  = CK;
  assign \DFF_43.CK  = CK;
  assign \DFF_430.CK  = CK;
  assign \DFF_431.CK  = CK;
  assign \DFF_432.CK  = CK;
  assign \DFF_433.CK  = CK;
  assign \DFF_434.CK  = CK;
  assign \DFF_435.CK  = CK;
  assign \DFF_436.CK  = CK;
  assign \DFF_437.CK  = CK;
  assign \DFF_438.CK  = CK;
  assign \DFF_439.CK  = CK;
  assign \DFF_44.CK  = CK;
  assign \DFF_440.CK  = CK;
  assign \DFF_441.CK  = CK;
  assign \DFF_442.CK  = CK;
  assign \DFF_443.CK  = CK;
  assign \DFF_444.CK  = CK;
  assign \DFF_445.CK  = CK;
  assign \DFF_446.CK  = CK;
  assign \DFF_447.CK  = CK;
  assign \DFF_448.CK  = CK;
  assign \DFF_449.CK  = CK;
  assign \DFF_45.CK  = CK;
  assign \DFF_450.CK  = CK;
  assign \DFF_451.CK  = CK;
  assign \DFF_452.CK  = CK;
  assign \DFF_453.CK  = CK;
  assign \DFF_454.CK  = CK;
  assign \DFF_455.CK  = CK;
  assign \DFF_456.CK  = CK;
  assign \DFF_457.CK  = CK;
  assign \DFF_458.CK  = CK;
  assign \DFF_459.CK  = CK;
  assign \DFF_46.CK  = CK;
  assign \DFF_460.CK  = CK;
  assign \DFF_461.CK  = CK;
  assign \DFF_462.CK  = CK;
  assign \DFF_463.CK  = CK;
  assign \DFF_464.CK  = CK;
  assign \DFF_465.CK  = CK;
  assign \DFF_466.CK  = CK;
  assign \DFF_467.CK  = CK;
  assign \DFF_468.CK  = CK;
  assign \DFF_469.CK  = CK;
  assign \DFF_47.CK  = CK;
  assign \DFF_470.CK  = CK;
  assign \DFF_471.CK  = CK;
  assign \DFF_472.CK  = CK;
  assign \DFF_473.CK  = CK;
  assign \DFF_474.CK  = CK;
  assign \DFF_475.CK  = CK;
  assign \DFF_476.CK  = CK;
  assign \DFF_477.CK  = CK;
  assign \DFF_478.CK  = CK;
  assign \DFF_479.CK  = CK;
  assign \DFF_48.CK  = CK;
  assign \DFF_480.CK  = CK;
  assign \DFF_481.CK  = CK;
  assign \DFF_482.CK  = CK;
  assign \DFF_483.CK  = CK;
  assign \DFF_484.CK  = CK;
  assign \DFF_485.CK  = CK;
  assign \DFF_486.CK  = CK;
  assign \DFF_487.CK  = CK;
  assign \DFF_488.CK  = CK;
  assign \DFF_489.CK  = CK;
  assign \DFF_49.CK  = CK;
  assign \DFF_490.CK  = CK;
  assign \DFF_491.CK  = CK;
  assign \DFF_492.CK  = CK;
  assign \DFF_493.CK  = CK;
  assign \DFF_494.CK  = CK;
  assign \DFF_495.CK  = CK;
  assign \DFF_496.CK  = CK;
  assign \DFF_497.CK  = CK;
  assign \DFF_498.CK  = CK;
  assign \DFF_499.CK  = CK;
  assign \DFF_5.CK  = CK;
  assign \DFF_50.CK  = CK;
  assign \DFF_500.CK  = CK;
  assign \DFF_501.CK  = CK;
  assign \DFF_502.CK  = CK;
  assign \DFF_503.CK  = CK;
  assign \DFF_504.CK  = CK;
  assign \DFF_505.CK  = CK;
  assign \DFF_506.CK  = CK;
  assign \DFF_507.CK  = CK;
  assign \DFF_508.CK  = CK;
  assign \DFF_509.CK  = CK;
  assign \DFF_51.CK  = CK;
  assign \DFF_510.CK  = CK;
  assign \DFF_511.CK  = CK;
  assign \DFF_512.CK  = CK;
  assign \DFF_513.CK  = CK;
  assign \DFF_514.CK  = CK;
  assign \DFF_515.CK  = CK;
  assign \DFF_516.CK  = CK;
  assign \DFF_517.CK  = CK;
  assign \DFF_518.CK  = CK;
  assign \DFF_519.CK  = CK;
  assign \DFF_52.CK  = CK;
  assign \DFF_520.CK  = CK;
  assign \DFF_521.CK  = CK;
  assign \DFF_522.CK  = CK;
  assign \DFF_523.CK  = CK;
  assign \DFF_524.CK  = CK;
  assign \DFF_525.CK  = CK;
  assign \DFF_526.CK  = CK;
  assign \DFF_527.CK  = CK;
  assign \DFF_528.CK  = CK;
  assign \DFF_529.CK  = CK;
  assign \DFF_53.CK  = CK;
  assign \DFF_530.CK  = CK;
  assign \DFF_531.CK  = CK;
  assign \DFF_532.CK  = CK;
  assign \DFF_533.CK  = CK;
  assign \DFF_534.CK  = CK;
  assign \DFF_535.CK  = CK;
  assign \DFF_536.CK  = CK;
  assign \DFF_537.CK  = CK;
  assign \DFF_538.CK  = CK;
  assign \DFF_539.CK  = CK;
  assign \DFF_54.CK  = CK;
  assign \DFF_540.CK  = CK;
  assign \DFF_541.CK  = CK;
  assign \DFF_542.CK  = CK;
  assign \DFF_543.CK  = CK;
  assign \DFF_544.CK  = CK;
  assign \DFF_545.CK  = CK;
  assign \DFF_546.CK  = CK;
  assign \DFF_547.CK  = CK;
  assign \DFF_548.CK  = CK;
  assign \DFF_549.CK  = CK;
  assign \DFF_55.CK  = CK;
  assign \DFF_550.CK  = CK;
  assign \DFF_551.CK  = CK;
  assign \DFF_552.CK  = CK;
  assign \DFF_553.CK  = CK;
  assign \DFF_554.CK  = CK;
  assign \DFF_555.CK  = CK;
  assign \DFF_556.CK  = CK;
  assign \DFF_557.CK  = CK;
  assign \DFF_558.CK  = CK;
  assign \DFF_559.CK  = CK;
  assign \DFF_56.CK  = CK;
  assign \DFF_560.CK  = CK;
  assign \DFF_561.CK  = CK;
  assign \DFF_562.CK  = CK;
  assign \DFF_563.CK  = CK;
  assign \DFF_564.CK  = CK;
  assign \DFF_565.CK  = CK;
  assign \DFF_566.CK  = CK;
  assign \DFF_567.CK  = CK;
  assign \DFF_568.CK  = CK;
  assign \DFF_569.CK  = CK;
  assign \DFF_57.CK  = CK;
  assign \DFF_570.CK  = CK;
  assign \DFF_571.CK  = CK;
  assign \DFF_572.CK  = CK;
  assign \DFF_573.CK  = CK;
  assign \DFF_574.CK  = CK;
  assign \DFF_575.CK  = CK;
  assign \DFF_576.CK  = CK;
  assign \DFF_577.CK  = CK;
  assign \DFF_578.CK  = CK;
  assign \DFF_579.CK  = CK;
  assign \DFF_58.CK  = CK;
  assign \DFF_580.CK  = CK;
  assign \DFF_581.CK  = CK;
  assign \DFF_582.CK  = CK;
  assign \DFF_583.CK  = CK;
  assign \DFF_584.CK  = CK;
  assign \DFF_585.CK  = CK;
  assign \DFF_586.CK  = CK;
  assign \DFF_587.CK  = CK;
  assign \DFF_588.CK  = CK;
  assign \DFF_589.CK  = CK;
  assign \DFF_59.CK  = CK;
  assign \DFF_590.CK  = CK;
  assign \DFF_591.CK  = CK;
  assign \DFF_592.CK  = CK;
  assign \DFF_593.CK  = CK;
  assign \DFF_594.CK  = CK;
  assign \DFF_595.CK  = CK;
  assign \DFF_596.CK  = CK;
  assign \DFF_597.CK  = CK;
  assign \DFF_598.CK  = CK;
  assign \DFF_599.CK  = CK;
  assign \DFF_6.CK  = CK;
  assign \DFF_60.CK  = CK;
  assign \DFF_600.CK  = CK;
  assign \DFF_601.CK  = CK;
  assign \DFF_602.CK  = CK;
  assign \DFF_603.CK  = CK;
  assign \DFF_604.CK  = CK;
  assign \DFF_605.CK  = CK;
  assign \DFF_606.CK  = CK;
  assign \DFF_607.CK  = CK;
  assign \DFF_608.CK  = CK;
  assign \DFF_609.CK  = CK;
  assign \DFF_61.CK  = CK;
  assign \DFF_610.CK  = CK;
  assign \DFF_611.CK  = CK;
  assign \DFF_612.CK  = CK;
  assign \DFF_613.CK  = CK;
  assign \DFF_614.CK  = CK;
  assign \DFF_615.CK  = CK;
  assign \DFF_616.CK  = CK;
  assign \DFF_617.CK  = CK;
  assign \DFF_618.CK  = CK;
  assign \DFF_619.CK  = CK;
  assign \DFF_62.CK  = CK;
  assign \DFF_620.CK  = CK;
  assign \DFF_621.CK  = CK;
  assign \DFF_622.CK  = CK;
  assign \DFF_623.CK  = CK;
  assign \DFF_624.CK  = CK;
  assign \DFF_625.CK  = CK;
  assign \DFF_626.CK  = CK;
  assign \DFF_627.CK  = CK;
  assign \DFF_628.CK  = CK;
  assign \DFF_629.CK  = CK;
  assign \DFF_63.CK  = CK;
  assign \DFF_630.CK  = CK;
  assign \DFF_631.CK  = CK;
  assign \DFF_632.CK  = CK;
  assign \DFF_633.CK  = CK;
  assign \DFF_634.CK  = CK;
  assign \DFF_635.CK  = CK;
  assign \DFF_636.CK  = CK;
  assign \DFF_637.CK  = CK;
  assign \DFF_638.CK  = CK;
  assign \DFF_639.CK  = CK;
  assign \DFF_64.CK  = CK;
  assign \DFF_640.CK  = CK;
  assign \DFF_641.CK  = CK;
  assign \DFF_642.CK  = CK;
  assign \DFF_643.CK  = CK;
  assign \DFF_644.CK  = CK;
  assign \DFF_645.CK  = CK;
  assign \DFF_646.CK  = CK;
  assign \DFF_647.CK  = CK;
  assign \DFF_648.CK  = CK;
  assign \DFF_649.CK  = CK;
  assign \DFF_65.CK  = CK;
  assign \DFF_650.CK  = CK;
  assign \DFF_651.CK  = CK;
  assign \DFF_652.CK  = CK;
  assign \DFF_653.CK  = CK;
  assign \DFF_654.CK  = CK;
  assign \DFF_655.CK  = CK;
  assign \DFF_656.CK  = CK;
  assign \DFF_657.CK  = CK;
  assign \DFF_658.CK  = CK;
  assign \DFF_659.CK  = CK;
  assign \DFF_66.CK  = CK;
  assign \DFF_660.CK  = CK;
  assign \DFF_661.CK  = CK;
  assign \DFF_662.CK  = CK;
  assign \DFF_663.CK  = CK;
  assign \DFF_664.CK  = CK;
  assign \DFF_665.CK  = CK;
  assign \DFF_666.CK  = CK;
  assign \DFF_667.CK  = CK;
  assign \DFF_668.CK  = CK;
  assign \DFF_669.CK  = CK;
  assign \DFF_67.CK  = CK;
  assign \DFF_670.CK  = CK;
  assign \DFF_671.CK  = CK;
  assign \DFF_672.CK  = CK;
  assign \DFF_673.CK  = CK;
  assign \DFF_674.CK  = CK;
  assign \DFF_675.CK  = CK;
  assign \DFF_676.CK  = CK;
  assign \DFF_677.CK  = CK;
  assign \DFF_678.CK  = CK;
  assign \DFF_679.CK  = CK;
  assign \DFF_68.CK  = CK;
  assign \DFF_680.CK  = CK;
  assign \DFF_681.CK  = CK;
  assign \DFF_682.CK  = CK;
  assign \DFF_683.CK  = CK;
  assign \DFF_684.CK  = CK;
  assign \DFF_685.CK  = CK;
  assign \DFF_686.CK  = CK;
  assign \DFF_687.CK  = CK;
  assign \DFF_688.CK  = CK;
  assign \DFF_689.CK  = CK;
  assign \DFF_69.CK  = CK;
  assign \DFF_690.CK  = CK;
  assign \DFF_691.CK  = CK;
  assign \DFF_692.CK  = CK;
  assign \DFF_693.CK  = CK;
  assign \DFF_694.CK  = CK;
  assign \DFF_695.CK  = CK;
  assign \DFF_696.CK  = CK;
  assign \DFF_697.CK  = CK;
  assign \DFF_698.CK  = CK;
  assign \DFF_699.CK  = CK;
  assign \DFF_7.CK  = CK;
  assign \DFF_70.CK  = CK;
  assign \DFF_700.CK  = CK;
  assign \DFF_701.CK  = CK;
  assign \DFF_702.CK  = CK;
  assign \DFF_703.CK  = CK;
  assign \DFF_704.CK  = CK;
  assign \DFF_705.CK  = CK;
  assign \DFF_706.CK  = CK;
  assign \DFF_707.CK  = CK;
  assign \DFF_708.CK  = CK;
  assign \DFF_709.CK  = CK;
  assign \DFF_71.CK  = CK;
  assign \DFF_710.CK  = CK;
  assign \DFF_711.CK  = CK;
  assign \DFF_712.CK  = CK;
  assign \DFF_713.CK  = CK;
  assign \DFF_714.CK  = CK;
  assign \DFF_715.CK  = CK;
  assign \DFF_716.CK  = CK;
  assign \DFF_717.CK  = CK;
  assign \DFF_718.CK  = CK;
  assign \DFF_719.CK  = CK;
  assign \DFF_72.CK  = CK;
  assign \DFF_720.CK  = CK;
  assign \DFF_721.CK  = CK;
  assign \DFF_722.CK  = CK;
  assign \DFF_723.CK  = CK;
  assign \DFF_724.CK  = CK;
  assign \DFF_725.CK  = CK;
  assign \DFF_726.CK  = CK;
  assign \DFF_727.CK  = CK;
  assign \DFF_728.CK  = CK;
  assign \DFF_729.CK  = CK;
  assign \DFF_73.CK  = CK;
  assign \DFF_730.CK  = CK;
  assign \DFF_731.CK  = CK;
  assign \DFF_732.CK  = CK;
  assign \DFF_733.CK  = CK;
  assign \DFF_734.CK  = CK;
  assign \DFF_735.CK  = CK;
  assign \DFF_736.CK  = CK;
  assign \DFF_737.CK  = CK;
  assign \DFF_738.CK  = CK;
  assign \DFF_739.CK  = CK;
  assign \DFF_74.CK  = CK;
  assign \DFF_740.CK  = CK;
  assign \DFF_741.CK  = CK;
  assign \DFF_742.CK  = CK;
  assign \DFF_743.CK  = CK;
  assign \DFF_744.CK  = CK;
  assign \DFF_745.CK  = CK;
  assign \DFF_746.CK  = CK;
  assign \DFF_747.CK  = CK;
  assign \DFF_748.CK  = CK;
  assign \DFF_749.CK  = CK;
  assign \DFF_75.CK  = CK;
  assign \DFF_750.CK  = CK;
  assign \DFF_751.CK  = CK;
  assign \DFF_752.CK  = CK;
  assign \DFF_753.CK  = CK;
  assign \DFF_754.CK  = CK;
  assign \DFF_755.CK  = CK;
  assign \DFF_756.CK  = CK;
  assign \DFF_757.CK  = CK;
  assign \DFF_758.CK  = CK;
  assign \DFF_759.CK  = CK;
  assign \DFF_76.CK  = CK;
  assign \DFF_760.CK  = CK;
  assign \DFF_761.CK  = CK;
  assign \DFF_762.CK  = CK;
  assign \DFF_763.CK  = CK;
  assign \DFF_764.CK  = CK;
  assign \DFF_765.CK  = CK;
  assign \DFF_766.CK  = CK;
  assign \DFF_767.CK  = CK;
  assign \DFF_768.CK  = CK;
  assign \DFF_769.CK  = CK;
  assign \DFF_77.CK  = CK;
  assign \DFF_770.CK  = CK;
  assign \DFF_771.CK  = CK;
  assign \DFF_772.CK  = CK;
  assign \DFF_773.CK  = CK;
  assign \DFF_774.CK  = CK;
  assign \DFF_775.CK  = CK;
  assign \DFF_776.CK  = CK;
  assign \DFF_777.CK  = CK;
  assign \DFF_778.CK  = CK;
  assign \DFF_779.CK  = CK;
  assign \DFF_78.CK  = CK;
  assign \DFF_780.CK  = CK;
  assign \DFF_781.CK  = CK;
  assign \DFF_782.CK  = CK;
  assign \DFF_783.CK  = CK;
  assign \DFF_784.CK  = CK;
  assign \DFF_785.CK  = CK;
  assign \DFF_786.CK  = CK;
  assign \DFF_787.CK  = CK;
  assign \DFF_788.CK  = CK;
  assign \DFF_789.CK  = CK;
  assign \DFF_79.CK  = CK;
  assign \DFF_790.CK  = CK;
  assign \DFF_791.CK  = CK;
  assign \DFF_792.CK  = CK;
  assign \DFF_793.CK  = CK;
  assign \DFF_794.CK  = CK;
  assign \DFF_795.CK  = CK;
  assign \DFF_796.CK  = CK;
  assign \DFF_797.CK  = CK;
  assign \DFF_798.CK  = CK;
  assign \DFF_799.CK  = CK;
  assign \DFF_8.CK  = CK;
  assign \DFF_80.CK  = CK;
  assign \DFF_800.CK  = CK;
  assign \DFF_801.CK  = CK;
  assign \DFF_802.CK  = CK;
  assign \DFF_803.CK  = CK;
  assign \DFF_804.CK  = CK;
  assign \DFF_805.CK  = CK;
  assign \DFF_806.CK  = CK;
  assign \DFF_807.CK  = CK;
  assign \DFF_808.CK  = CK;
  assign \DFF_809.CK  = CK;
  assign \DFF_81.CK  = CK;
  assign \DFF_810.CK  = CK;
  assign \DFF_811.CK  = CK;
  assign \DFF_812.CK  = CK;
  assign \DFF_813.CK  = CK;
  assign \DFF_814.CK  = CK;
  assign \DFF_815.CK  = CK;
  assign \DFF_816.CK  = CK;
  assign \DFF_817.CK  = CK;
  assign \DFF_818.CK  = CK;
  assign \DFF_819.CK  = CK;
  assign \DFF_82.CK  = CK;
  assign \DFF_820.CK  = CK;
  assign \DFF_821.CK  = CK;
  assign \DFF_822.CK  = CK;
  assign \DFF_823.CK  = CK;
  assign \DFF_824.CK  = CK;
  assign \DFF_825.CK  = CK;
  assign \DFF_826.CK  = CK;
  assign \DFF_827.CK  = CK;
  assign \DFF_828.CK  = CK;
  assign \DFF_829.CK  = CK;
  assign \DFF_83.CK  = CK;
  assign \DFF_830.CK  = CK;
  assign \DFF_831.CK  = CK;
  assign \DFF_832.CK  = CK;
  assign \DFF_833.CK  = CK;
  assign \DFF_834.CK  = CK;
  assign \DFF_835.CK  = CK;
  assign \DFF_836.CK  = CK;
  assign \DFF_837.CK  = CK;
  assign \DFF_838.CK  = CK;
  assign \DFF_839.CK  = CK;
  assign \DFF_84.CK  = CK;
  assign \DFF_840.CK  = CK;
  assign \DFF_841.CK  = CK;
  assign \DFF_842.CK  = CK;
  assign \DFF_843.CK  = CK;
  assign \DFF_844.CK  = CK;
  assign \DFF_845.CK  = CK;
  assign \DFF_846.CK  = CK;
  assign \DFF_847.CK  = CK;
  assign \DFF_848.CK  = CK;
  assign \DFF_849.CK  = CK;
  assign \DFF_85.CK  = CK;
  assign \DFF_850.CK  = CK;
  assign \DFF_851.CK  = CK;
  assign \DFF_852.CK  = CK;
  assign \DFF_853.CK  = CK;
  assign \DFF_854.CK  = CK;
  assign \DFF_855.CK  = CK;
  assign \DFF_856.CK  = CK;
  assign \DFF_857.CK  = CK;
  assign \DFF_858.CK  = CK;
  assign \DFF_859.CK  = CK;
  assign \DFF_86.CK  = CK;
  assign \DFF_860.CK  = CK;
  assign \DFF_861.CK  = CK;
  assign \DFF_862.CK  = CK;
  assign \DFF_863.CK  = CK;
  assign \DFF_864.CK  = CK;
  assign \DFF_865.CK  = CK;
  assign \DFF_866.CK  = CK;
  assign \DFF_867.CK  = CK;
  assign \DFF_868.CK  = CK;
  assign \DFF_869.CK  = CK;
  assign \DFF_87.CK  = CK;
  assign \DFF_870.CK  = CK;
  assign \DFF_871.CK  = CK;
  assign \DFF_872.CK  = CK;
  assign \DFF_873.CK  = CK;
  assign \DFF_874.CK  = CK;
  assign \DFF_875.CK  = CK;
  assign \DFF_876.CK  = CK;
  assign \DFF_877.CK  = CK;
  assign \DFF_878.CK  = CK;
  assign \DFF_879.CK  = CK;
  assign \DFF_88.CK  = CK;
  assign \DFF_880.CK  = CK;
  assign \DFF_881.CK  = CK;
  assign \DFF_882.CK  = CK;
  assign \DFF_883.CK  = CK;
  assign \DFF_884.CK  = CK;
  assign \DFF_885.CK  = CK;
  assign \DFF_886.CK  = CK;
  assign \DFF_887.CK  = CK;
  assign \DFF_888.CK  = CK;
  assign \DFF_889.CK  = CK;
  assign \DFF_89.CK  = CK;
  assign \DFF_890.CK  = CK;
  assign \DFF_891.CK  = CK;
  assign \DFF_892.CK  = CK;
  assign \DFF_893.CK  = CK;
  assign \DFF_894.CK  = CK;
  assign \DFF_895.CK  = CK;
  assign \DFF_896.CK  = CK;
  assign \DFF_897.CK  = CK;
  assign \DFF_898.CK  = CK;
  assign \DFF_899.CK  = CK;
  assign \DFF_9.CK  = CK;
  assign \DFF_90.CK  = CK;
  assign \DFF_900.CK  = CK;
  assign \DFF_901.CK  = CK;
  assign \DFF_902.CK  = CK;
  assign \DFF_903.CK  = CK;
  assign \DFF_904.CK  = CK;
  assign \DFF_905.CK  = CK;
  assign \DFF_906.CK  = CK;
  assign \DFF_907.CK  = CK;
  assign \DFF_908.CK  = CK;
  assign \DFF_909.CK  = CK;
  assign \DFF_91.CK  = CK;
  assign \DFF_910.CK  = CK;
  assign \DFF_911.CK  = CK;
  assign \DFF_912.CK  = CK;
  assign \DFF_913.CK  = CK;
  assign \DFF_914.CK  = CK;
  assign \DFF_915.CK  = CK;
  assign \DFF_916.CK  = CK;
  assign \DFF_917.CK  = CK;
  assign \DFF_918.CK  = CK;
  assign \DFF_919.CK  = CK;
  assign \DFF_92.CK  = CK;
  assign \DFF_920.CK  = CK;
  assign \DFF_921.CK  = CK;
  assign \DFF_922.CK  = CK;
  assign \DFF_923.CK  = CK;
  assign \DFF_924.CK  = CK;
  assign \DFF_925.CK  = CK;
  assign \DFF_926.CK  = CK;
  assign \DFF_927.CK  = CK;
  assign \DFF_928.CK  = CK;
  assign \DFF_929.CK  = CK;
  assign \DFF_93.CK  = CK;
  assign \DFF_930.CK  = CK;
  assign \DFF_931.CK  = CK;
  assign \DFF_932.CK  = CK;
  assign \DFF_933.CK  = CK;
  assign \DFF_934.CK  = CK;
  assign \DFF_935.CK  = CK;
  assign \DFF_936.CK  = CK;
  assign \DFF_937.CK  = CK;
  assign \DFF_938.CK  = CK;
  assign \DFF_939.CK  = CK;
  assign \DFF_94.CK  = CK;
  assign \DFF_940.CK  = CK;
  assign \DFF_941.CK  = CK;
  assign \DFF_942.CK  = CK;
  assign \DFF_943.CK  = CK;
  assign \DFF_944.CK  = CK;
  assign \DFF_945.CK  = CK;
  assign \DFF_946.CK  = CK;
  assign \DFF_947.CK  = CK;
  assign \DFF_948.CK  = CK;
  assign \DFF_949.CK  = CK;
  assign \DFF_95.CK  = CK;
  assign \DFF_950.CK  = CK;
  assign \DFF_951.CK  = CK;
  assign \DFF_952.CK  = CK;
  assign \DFF_953.CK  = CK;
  assign \DFF_954.CK  = CK;
  assign \DFF_955.CK  = CK;
  assign \DFF_956.CK  = CK;
  assign \DFF_957.CK  = CK;
  assign \DFF_958.CK  = CK;
  assign \DFF_959.CK  = CK;
  assign \DFF_96.CK  = CK;
  assign \DFF_960.CK  = CK;
  assign \DFF_961.CK  = CK;
  assign \DFF_962.CK  = CK;
  assign \DFF_963.CK  = CK;
  assign \DFF_964.CK  = CK;
  assign \DFF_965.CK  = CK;
  assign \DFF_966.CK  = CK;
  assign \DFF_967.CK  = CK;
  assign \DFF_968.CK  = CK;
  assign \DFF_969.CK  = CK;
  assign \DFF_97.CK  = CK;
  assign \DFF_970.CK  = CK;
  assign \DFF_971.CK  = CK;
  assign \DFF_972.CK  = CK;
  assign \DFF_973.CK  = CK;
  assign \DFF_974.CK  = CK;
  assign \DFF_975.CK  = CK;
  assign \DFF_976.CK  = CK;
  assign \DFF_977.CK  = CK;
  assign \DFF_978.CK  = CK;
  assign \DFF_979.CK  = CK;
  assign \DFF_98.CK  = CK;
  assign \DFF_980.CK  = CK;
  assign \DFF_981.CK  = CK;
  assign \DFF_982.CK  = CK;
  assign \DFF_983.CK  = CK;
  assign \DFF_984.CK  = CK;
  assign \DFF_985.CK  = CK;
  assign \DFF_986.CK  = CK;
  assign \DFF_987.CK  = CK;
  assign \DFF_988.CK  = CK;
  assign \DFF_989.CK  = CK;
  assign \DFF_99.CK  = CK;
  assign \DFF_990.CK  = CK;
  assign \DFF_991.CK  = CK;
  assign \DFF_992.CK  = CK;
  assign \DFF_993.CK  = CK;
  assign \DFF_994.CK  = CK;
  assign \DFF_995.CK  = CK;
  assign \DFF_996.CK  = CK;
  assign \DFF_997.CK  = CK;
  assign \DFF_998.CK  = CK;
  assign \DFF_999.CK  = CK;
  assign WX1001 = TM1;
  assign WX1002 = TM0;
  assign WX1003 = TM1;
  assign WX1004 = TM0;
  assign WX1005 = TM0;
  assign WX10052 = TM1;
  assign WX10053 = TM0;
  assign WX10054 = TM1;
  assign WX10055 = TM0;
  assign WX10056 = TM0;
  assign WX1010 = DATA_9_31;
  assign WX1017 = DATA_9_30;
  assign WX1024 = DATA_9_29;
  assign WX1031 = DATA_9_28;
  assign WX10314 = RESET;
  assign WX10315 = \DFF_1504.D ;
  assign WX10317 = \DFF_1505.D ;
  assign WX10319 = \DFF_1506.D ;
  assign WX10321 = \DFF_1507.D ;
  assign WX10323 = \DFF_1508.D ;
  assign WX10325 = \DFF_1509.D ;
  assign WX10327 = \DFF_1510.D ;
  assign WX10329 = \DFF_1511.D ;
  assign WX10331 = \DFF_1512.D ;
  assign WX10333 = \DFF_1513.D ;
  assign WX10335 = \DFF_1514.D ;
  assign WX10337 = \DFF_1515.D ;
  assign WX10339 = \DFF_1516.D ;
  assign WX10341 = \DFF_1517.D ;
  assign WX10343 = \DFF_1518.D ;
  assign WX10345 = \DFF_1519.D ;
  assign WX10347 = \DFF_1520.D ;
  assign WX10349 = \DFF_1521.D ;
  assign WX10351 = \DFF_1522.D ;
  assign WX10353 = \DFF_1523.D ;
  assign WX10355 = \DFF_1524.D ;
  assign WX10357 = \DFF_1525.D ;
  assign WX10359 = \DFF_1526.D ;
  assign WX10361 = \DFF_1527.D ;
  assign WX10363 = \DFF_1528.D ;
  assign WX10365 = \DFF_1529.D ;
  assign WX10367 = \DFF_1530.D ;
  assign WX10369 = \DFF_1531.D ;
  assign WX10371 = \DFF_1532.D ;
  assign WX10373 = \DFF_1533.D ;
  assign WX10375 = \DFF_1534.D ;
  assign WX10377 = \DFF_1535.D ;
  assign WX1038 = DATA_9_27;
  assign WX1045 = DATA_9_26;
  assign WX1052 = DATA_9_25;
  assign WX1059 = DATA_9_24;
  assign WX1066 = DATA_9_23;
  assign WX1073 = DATA_9_22;
  assign WX1080 = DATA_9_21;
  assign WX10828 = \DFF_1536.D ;
  assign WX10829 = \DFF_1536.Q ;
  assign WX10830 = \DFF_1537.D ;
  assign WX10831 = \DFF_1537.Q ;
  assign WX10832 = \DFF_1538.D ;
  assign WX10833 = \DFF_1538.Q ;
  assign WX10834 = \DFF_1539.D ;
  assign WX10835 = \DFF_1539.Q ;
  assign WX10836 = \DFF_1540.D ;
  assign WX10837 = \DFF_1540.Q ;
  assign WX10838 = \DFF_1541.D ;
  assign WX10839 = \DFF_1541.Q ;
  assign WX10840 = \DFF_1542.D ;
  assign WX10841 = \DFF_1542.Q ;
  assign WX10842 = \DFF_1543.D ;
  assign WX10843 = \DFF_1543.Q ;
  assign WX10844 = \DFF_1544.D ;
  assign WX10845 = \DFF_1544.Q ;
  assign WX10846 = \DFF_1545.D ;
  assign WX10847 = \DFF_1545.Q ;
  assign WX10848 = \DFF_1546.D ;
  assign WX10849 = \DFF_1546.Q ;
  assign WX10850 = \DFF_1547.D ;
  assign WX10851 = \DFF_1547.Q ;
  assign WX10852 = \DFF_1548.D ;
  assign WX10853 = \DFF_1548.Q ;
  assign WX10854 = \DFF_1549.D ;
  assign WX10855 = \DFF_1549.Q ;
  assign WX10856 = \DFF_1550.D ;
  assign WX10857 = \DFF_1550.Q ;
  assign WX10858 = \DFF_1551.D ;
  assign WX10859 = \DFF_1551.Q ;
  assign WX10860 = \DFF_1552.D ;
  assign WX10861 = \DFF_1552.Q ;
  assign WX10862 = \DFF_1553.D ;
  assign WX10863 = \DFF_1553.Q ;
  assign WX10864 = \DFF_1554.D ;
  assign WX10865 = \DFF_1554.Q ;
  assign WX10866 = \DFF_1555.D ;
  assign WX10867 = \DFF_1555.Q ;
  assign WX10868 = \DFF_1556.D ;
  assign WX10869 = \DFF_1556.Q ;
  assign WX1087 = DATA_9_20;
  assign WX10870 = \DFF_1557.D ;
  assign WX10871 = \DFF_1557.Q ;
  assign WX10872 = \DFF_1558.D ;
  assign WX10873 = \DFF_1558.Q ;
  assign WX10874 = \DFF_1559.D ;
  assign WX10875 = \DFF_1559.Q ;
  assign WX10876 = \DFF_1560.D ;
  assign WX10877 = \DFF_1560.Q ;
  assign WX10878 = \DFF_1561.D ;
  assign WX10879 = \DFF_1561.Q ;
  assign WX10880 = \DFF_1562.D ;
  assign WX10881 = \DFF_1562.Q ;
  assign WX10882 = \DFF_1563.D ;
  assign WX10883 = \DFF_1563.Q ;
  assign WX10884 = \DFF_1564.D ;
  assign WX10885 = \DFF_1564.Q ;
  assign WX10886 = \DFF_1565.D ;
  assign WX10887 = \DFF_1565.Q ;
  assign WX10888 = \DFF_1566.D ;
  assign WX10889 = \DFF_1566.Q ;
  assign WX10890 = \DFF_1567.D ;
  assign WX10891 = \DFF_1567.Q ;
  assign WX1094 = DATA_9_19;
  assign WX10988 = \DFF_1568.D ;
  assign WX10989 = \DFF_1568.Q ;
  assign WX10990 = \DFF_1569.D ;
  assign WX10991 = \DFF_1569.Q ;
  assign WX10992 = \DFF_1570.D ;
  assign WX10993 = \DFF_1570.Q ;
  assign WX10994 = \DFF_1571.D ;
  assign WX10995 = \DFF_1571.Q ;
  assign WX10996 = \DFF_1572.D ;
  assign WX10997 = \DFF_1572.Q ;
  assign WX10998 = \DFF_1573.D ;
  assign WX10999 = \DFF_1573.Q ;
  assign WX11000 = \DFF_1574.D ;
  assign WX11001 = \DFF_1574.Q ;
  assign WX11002 = \DFF_1575.D ;
  assign WX11003 = \DFF_1575.Q ;
  assign WX11004 = \DFF_1576.D ;
  assign WX11005 = \DFF_1576.Q ;
  assign WX11006 = \DFF_1577.D ;
  assign WX11007 = \DFF_1577.Q ;
  assign WX11008 = \DFF_1578.D ;
  assign WX11009 = \DFF_1578.Q ;
  assign WX1101 = DATA_9_18;
  assign WX11010 = \DFF_1579.D ;
  assign WX11011 = \DFF_1579.Q ;
  assign WX11012 = \DFF_1580.D ;
  assign WX11013 = \DFF_1580.Q ;
  assign WX11014 = \DFF_1581.D ;
  assign WX11015 = \DFF_1581.Q ;
  assign WX11016 = \DFF_1582.D ;
  assign WX11017 = \DFF_1582.Q ;
  assign WX11018 = \DFF_1583.D ;
  assign WX11019 = \DFF_1583.Q ;
  assign WX11020 = \DFF_1584.D ;
  assign WX11021 = \DFF_1584.Q ;
  assign WX11022 = \DFF_1585.D ;
  assign WX11023 = \DFF_1585.Q ;
  assign WX11024 = \DFF_1586.D ;
  assign WX11025 = \DFF_1586.Q ;
  assign WX11026 = \DFF_1587.D ;
  assign WX11027 = \DFF_1587.Q ;
  assign WX11028 = \DFF_1588.D ;
  assign WX11029 = \DFF_1588.Q ;
  assign WX11030 = \DFF_1589.D ;
  assign WX11031 = \DFF_1589.Q ;
  assign WX11032 = \DFF_1590.D ;
  assign WX11033 = \DFF_1590.Q ;
  assign WX11034 = \DFF_1591.D ;
  assign WX11035 = \DFF_1591.Q ;
  assign WX11036 = \DFF_1592.D ;
  assign WX11037 = \DFF_1592.Q ;
  assign WX11038 = \DFF_1593.D ;
  assign WX11039 = \DFF_1593.Q ;
  assign WX11040 = \DFF_1594.D ;
  assign WX11041 = \DFF_1594.Q ;
  assign WX11042 = \DFF_1595.D ;
  assign WX11043 = \DFF_1595.Q ;
  assign WX11044 = \DFF_1596.D ;
  assign WX11045 = \DFF_1596.Q ;
  assign WX11046 = \DFF_1597.D ;
  assign WX11047 = \DFF_1597.Q ;
  assign WX11048 = \DFF_1598.D ;
  assign WX11049 = \DFF_1598.Q ;
  assign WX11050 = \DFF_1599.D ;
  assign WX11051 = \DFF_1599.Q ;
  assign WX11052 = \DFF_1600.D ;
  assign WX11053 = \DFF_1600.Q ;
  assign WX11054 = \DFF_1601.D ;
  assign WX11055 = \DFF_1601.Q ;
  assign WX11056 = \DFF_1602.D ;
  assign WX11057 = \DFF_1602.Q ;
  assign WX11058 = \DFF_1603.D ;
  assign WX11059 = \DFF_1603.Q ;
  assign WX11060 = \DFF_1604.D ;
  assign WX11061 = \DFF_1604.Q ;
  assign WX11062 = \DFF_1605.D ;
  assign WX11063 = \DFF_1605.Q ;
  assign WX11064 = \DFF_1606.D ;
  assign WX11065 = \DFF_1606.Q ;
  assign WX11066 = \DFF_1607.D ;
  assign WX11067 = \DFF_1607.Q ;
  assign WX11068 = \DFF_1608.D ;
  assign WX11069 = \DFF_1608.Q ;
  assign WX11070 = \DFF_1609.D ;
  assign WX11071 = \DFF_1609.Q ;
  assign WX11072 = \DFF_1610.D ;
  assign WX11073 = \DFF_1610.Q ;
  assign WX11074 = \DFF_1611.D ;
  assign WX11075 = \DFF_1611.Q ;
  assign WX11076 = \DFF_1612.D ;
  assign WX11077 = \DFF_1612.Q ;
  assign WX11078 = \DFF_1613.D ;
  assign WX11079 = \DFF_1613.Q ;
  assign WX1108 = DATA_9_17;
  assign WX11080 = \DFF_1614.D ;
  assign WX11081 = \DFF_1614.Q ;
  assign WX11082 = \DFF_1615.D ;
  assign WX11083 = \DFF_1615.Q ;
  assign WX11084 = \DFF_1616.D ;
  assign WX11085 = \DFF_1616.Q ;
  assign WX11086 = \DFF_1617.D ;
  assign WX11087 = \DFF_1617.Q ;
  assign WX11088 = \DFF_1618.D ;
  assign WX11089 = \DFF_1618.Q ;
  assign WX11090 = \DFF_1619.D ;
  assign WX11091 = \DFF_1619.Q ;
  assign WX11092 = \DFF_1620.D ;
  assign WX11093 = \DFF_1620.Q ;
  assign WX11094 = \DFF_1621.D ;
  assign WX11095 = \DFF_1621.Q ;
  assign WX11096 = \DFF_1622.D ;
  assign WX11097 = \DFF_1622.Q ;
  assign WX11098 = \DFF_1623.D ;
  assign WX11099 = \DFF_1623.Q ;
  assign WX11100 = \DFF_1624.D ;
  assign WX11101 = \DFF_1624.Q ;
  assign WX11102 = \DFF_1625.D ;
  assign WX11103 = \DFF_1625.Q ;
  assign WX11104 = \DFF_1626.D ;
  assign WX11105 = \DFF_1626.Q ;
  assign WX11106 = \DFF_1627.D ;
  assign WX11107 = \DFF_1627.Q ;
  assign WX11108 = \DFF_1628.D ;
  assign WX11109 = \DFF_1628.Q ;
  assign WX11110 = \DFF_1629.D ;
  assign WX11111 = \DFF_1629.Q ;
  assign WX11112 = \DFF_1630.D ;
  assign WX11113 = \DFF_1630.Q ;
  assign WX11114 = \DFF_1631.D ;
  assign WX11115 = \DFF_1631.Q ;
  assign WX11116 = \DFF_1632.D ;
  assign WX11117 = \DFF_1632.Q ;
  assign WX11118 = \DFF_1633.D ;
  assign WX11119 = \DFF_1633.Q ;
  assign WX11120 = \DFF_1634.D ;
  assign WX11121 = \DFF_1634.Q ;
  assign WX11122 = \DFF_1635.D ;
  assign WX11123 = \DFF_1635.Q ;
  assign WX11124 = \DFF_1636.D ;
  assign WX11125 = \DFF_1636.Q ;
  assign WX11126 = \DFF_1637.D ;
  assign WX11127 = \DFF_1637.Q ;
  assign WX11128 = \DFF_1638.D ;
  assign WX11129 = \DFF_1638.Q ;
  assign WX11130 = \DFF_1639.D ;
  assign WX11131 = \DFF_1639.Q ;
  assign WX11132 = \DFF_1640.D ;
  assign WX11133 = \DFF_1640.Q ;
  assign WX11134 = \DFF_1641.D ;
  assign WX11135 = \DFF_1641.Q ;
  assign WX11136 = \DFF_1642.D ;
  assign WX11137 = \DFF_1642.Q ;
  assign WX11138 = \DFF_1643.D ;
  assign WX11139 = \DFF_1643.Q ;
  assign WX11140 = \DFF_1644.D ;
  assign WX11141 = \DFF_1644.Q ;
  assign WX11142 = \DFF_1645.D ;
  assign WX11143 = \DFF_1645.Q ;
  assign WX11144 = \DFF_1646.D ;
  assign WX11145 = \DFF_1646.Q ;
  assign WX11146 = \DFF_1647.D ;
  assign WX11147 = \DFF_1647.Q ;
  assign WX11148 = \DFF_1648.D ;
  assign WX11149 = \DFF_1648.Q ;
  assign WX1115 = DATA_9_16;
  assign WX11150 = \DFF_1649.D ;
  assign WX11151 = \DFF_1649.Q ;
  assign WX11152 = \DFF_1650.D ;
  assign WX11153 = \DFF_1650.Q ;
  assign WX11154 = \DFF_1651.D ;
  assign WX11155 = \DFF_1651.Q ;
  assign WX11156 = \DFF_1652.D ;
  assign WX11157 = \DFF_1652.Q ;
  assign WX11158 = \DFF_1653.D ;
  assign WX11159 = \DFF_1653.Q ;
  assign WX11160 = \DFF_1654.D ;
  assign WX11161 = \DFF_1654.Q ;
  assign WX11162 = \DFF_1655.D ;
  assign WX11163 = \DFF_1655.Q ;
  assign WX11164 = \DFF_1656.D ;
  assign WX11165 = \DFF_1656.Q ;
  assign WX11166 = \DFF_1657.D ;
  assign WX11167 = \DFF_1657.Q ;
  assign WX11168 = \DFF_1658.D ;
  assign WX11169 = \DFF_1658.Q ;
  assign WX11170 = \DFF_1659.D ;
  assign WX11171 = \DFF_1659.Q ;
  assign WX11172 = \DFF_1660.D ;
  assign WX11173 = \DFF_1660.Q ;
  assign WX11174 = \DFF_1661.D ;
  assign WX11175 = \DFF_1661.Q ;
  assign WX11176 = \DFF_1662.D ;
  assign WX11177 = \DFF_1662.Q ;
  assign WX11178 = \DFF_1663.D ;
  assign WX11179 = \DFF_1663.Q ;
  assign WX11180 = \DFF_1664.D ;
  assign WX11181 = \DFF_1664.Q ;
  assign WX11182 = \DFF_1665.D ;
  assign WX11183 = \DFF_1665.Q ;
  assign WX11184 = \DFF_1666.D ;
  assign WX11185 = \DFF_1666.Q ;
  assign WX11186 = \DFF_1667.D ;
  assign WX11187 = \DFF_1667.Q ;
  assign WX11188 = \DFF_1668.D ;
  assign WX11189 = \DFF_1668.Q ;
  assign WX11190 = \DFF_1669.D ;
  assign WX11191 = \DFF_1669.Q ;
  assign WX11192 = \DFF_1670.D ;
  assign WX11193 = \DFF_1670.Q ;
  assign WX11194 = \DFF_1671.D ;
  assign WX11195 = \DFF_1671.Q ;
  assign WX11196 = \DFF_1672.D ;
  assign WX11197 = \DFF_1672.Q ;
  assign WX11198 = \DFF_1673.D ;
  assign WX11199 = \DFF_1673.Q ;
  assign WX11200 = \DFF_1674.D ;
  assign WX11201 = \DFF_1674.Q ;
  assign WX11202 = \DFF_1675.D ;
  assign WX11203 = \DFF_1675.Q ;
  assign WX11204 = \DFF_1676.D ;
  assign WX11205 = \DFF_1676.Q ;
  assign WX11206 = \DFF_1677.D ;
  assign WX11207 = \DFF_1677.Q ;
  assign WX11208 = \DFF_1678.D ;
  assign WX11209 = \DFF_1678.Q ;
  assign WX11210 = \DFF_1679.D ;
  assign WX11211 = \DFF_1679.Q ;
  assign WX11212 = \DFF_1680.D ;
  assign WX11213 = \DFF_1680.Q ;
  assign WX11214 = \DFF_1681.D ;
  assign WX11215 = \DFF_1681.Q ;
  assign WX11216 = \DFF_1682.D ;
  assign WX11217 = \DFF_1682.Q ;
  assign WX11218 = \DFF_1683.D ;
  assign WX11219 = \DFF_1683.Q ;
  assign WX1122 = DATA_9_15;
  assign WX11220 = \DFF_1684.D ;
  assign WX11221 = \DFF_1684.Q ;
  assign WX11222 = \DFF_1685.D ;
  assign WX11223 = \DFF_1685.Q ;
  assign WX11224 = \DFF_1686.D ;
  assign WX11225 = \DFF_1686.Q ;
  assign WX11226 = \DFF_1687.D ;
  assign WX11227 = \DFF_1687.Q ;
  assign WX11228 = \DFF_1688.D ;
  assign WX11229 = \DFF_1688.Q ;
  assign WX11230 = \DFF_1689.D ;
  assign WX11231 = \DFF_1689.Q ;
  assign WX11232 = \DFF_1690.D ;
  assign WX11233 = \DFF_1690.Q ;
  assign WX11234 = \DFF_1691.D ;
  assign WX11235 = \DFF_1691.Q ;
  assign WX11236 = \DFF_1692.D ;
  assign WX11237 = \DFF_1692.Q ;
  assign WX11238 = \DFF_1693.D ;
  assign WX11239 = \DFF_1693.Q ;
  assign WX11240 = \DFF_1694.D ;
  assign WX11241 = \DFF_1694.Q ;
  assign WX11242 = \DFF_1695.D ;
  assign WX11243 = \DFF_1695.Q ;
  assign WX1129 = DATA_9_14;
  assign WX11345 = TM1;
  assign WX11346 = TM0;
  assign WX11347 = TM1;
  assign WX11348 = TM0;
  assign WX11349 = TM0;
  assign WX1136 = DATA_9_13;
  assign WX1143 = DATA_9_12;
  assign WX1150 = DATA_9_11;
  assign WX1157 = DATA_9_10;
  assign WX11607 = RESET;
  assign WX11608 = \DFF_1696.D ;
  assign WX11610 = \DFF_1697.D ;
  assign WX11612 = \DFF_1698.D ;
  assign WX11614 = \DFF_1699.D ;
  assign WX11616 = \DFF_1700.D ;
  assign WX11618 = \DFF_1701.D ;
  assign WX11620 = \DFF_1702.D ;
  assign WX11622 = \DFF_1703.D ;
  assign WX11624 = \DFF_1704.D ;
  assign WX11626 = \DFF_1705.D ;
  assign WX11628 = \DFF_1706.D ;
  assign WX11630 = \DFF_1707.D ;
  assign WX11632 = \DFF_1708.D ;
  assign WX11634 = \DFF_1709.D ;
  assign WX11636 = \DFF_1710.D ;
  assign WX11638 = \DFF_1711.D ;
  assign WX1164 = DATA_9_9;
  assign WX11640 = \DFF_1712.D ;
  assign WX11642 = \DFF_1713.D ;
  assign WX11644 = \DFF_1714.D ;
  assign WX11646 = \DFF_1715.D ;
  assign WX11648 = \DFF_1716.D ;
  assign WX11650 = \DFF_1717.D ;
  assign WX11652 = \DFF_1718.D ;
  assign WX11654 = \DFF_1719.D ;
  assign WX11656 = \DFF_1720.D ;
  assign WX11658 = \DFF_1721.D ;
  assign WX11660 = \DFF_1722.D ;
  assign WX11662 = \DFF_1723.D ;
  assign WX11664 = \DFF_1724.D ;
  assign WX11666 = \DFF_1725.D ;
  assign WX11668 = \DFF_1726.D ;
  assign WX11670 = \DFF_1727.D ;
  assign WX1171 = DATA_9_8;
  assign WX1178 = DATA_9_7;
  assign WX1185 = DATA_9_6;
  assign WX1192 = DATA_9_5;
  assign WX1199 = DATA_9_4;
  assign WX1206 = DATA_9_3;
  assign WX1213 = DATA_9_2;
  assign WX1220 = DATA_9_1;
  assign WX1227 = DATA_9_0;
  assign WX1263 = RESET;
  assign WX1264 = \DFF_160.D ;
  assign WX1266 = \DFF_161.D ;
  assign WX1268 = \DFF_162.D ;
  assign WX1270 = \DFF_163.D ;
  assign WX1272 = \DFF_164.D ;
  assign WX1274 = \DFF_165.D ;
  assign WX1276 = \DFF_166.D ;
  assign WX1278 = \DFF_167.D ;
  assign WX1280 = \DFF_168.D ;
  assign WX1282 = \DFF_169.D ;
  assign WX1284 = \DFF_170.D ;
  assign WX1286 = \DFF_171.D ;
  assign WX1288 = \DFF_172.D ;
  assign WX1290 = \DFF_173.D ;
  assign WX1292 = \DFF_174.D ;
  assign WX1294 = \DFF_175.D ;
  assign WX1296 = \DFF_176.D ;
  assign WX1298 = \DFF_177.D ;
  assign WX1300 = \DFF_178.D ;
  assign WX1302 = \DFF_179.D ;
  assign WX1304 = \DFF_180.D ;
  assign WX1306 = \DFF_181.D ;
  assign WX1308 = \DFF_182.D ;
  assign WX1310 = \DFF_183.D ;
  assign WX1312 = \DFF_184.D ;
  assign WX1314 = \DFF_185.D ;
  assign WX1316 = \DFF_186.D ;
  assign WX1318 = \DFF_187.D ;
  assign WX1320 = \DFF_188.D ;
  assign WX1322 = \DFF_189.D ;
  assign WX1324 = \DFF_190.D ;
  assign WX1326 = \DFF_191.D ;
  assign WX1777 = \DFF_192.D ;
  assign WX1778 = \DFF_192.Q ;
  assign WX1779 = \DFF_193.D ;
  assign WX1780 = \DFF_193.Q ;
  assign WX1781 = \DFF_194.D ;
  assign WX1782 = \DFF_194.Q ;
  assign WX1783 = \DFF_195.D ;
  assign WX1784 = \DFF_195.Q ;
  assign WX1785 = \DFF_196.D ;
  assign WX1786 = \DFF_196.Q ;
  assign WX1787 = \DFF_197.D ;
  assign WX1788 = \DFF_197.Q ;
  assign WX1789 = \DFF_198.D ;
  assign WX1790 = \DFF_198.Q ;
  assign WX1791 = \DFF_199.D ;
  assign WX1792 = \DFF_199.Q ;
  assign WX1793 = \DFF_200.D ;
  assign WX1794 = \DFF_200.Q ;
  assign WX1795 = \DFF_201.D ;
  assign WX1796 = \DFF_201.Q ;
  assign WX1797 = \DFF_202.D ;
  assign WX1798 = \DFF_202.Q ;
  assign WX1799 = \DFF_203.D ;
  assign WX1800 = \DFF_203.Q ;
  assign WX1801 = \DFF_204.D ;
  assign WX1802 = \DFF_204.Q ;
  assign WX1803 = \DFF_205.D ;
  assign WX1804 = \DFF_205.Q ;
  assign WX1805 = \DFF_206.D ;
  assign WX1806 = \DFF_206.Q ;
  assign WX1807 = \DFF_207.D ;
  assign WX1808 = \DFF_207.Q ;
  assign WX1809 = \DFF_208.D ;
  assign WX1810 = \DFF_208.Q ;
  assign WX1811 = \DFF_209.D ;
  assign WX1812 = \DFF_209.Q ;
  assign WX1813 = \DFF_210.D ;
  assign WX1814 = \DFF_210.Q ;
  assign WX1815 = \DFF_211.D ;
  assign WX1816 = \DFF_211.Q ;
  assign WX1817 = \DFF_212.D ;
  assign WX1818 = \DFF_212.Q ;
  assign WX1819 = \DFF_213.D ;
  assign WX1820 = \DFF_213.Q ;
  assign WX1821 = \DFF_214.D ;
  assign WX1822 = \DFF_214.Q ;
  assign WX1823 = \DFF_215.D ;
  assign WX1824 = \DFF_215.Q ;
  assign WX1825 = \DFF_216.D ;
  assign WX1826 = \DFF_216.Q ;
  assign WX1827 = \DFF_217.D ;
  assign WX1828 = \DFF_217.Q ;
  assign WX1829 = \DFF_218.D ;
  assign WX1830 = \DFF_218.Q ;
  assign WX1831 = \DFF_219.D ;
  assign WX1832 = \DFF_219.Q ;
  assign WX1833 = \DFF_220.D ;
  assign WX1834 = \DFF_220.Q ;
  assign WX1835 = \DFF_221.D ;
  assign WX1836 = \DFF_221.Q ;
  assign WX1837 = \DFF_222.D ;
  assign WX1838 = \DFF_222.Q ;
  assign WX1839 = \DFF_223.D ;
  assign WX1840 = \DFF_223.Q ;
  assign WX1937 = \DFF_224.D ;
  assign WX1938 = \DFF_224.Q ;
  assign WX1939 = \DFF_225.D ;
  assign WX1940 = \DFF_225.Q ;
  assign WX1941 = \DFF_226.D ;
  assign WX1942 = \DFF_226.Q ;
  assign WX1943 = \DFF_227.D ;
  assign WX1944 = \DFF_227.Q ;
  assign WX1945 = \DFF_228.D ;
  assign WX1946 = \DFF_228.Q ;
  assign WX1947 = \DFF_229.D ;
  assign WX1948 = \DFF_229.Q ;
  assign WX1949 = \DFF_230.D ;
  assign WX1950 = \DFF_230.Q ;
  assign WX1951 = \DFF_231.D ;
  assign WX1952 = \DFF_231.Q ;
  assign WX1953 = \DFF_232.D ;
  assign WX1954 = \DFF_232.Q ;
  assign WX1955 = \DFF_233.D ;
  assign WX1956 = \DFF_233.Q ;
  assign WX1957 = \DFF_234.D ;
  assign WX1958 = \DFF_234.Q ;
  assign WX1959 = \DFF_235.D ;
  assign WX1960 = \DFF_235.Q ;
  assign WX1961 = \DFF_236.D ;
  assign WX1962 = \DFF_236.Q ;
  assign WX1963 = \DFF_237.D ;
  assign WX1964 = \DFF_237.Q ;
  assign WX1965 = \DFF_238.D ;
  assign WX1966 = \DFF_238.Q ;
  assign WX1967 = \DFF_239.D ;
  assign WX1968 = \DFF_239.Q ;
  assign WX1969 = \DFF_240.D ;
  assign WX1970 = \DFF_240.Q ;
  assign WX1971 = \DFF_241.D ;
  assign WX1972 = \DFF_241.Q ;
  assign WX1973 = \DFF_242.D ;
  assign WX1974 = \DFF_242.Q ;
  assign WX1975 = \DFF_243.D ;
  assign WX1976 = \DFF_243.Q ;
  assign WX1977 = \DFF_244.D ;
  assign WX1978 = \DFF_244.Q ;
  assign WX1979 = \DFF_245.D ;
  assign WX1980 = \DFF_245.Q ;
  assign WX1981 = \DFF_246.D ;
  assign WX1982 = \DFF_246.Q ;
  assign WX1983 = \DFF_247.D ;
  assign WX1984 = \DFF_247.Q ;
  assign WX1985 = \DFF_248.D ;
  assign WX1986 = \DFF_248.Q ;
  assign WX1987 = \DFF_249.D ;
  assign WX1988 = \DFF_249.Q ;
  assign WX1989 = \DFF_250.D ;
  assign WX1990 = \DFF_250.Q ;
  assign WX1991 = \DFF_251.D ;
  assign WX1992 = \DFF_251.Q ;
  assign WX1993 = \DFF_252.D ;
  assign WX1994 = \DFF_252.Q ;
  assign WX1995 = \DFF_253.D ;
  assign WX1996 = \DFF_253.Q ;
  assign WX1997 = \DFF_254.D ;
  assign WX1998 = \DFF_254.Q ;
  assign WX1999 = \DFF_255.D ;
  assign WX2000 = \DFF_255.Q ;
  assign WX2001 = \DFF_256.D ;
  assign WX2002 = \DFF_256.Q ;
  assign WX2003 = \DFF_257.D ;
  assign WX2004 = \DFF_257.Q ;
  assign WX2005 = \DFF_258.D ;
  assign WX2006 = \DFF_258.Q ;
  assign WX2007 = \DFF_259.D ;
  assign WX2008 = \DFF_259.Q ;
  assign WX2009 = \DFF_260.D ;
  assign WX2010 = \DFF_260.Q ;
  assign WX2011 = \DFF_261.D ;
  assign WX2012 = \DFF_261.Q ;
  assign WX2013 = \DFF_262.D ;
  assign WX2014 = \DFF_262.Q ;
  assign WX2015 = \DFF_263.D ;
  assign WX2016 = \DFF_263.Q ;
  assign WX2017 = \DFF_264.D ;
  assign WX2018 = \DFF_264.Q ;
  assign WX2019 = \DFF_265.D ;
  assign WX2020 = \DFF_265.Q ;
  assign WX2021 = \DFF_266.D ;
  assign WX2022 = \DFF_266.Q ;
  assign WX2023 = \DFF_267.D ;
  assign WX2024 = \DFF_267.Q ;
  assign WX2025 = \DFF_268.D ;
  assign WX2026 = \DFF_268.Q ;
  assign WX2027 = \DFF_269.D ;
  assign WX2028 = \DFF_269.Q ;
  assign WX2029 = \DFF_270.D ;
  assign WX2030 = \DFF_270.Q ;
  assign WX2031 = \DFF_271.D ;
  assign WX2032 = \DFF_271.Q ;
  assign WX2033 = \DFF_272.D ;
  assign WX2034 = \DFF_272.Q ;
  assign WX2035 = \DFF_273.D ;
  assign WX2036 = \DFF_273.Q ;
  assign WX2037 = \DFF_274.D ;
  assign WX2038 = \DFF_274.Q ;
  assign WX2039 = \DFF_275.D ;
  assign WX2040 = \DFF_275.Q ;
  assign WX2041 = \DFF_276.D ;
  assign WX2042 = \DFF_276.Q ;
  assign WX2043 = \DFF_277.D ;
  assign WX2044 = \DFF_277.Q ;
  assign WX2045 = \DFF_278.D ;
  assign WX2046 = \DFF_278.Q ;
  assign WX2047 = \DFF_279.D ;
  assign WX2048 = \DFF_279.Q ;
  assign WX2049 = \DFF_280.D ;
  assign WX2050 = \DFF_280.Q ;
  assign WX2051 = \DFF_281.D ;
  assign WX2052 = \DFF_281.Q ;
  assign WX2053 = \DFF_282.D ;
  assign WX2054 = \DFF_282.Q ;
  assign WX2055 = \DFF_283.D ;
  assign WX2056 = \DFF_283.Q ;
  assign WX2057 = \DFF_284.D ;
  assign WX2058 = \DFF_284.Q ;
  assign WX2059 = \DFF_285.D ;
  assign WX2060 = \DFF_285.Q ;
  assign WX2061 = \DFF_286.D ;
  assign WX2062 = \DFF_286.Q ;
  assign WX2063 = \DFF_287.D ;
  assign WX2064 = \DFF_287.Q ;
  assign WX2065 = \DFF_288.D ;
  assign WX2066 = \DFF_288.Q ;
  assign WX2067 = \DFF_289.D ;
  assign WX2068 = \DFF_289.Q ;
  assign WX2069 = \DFF_290.D ;
  assign WX2070 = \DFF_290.Q ;
  assign WX2071 = \DFF_291.D ;
  assign WX2072 = \DFF_291.Q ;
  assign WX2073 = \DFF_292.D ;
  assign WX2074 = \DFF_292.Q ;
  assign WX2075 = \DFF_293.D ;
  assign WX2076 = \DFF_293.Q ;
  assign WX2077 = \DFF_294.D ;
  assign WX2078 = \DFF_294.Q ;
  assign WX2079 = \DFF_295.D ;
  assign WX2080 = \DFF_295.Q ;
  assign WX2081 = \DFF_296.D ;
  assign WX2082 = \DFF_296.Q ;
  assign WX2083 = \DFF_297.D ;
  assign WX2084 = \DFF_297.Q ;
  assign WX2085 = \DFF_298.D ;
  assign WX2086 = \DFF_298.Q ;
  assign WX2087 = \DFF_299.D ;
  assign WX2088 = \DFF_299.Q ;
  assign WX2089 = \DFF_300.D ;
  assign WX2090 = \DFF_300.Q ;
  assign WX2091 = \DFF_301.D ;
  assign WX2092 = \DFF_301.Q ;
  assign WX2093 = \DFF_302.D ;
  assign WX2094 = \DFF_302.Q ;
  assign WX2095 = \DFF_303.D ;
  assign WX2096 = \DFF_303.Q ;
  assign WX2097 = \DFF_304.D ;
  assign WX2098 = \DFF_304.Q ;
  assign WX2099 = \DFF_305.D ;
  assign WX2100 = \DFF_305.Q ;
  assign WX2101 = \DFF_306.D ;
  assign WX2102 = \DFF_306.Q ;
  assign WX2103 = \DFF_307.D ;
  assign WX2104 = \DFF_307.Q ;
  assign WX2105 = \DFF_308.D ;
  assign WX2106 = \DFF_308.Q ;
  assign WX2107 = \DFF_309.D ;
  assign WX2108 = \DFF_309.Q ;
  assign WX2109 = \DFF_310.D ;
  assign WX2110 = \DFF_310.Q ;
  assign WX2111 = \DFF_311.D ;
  assign WX2112 = \DFF_311.Q ;
  assign WX2113 = \DFF_312.D ;
  assign WX2114 = \DFF_312.Q ;
  assign WX2115 = \DFF_313.D ;
  assign WX2116 = \DFF_313.Q ;
  assign WX2117 = \DFF_314.D ;
  assign WX2118 = \DFF_314.Q ;
  assign WX2119 = \DFF_315.D ;
  assign WX2120 = \DFF_315.Q ;
  assign WX2121 = \DFF_316.D ;
  assign WX2122 = \DFF_316.Q ;
  assign WX2123 = \DFF_317.D ;
  assign WX2124 = \DFF_317.Q ;
  assign WX2125 = \DFF_318.D ;
  assign WX2126 = \DFF_318.Q ;
  assign WX2127 = \DFF_319.D ;
  assign WX2128 = \DFF_319.Q ;
  assign WX2129 = \DFF_320.D ;
  assign WX2130 = \DFF_320.Q ;
  assign WX2131 = \DFF_321.D ;
  assign WX2132 = \DFF_321.Q ;
  assign WX2133 = \DFF_322.D ;
  assign WX2134 = \DFF_322.Q ;
  assign WX2135 = \DFF_323.D ;
  assign WX2136 = \DFF_323.Q ;
  assign WX2137 = \DFF_324.D ;
  assign WX2138 = \DFF_324.Q ;
  assign WX2139 = \DFF_325.D ;
  assign WX2140 = \DFF_325.Q ;
  assign WX2141 = \DFF_326.D ;
  assign WX2142 = \DFF_326.Q ;
  assign WX2143 = \DFF_327.D ;
  assign WX2144 = \DFF_327.Q ;
  assign WX2145 = \DFF_328.D ;
  assign WX2146 = \DFF_328.Q ;
  assign WX2147 = \DFF_329.D ;
  assign WX2148 = \DFF_329.Q ;
  assign WX2149 = \DFF_330.D ;
  assign WX2150 = \DFF_330.Q ;
  assign WX2151 = \DFF_331.D ;
  assign WX2152 = \DFF_331.Q ;
  assign WX2153 = \DFF_332.D ;
  assign WX2154 = \DFF_332.Q ;
  assign WX2155 = \DFF_333.D ;
  assign WX2156 = \DFF_333.Q ;
  assign WX2157 = \DFF_334.D ;
  assign WX2158 = \DFF_334.Q ;
  assign WX2159 = \DFF_335.D ;
  assign WX2160 = \DFF_335.Q ;
  assign WX2161 = \DFF_336.D ;
  assign WX2162 = \DFF_336.Q ;
  assign WX2163 = \DFF_337.D ;
  assign WX2164 = \DFF_337.Q ;
  assign WX2165 = \DFF_338.D ;
  assign WX2166 = \DFF_338.Q ;
  assign WX2167 = \DFF_339.D ;
  assign WX2168 = \DFF_339.Q ;
  assign WX2169 = \DFF_340.D ;
  assign WX2170 = \DFF_340.Q ;
  assign WX2171 = \DFF_341.D ;
  assign WX2172 = \DFF_341.Q ;
  assign WX2173 = \DFF_342.D ;
  assign WX2174 = \DFF_342.Q ;
  assign WX2175 = \DFF_343.D ;
  assign WX2176 = \DFF_343.Q ;
  assign WX2177 = \DFF_344.D ;
  assign WX2178 = \DFF_344.Q ;
  assign WX2179 = \DFF_345.D ;
  assign WX2180 = \DFF_345.Q ;
  assign WX2181 = \DFF_346.D ;
  assign WX2182 = \DFF_346.Q ;
  assign WX2183 = \DFF_347.D ;
  assign WX2184 = \DFF_347.Q ;
  assign WX2185 = \DFF_348.D ;
  assign WX2186 = \DFF_348.Q ;
  assign WX2187 = \DFF_349.D ;
  assign WX2188 = \DFF_349.Q ;
  assign WX2189 = \DFF_350.D ;
  assign WX2190 = \DFF_350.Q ;
  assign WX2191 = \DFF_351.D ;
  assign WX2192 = \DFF_351.Q ;
  assign WX2294 = TM1;
  assign WX2295 = TM0;
  assign WX2296 = TM1;
  assign WX2297 = TM0;
  assign WX2298 = TM0;
  assign WX2556 = RESET;
  assign WX2557 = \DFF_352.D ;
  assign WX2559 = \DFF_353.D ;
  assign WX2561 = \DFF_354.D ;
  assign WX2563 = \DFF_355.D ;
  assign WX2565 = \DFF_356.D ;
  assign WX2567 = \DFF_357.D ;
  assign WX2569 = \DFF_358.D ;
  assign WX2571 = \DFF_359.D ;
  assign WX2573 = \DFF_360.D ;
  assign WX2575 = \DFF_361.D ;
  assign WX2577 = \DFF_362.D ;
  assign WX2579 = \DFF_363.D ;
  assign WX2581 = \DFF_364.D ;
  assign WX2583 = \DFF_365.D ;
  assign WX2585 = \DFF_366.D ;
  assign WX2587 = \DFF_367.D ;
  assign WX2589 = \DFF_368.D ;
  assign WX2591 = \DFF_369.D ;
  assign WX2593 = \DFF_370.D ;
  assign WX2595 = \DFF_371.D ;
  assign WX2597 = \DFF_372.D ;
  assign WX2599 = \DFF_373.D ;
  assign WX2601 = \DFF_374.D ;
  assign WX2603 = \DFF_375.D ;
  assign WX2605 = \DFF_376.D ;
  assign WX2607 = \DFF_377.D ;
  assign WX2609 = \DFF_378.D ;
  assign WX2611 = \DFF_379.D ;
  assign WX2613 = \DFF_380.D ;
  assign WX2615 = \DFF_381.D ;
  assign WX2617 = \DFF_382.D ;
  assign WX2619 = \DFF_383.D ;
  assign WX3070 = \DFF_384.D ;
  assign WX3071 = \DFF_384.Q ;
  assign WX3072 = \DFF_385.D ;
  assign WX3073 = \DFF_385.Q ;
  assign WX3074 = \DFF_386.D ;
  assign WX3075 = \DFF_386.Q ;
  assign WX3076 = \DFF_387.D ;
  assign WX3077 = \DFF_387.Q ;
  assign WX3078 = \DFF_388.D ;
  assign WX3079 = \DFF_388.Q ;
  assign WX3080 = \DFF_389.D ;
  assign WX3081 = \DFF_389.Q ;
  assign WX3082 = \DFF_390.D ;
  assign WX3083 = \DFF_390.Q ;
  assign WX3084 = \DFF_391.D ;
  assign WX3085 = \DFF_391.Q ;
  assign WX3086 = \DFF_392.D ;
  assign WX3087 = \DFF_392.Q ;
  assign WX3088 = \DFF_393.D ;
  assign WX3089 = \DFF_393.Q ;
  assign WX3090 = \DFF_394.D ;
  assign WX3091 = \DFF_394.Q ;
  assign WX3092 = \DFF_395.D ;
  assign WX3093 = \DFF_395.Q ;
  assign WX3094 = \DFF_396.D ;
  assign WX3095 = \DFF_396.Q ;
  assign WX3096 = \DFF_397.D ;
  assign WX3097 = \DFF_397.Q ;
  assign WX3098 = \DFF_398.D ;
  assign WX3099 = \DFF_398.Q ;
  assign WX3100 = \DFF_399.D ;
  assign WX3101 = \DFF_399.Q ;
  assign WX3102 = \DFF_400.D ;
  assign WX3103 = \DFF_400.Q ;
  assign WX3104 = \DFF_401.D ;
  assign WX3105 = \DFF_401.Q ;
  assign WX3106 = \DFF_402.D ;
  assign WX3107 = \DFF_402.Q ;
  assign WX3108 = \DFF_403.D ;
  assign WX3109 = \DFF_403.Q ;
  assign WX3110 = \DFF_404.D ;
  assign WX3111 = \DFF_404.Q ;
  assign WX3112 = \DFF_405.D ;
  assign WX3113 = \DFF_405.Q ;
  assign WX3114 = \DFF_406.D ;
  assign WX3115 = \DFF_406.Q ;
  assign WX3116 = \DFF_407.D ;
  assign WX3117 = \DFF_407.Q ;
  assign WX3118 = \DFF_408.D ;
  assign WX3119 = \DFF_408.Q ;
  assign WX3120 = \DFF_409.D ;
  assign WX3121 = \DFF_409.Q ;
  assign WX3122 = \DFF_410.D ;
  assign WX3123 = \DFF_410.Q ;
  assign WX3124 = \DFF_411.D ;
  assign WX3125 = \DFF_411.Q ;
  assign WX3126 = \DFF_412.D ;
  assign WX3127 = \DFF_412.Q ;
  assign WX3128 = \DFF_413.D ;
  assign WX3129 = \DFF_413.Q ;
  assign WX3130 = \DFF_414.D ;
  assign WX3131 = \DFF_414.Q ;
  assign WX3132 = \DFF_415.D ;
  assign WX3133 = \DFF_415.Q ;
  assign WX3230 = \DFF_416.D ;
  assign WX3231 = \DFF_416.Q ;
  assign WX3232 = \DFF_417.D ;
  assign WX3233 = \DFF_417.Q ;
  assign WX3234 = \DFF_418.D ;
  assign WX3235 = \DFF_418.Q ;
  assign WX3236 = \DFF_419.D ;
  assign WX3237 = \DFF_419.Q ;
  assign WX3238 = \DFF_420.D ;
  assign WX3239 = \DFF_420.Q ;
  assign WX3240 = \DFF_421.D ;
  assign WX3241 = \DFF_421.Q ;
  assign WX3242 = \DFF_422.D ;
  assign WX3243 = \DFF_422.Q ;
  assign WX3244 = \DFF_423.D ;
  assign WX3245 = \DFF_423.Q ;
  assign WX3246 = \DFF_424.D ;
  assign WX3247 = \DFF_424.Q ;
  assign WX3248 = \DFF_425.D ;
  assign WX3249 = \DFF_425.Q ;
  assign WX3250 = \DFF_426.D ;
  assign WX3251 = \DFF_426.Q ;
  assign WX3252 = \DFF_427.D ;
  assign WX3253 = \DFF_427.Q ;
  assign WX3254 = \DFF_428.D ;
  assign WX3255 = \DFF_428.Q ;
  assign WX3256 = \DFF_429.D ;
  assign WX3257 = \DFF_429.Q ;
  assign WX3258 = \DFF_430.D ;
  assign WX3259 = \DFF_430.Q ;
  assign WX3260 = \DFF_431.D ;
  assign WX3261 = \DFF_431.Q ;
  assign WX3262 = \DFF_432.D ;
  assign WX3263 = \DFF_432.Q ;
  assign WX3264 = \DFF_433.D ;
  assign WX3265 = \DFF_433.Q ;
  assign WX3266 = \DFF_434.D ;
  assign WX3267 = \DFF_434.Q ;
  assign WX3268 = \DFF_435.D ;
  assign WX3269 = \DFF_435.Q ;
  assign WX3270 = \DFF_436.D ;
  assign WX3271 = \DFF_436.Q ;
  assign WX3272 = \DFF_437.D ;
  assign WX3273 = \DFF_437.Q ;
  assign WX3274 = \DFF_438.D ;
  assign WX3275 = \DFF_438.Q ;
  assign WX3276 = \DFF_439.D ;
  assign WX3277 = \DFF_439.Q ;
  assign WX3278 = \DFF_440.D ;
  assign WX3279 = \DFF_440.Q ;
  assign WX3280 = \DFF_441.D ;
  assign WX3281 = \DFF_441.Q ;
  assign WX3282 = \DFF_442.D ;
  assign WX3283 = \DFF_442.Q ;
  assign WX3284 = \DFF_443.D ;
  assign WX3285 = \DFF_443.Q ;
  assign WX3286 = \DFF_444.D ;
  assign WX3287 = \DFF_444.Q ;
  assign WX3288 = \DFF_445.D ;
  assign WX3289 = \DFF_445.Q ;
  assign WX3290 = \DFF_446.D ;
  assign WX3291 = \DFF_446.Q ;
  assign WX3292 = \DFF_447.D ;
  assign WX3293 = \DFF_447.Q ;
  assign WX3294 = \DFF_448.D ;
  assign WX3295 = \DFF_448.Q ;
  assign WX3296 = \DFF_449.D ;
  assign WX3297 = \DFF_449.Q ;
  assign WX3298 = \DFF_450.D ;
  assign WX3299 = \DFF_450.Q ;
  assign WX3300 = \DFF_451.D ;
  assign WX3301 = \DFF_451.Q ;
  assign WX3302 = \DFF_452.D ;
  assign WX3303 = \DFF_452.Q ;
  assign WX3304 = \DFF_453.D ;
  assign WX3305 = \DFF_453.Q ;
  assign WX3306 = \DFF_454.D ;
  assign WX3307 = \DFF_454.Q ;
  assign WX3308 = \DFF_455.D ;
  assign WX3309 = \DFF_455.Q ;
  assign WX3310 = \DFF_456.D ;
  assign WX3311 = \DFF_456.Q ;
  assign WX3312 = \DFF_457.D ;
  assign WX3313 = \DFF_457.Q ;
  assign WX3314 = \DFF_458.D ;
  assign WX3315 = \DFF_458.Q ;
  assign WX3316 = \DFF_459.D ;
  assign WX3317 = \DFF_459.Q ;
  assign WX3318 = \DFF_460.D ;
  assign WX3319 = \DFF_460.Q ;
  assign WX3320 = \DFF_461.D ;
  assign WX3321 = \DFF_461.Q ;
  assign WX3322 = \DFF_462.D ;
  assign WX3323 = \DFF_462.Q ;
  assign WX3324 = \DFF_463.D ;
  assign WX3325 = \DFF_463.Q ;
  assign WX3326 = \DFF_464.D ;
  assign WX3327 = \DFF_464.Q ;
  assign WX3328 = \DFF_465.D ;
  assign WX3329 = \DFF_465.Q ;
  assign WX3330 = \DFF_466.D ;
  assign WX3331 = \DFF_466.Q ;
  assign WX3332 = \DFF_467.D ;
  assign WX3333 = \DFF_467.Q ;
  assign WX3334 = \DFF_468.D ;
  assign WX3335 = \DFF_468.Q ;
  assign WX3336 = \DFF_469.D ;
  assign WX3337 = \DFF_469.Q ;
  assign WX3338 = \DFF_470.D ;
  assign WX3339 = \DFF_470.Q ;
  assign WX3340 = \DFF_471.D ;
  assign WX3341 = \DFF_471.Q ;
  assign WX3342 = \DFF_472.D ;
  assign WX3343 = \DFF_472.Q ;
  assign WX3344 = \DFF_473.D ;
  assign WX3345 = \DFF_473.Q ;
  assign WX3346 = \DFF_474.D ;
  assign WX3347 = \DFF_474.Q ;
  assign WX3348 = \DFF_475.D ;
  assign WX3349 = \DFF_475.Q ;
  assign WX3350 = \DFF_476.D ;
  assign WX3351 = \DFF_476.Q ;
  assign WX3352 = \DFF_477.D ;
  assign WX3353 = \DFF_477.Q ;
  assign WX3354 = \DFF_478.D ;
  assign WX3355 = \DFF_478.Q ;
  assign WX3356 = \DFF_479.D ;
  assign WX3357 = \DFF_479.Q ;
  assign WX3358 = \DFF_480.D ;
  assign WX3359 = \DFF_480.Q ;
  assign WX3360 = \DFF_481.D ;
  assign WX3361 = \DFF_481.Q ;
  assign WX3362 = \DFF_482.D ;
  assign WX3363 = \DFF_482.Q ;
  assign WX3364 = \DFF_483.D ;
  assign WX3365 = \DFF_483.Q ;
  assign WX3366 = \DFF_484.D ;
  assign WX3367 = \DFF_484.Q ;
  assign WX3368 = \DFF_485.D ;
  assign WX3369 = \DFF_485.Q ;
  assign WX3370 = \DFF_486.D ;
  assign WX3371 = \DFF_486.Q ;
  assign WX3372 = \DFF_487.D ;
  assign WX3373 = \DFF_487.Q ;
  assign WX3374 = \DFF_488.D ;
  assign WX3375 = \DFF_488.Q ;
  assign WX3376 = \DFF_489.D ;
  assign WX3377 = \DFF_489.Q ;
  assign WX3378 = \DFF_490.D ;
  assign WX3379 = \DFF_490.Q ;
  assign WX3380 = \DFF_491.D ;
  assign WX3381 = \DFF_491.Q ;
  assign WX3382 = \DFF_492.D ;
  assign WX3383 = \DFF_492.Q ;
  assign WX3384 = \DFF_493.D ;
  assign WX3385 = \DFF_493.Q ;
  assign WX3386 = \DFF_494.D ;
  assign WX3387 = \DFF_494.Q ;
  assign WX3388 = \DFF_495.D ;
  assign WX3389 = \DFF_495.Q ;
  assign WX3390 = \DFF_496.D ;
  assign WX3391 = \DFF_496.Q ;
  assign WX3392 = \DFF_497.D ;
  assign WX3393 = \DFF_497.Q ;
  assign WX3394 = \DFF_498.D ;
  assign WX3395 = \DFF_498.Q ;
  assign WX3396 = \DFF_499.D ;
  assign WX3397 = \DFF_499.Q ;
  assign WX3398 = \DFF_500.D ;
  assign WX3399 = \DFF_500.Q ;
  assign WX3400 = \DFF_501.D ;
  assign WX3401 = \DFF_501.Q ;
  assign WX3402 = \DFF_502.D ;
  assign WX3403 = \DFF_502.Q ;
  assign WX3404 = \DFF_503.D ;
  assign WX3405 = \DFF_503.Q ;
  assign WX3406 = \DFF_504.D ;
  assign WX3407 = \DFF_504.Q ;
  assign WX3408 = \DFF_505.D ;
  assign WX3409 = \DFF_505.Q ;
  assign WX3410 = \DFF_506.D ;
  assign WX3411 = \DFF_506.Q ;
  assign WX3412 = \DFF_507.D ;
  assign WX3413 = \DFF_507.Q ;
  assign WX3414 = \DFF_508.D ;
  assign WX3415 = \DFF_508.Q ;
  assign WX3416 = \DFF_509.D ;
  assign WX3417 = \DFF_509.Q ;
  assign WX3418 = \DFF_510.D ;
  assign WX3419 = \DFF_510.Q ;
  assign WX3420 = \DFF_511.D ;
  assign WX3421 = \DFF_511.Q ;
  assign WX3422 = \DFF_512.D ;
  assign WX3423 = \DFF_512.Q ;
  assign WX3424 = \DFF_513.D ;
  assign WX3425 = \DFF_513.Q ;
  assign WX3426 = \DFF_514.D ;
  assign WX3427 = \DFF_514.Q ;
  assign WX3428 = \DFF_515.D ;
  assign WX3429 = \DFF_515.Q ;
  assign WX3430 = \DFF_516.D ;
  assign WX3431 = \DFF_516.Q ;
  assign WX3432 = \DFF_517.D ;
  assign WX3433 = \DFF_517.Q ;
  assign WX3434 = \DFF_518.D ;
  assign WX3435 = \DFF_518.Q ;
  assign WX3436 = \DFF_519.D ;
  assign WX3437 = \DFF_519.Q ;
  assign WX3438 = \DFF_520.D ;
  assign WX3439 = \DFF_520.Q ;
  assign WX3440 = \DFF_521.D ;
  assign WX3441 = \DFF_521.Q ;
  assign WX3442 = \DFF_522.D ;
  assign WX3443 = \DFF_522.Q ;
  assign WX3444 = \DFF_523.D ;
  assign WX3445 = \DFF_523.Q ;
  assign WX3446 = \DFF_524.D ;
  assign WX3447 = \DFF_524.Q ;
  assign WX3448 = \DFF_525.D ;
  assign WX3449 = \DFF_525.Q ;
  assign WX3450 = \DFF_526.D ;
  assign WX3451 = \DFF_526.Q ;
  assign WX3452 = \DFF_527.D ;
  assign WX3453 = \DFF_527.Q ;
  assign WX3454 = \DFF_528.D ;
  assign WX3455 = \DFF_528.Q ;
  assign WX3456 = \DFF_529.D ;
  assign WX3457 = \DFF_529.Q ;
  assign WX3458 = \DFF_530.D ;
  assign WX3459 = \DFF_530.Q ;
  assign WX3460 = \DFF_531.D ;
  assign WX3461 = \DFF_531.Q ;
  assign WX3462 = \DFF_532.D ;
  assign WX3463 = \DFF_532.Q ;
  assign WX3464 = \DFF_533.D ;
  assign WX3465 = \DFF_533.Q ;
  assign WX3466 = \DFF_534.D ;
  assign WX3467 = \DFF_534.Q ;
  assign WX3468 = \DFF_535.D ;
  assign WX3469 = \DFF_535.Q ;
  assign WX3470 = \DFF_536.D ;
  assign WX3471 = \DFF_536.Q ;
  assign WX3472 = \DFF_537.D ;
  assign WX3473 = \DFF_537.Q ;
  assign WX3474 = \DFF_538.D ;
  assign WX3475 = \DFF_538.Q ;
  assign WX3476 = \DFF_539.D ;
  assign WX3477 = \DFF_539.Q ;
  assign WX3478 = \DFF_540.D ;
  assign WX3479 = \DFF_540.Q ;
  assign WX3480 = \DFF_541.D ;
  assign WX3481 = \DFF_541.Q ;
  assign WX3482 = \DFF_542.D ;
  assign WX3483 = \DFF_542.Q ;
  assign WX3484 = \DFF_543.D ;
  assign WX3485 = \DFF_543.Q ;
  assign WX3587 = TM1;
  assign WX3588 = TM0;
  assign WX3589 = TM1;
  assign WX3590 = TM0;
  assign WX3591 = TM0;
  assign WX3849 = RESET;
  assign WX3850 = \DFF_544.D ;
  assign WX3852 = \DFF_545.D ;
  assign WX3854 = \DFF_546.D ;
  assign WX3856 = \DFF_547.D ;
  assign WX3858 = \DFF_548.D ;
  assign WX3860 = \DFF_549.D ;
  assign WX3862 = \DFF_550.D ;
  assign WX3864 = \DFF_551.D ;
  assign WX3866 = \DFF_552.D ;
  assign WX3868 = \DFF_553.D ;
  assign WX3870 = \DFF_554.D ;
  assign WX3872 = \DFF_555.D ;
  assign WX3874 = \DFF_556.D ;
  assign WX3876 = \DFF_557.D ;
  assign WX3878 = \DFF_558.D ;
  assign WX3880 = \DFF_559.D ;
  assign WX3882 = \DFF_560.D ;
  assign WX3884 = \DFF_561.D ;
  assign WX3886 = \DFF_562.D ;
  assign WX3888 = \DFF_563.D ;
  assign WX3890 = \DFF_564.D ;
  assign WX3892 = \DFF_565.D ;
  assign WX3894 = \DFF_566.D ;
  assign WX3896 = \DFF_567.D ;
  assign WX3898 = \DFF_568.D ;
  assign WX3900 = \DFF_569.D ;
  assign WX3902 = \DFF_570.D ;
  assign WX3904 = \DFF_571.D ;
  assign WX3906 = \DFF_572.D ;
  assign WX3908 = \DFF_573.D ;
  assign WX3910 = \DFF_574.D ;
  assign WX3912 = \DFF_575.D ;
  assign WX4363 = \DFF_576.D ;
  assign WX4364 = \DFF_576.Q ;
  assign WX4365 = \DFF_577.D ;
  assign WX4366 = \DFF_577.Q ;
  assign WX4367 = \DFF_578.D ;
  assign WX4368 = \DFF_578.Q ;
  assign WX4369 = \DFF_579.D ;
  assign WX4370 = \DFF_579.Q ;
  assign WX4371 = \DFF_580.D ;
  assign WX4372 = \DFF_580.Q ;
  assign WX4373 = \DFF_581.D ;
  assign WX4374 = \DFF_581.Q ;
  assign WX4375 = \DFF_582.D ;
  assign WX4376 = \DFF_582.Q ;
  assign WX4377 = \DFF_583.D ;
  assign WX4378 = \DFF_583.Q ;
  assign WX4379 = \DFF_584.D ;
  assign WX4380 = \DFF_584.Q ;
  assign WX4381 = \DFF_585.D ;
  assign WX4382 = \DFF_585.Q ;
  assign WX4383 = \DFF_586.D ;
  assign WX4384 = \DFF_586.Q ;
  assign WX4385 = \DFF_587.D ;
  assign WX4386 = \DFF_587.Q ;
  assign WX4387 = \DFF_588.D ;
  assign WX4388 = \DFF_588.Q ;
  assign WX4389 = \DFF_589.D ;
  assign WX4390 = \DFF_589.Q ;
  assign WX4391 = \DFF_590.D ;
  assign WX4392 = \DFF_590.Q ;
  assign WX4393 = \DFF_591.D ;
  assign WX4394 = \DFF_591.Q ;
  assign WX4395 = \DFF_592.D ;
  assign WX4396 = \DFF_592.Q ;
  assign WX4397 = \DFF_593.D ;
  assign WX4398 = \DFF_593.Q ;
  assign WX4399 = \DFF_594.D ;
  assign WX4400 = \DFF_594.Q ;
  assign WX4401 = \DFF_595.D ;
  assign WX4402 = \DFF_595.Q ;
  assign WX4403 = \DFF_596.D ;
  assign WX4404 = \DFF_596.Q ;
  assign WX4405 = \DFF_597.D ;
  assign WX4406 = \DFF_597.Q ;
  assign WX4407 = \DFF_598.D ;
  assign WX4408 = \DFF_598.Q ;
  assign WX4409 = \DFF_599.D ;
  assign WX4410 = \DFF_599.Q ;
  assign WX4411 = \DFF_600.D ;
  assign WX4412 = \DFF_600.Q ;
  assign WX4413 = \DFF_601.D ;
  assign WX4414 = \DFF_601.Q ;
  assign WX4415 = \DFF_602.D ;
  assign WX4416 = \DFF_602.Q ;
  assign WX4417 = \DFF_603.D ;
  assign WX4418 = \DFF_603.Q ;
  assign WX4419 = \DFF_604.D ;
  assign WX4420 = \DFF_604.Q ;
  assign WX4421 = \DFF_605.D ;
  assign WX4422 = \DFF_605.Q ;
  assign WX4423 = \DFF_606.D ;
  assign WX4424 = \DFF_606.Q ;
  assign WX4425 = \DFF_607.D ;
  assign WX4426 = \DFF_607.Q ;
  assign WX4523 = \DFF_608.D ;
  assign WX4524 = \DFF_608.Q ;
  assign WX4525 = \DFF_609.D ;
  assign WX4526 = \DFF_609.Q ;
  assign WX4527 = \DFF_610.D ;
  assign WX4528 = \DFF_610.Q ;
  assign WX4529 = \DFF_611.D ;
  assign WX4530 = \DFF_611.Q ;
  assign WX4531 = \DFF_612.D ;
  assign WX4532 = \DFF_612.Q ;
  assign WX4533 = \DFF_613.D ;
  assign WX4534 = \DFF_613.Q ;
  assign WX4535 = \DFF_614.D ;
  assign WX4536 = \DFF_614.Q ;
  assign WX4537 = \DFF_615.D ;
  assign WX4538 = \DFF_615.Q ;
  assign WX4539 = \DFF_616.D ;
  assign WX4540 = \DFF_616.Q ;
  assign WX4541 = \DFF_617.D ;
  assign WX4542 = \DFF_617.Q ;
  assign WX4543 = \DFF_618.D ;
  assign WX4544 = \DFF_618.Q ;
  assign WX4545 = \DFF_619.D ;
  assign WX4546 = \DFF_619.Q ;
  assign WX4547 = \DFF_620.D ;
  assign WX4548 = \DFF_620.Q ;
  assign WX4549 = \DFF_621.D ;
  assign WX4550 = \DFF_621.Q ;
  assign WX4551 = \DFF_622.D ;
  assign WX4552 = \DFF_622.Q ;
  assign WX4553 = \DFF_623.D ;
  assign WX4554 = \DFF_623.Q ;
  assign WX4555 = \DFF_624.D ;
  assign WX4556 = \DFF_624.Q ;
  assign WX4557 = \DFF_625.D ;
  assign WX4558 = \DFF_625.Q ;
  assign WX4559 = \DFF_626.D ;
  assign WX4560 = \DFF_626.Q ;
  assign WX4561 = \DFF_627.D ;
  assign WX4562 = \DFF_627.Q ;
  assign WX4563 = \DFF_628.D ;
  assign WX4564 = \DFF_628.Q ;
  assign WX4565 = \DFF_629.D ;
  assign WX4566 = \DFF_629.Q ;
  assign WX4567 = \DFF_630.D ;
  assign WX4568 = \DFF_630.Q ;
  assign WX4569 = \DFF_631.D ;
  assign WX4570 = \DFF_631.Q ;
  assign WX4571 = \DFF_632.D ;
  assign WX4572 = \DFF_632.Q ;
  assign WX4573 = \DFF_633.D ;
  assign WX4574 = \DFF_633.Q ;
  assign WX4575 = \DFF_634.D ;
  assign WX4576 = \DFF_634.Q ;
  assign WX4577 = \DFF_635.D ;
  assign WX4578 = \DFF_635.Q ;
  assign WX4579 = \DFF_636.D ;
  assign WX4580 = \DFF_636.Q ;
  assign WX4581 = \DFF_637.D ;
  assign WX4582 = \DFF_637.Q ;
  assign WX4583 = \DFF_638.D ;
  assign WX4584 = \DFF_638.Q ;
  assign WX4585 = \DFF_639.D ;
  assign WX4586 = \DFF_639.Q ;
  assign WX4587 = \DFF_640.D ;
  assign WX4588 = \DFF_640.Q ;
  assign WX4589 = \DFF_641.D ;
  assign WX4590 = \DFF_641.Q ;
  assign WX4591 = \DFF_642.D ;
  assign WX4592 = \DFF_642.Q ;
  assign WX4593 = \DFF_643.D ;
  assign WX4594 = \DFF_643.Q ;
  assign WX4595 = \DFF_644.D ;
  assign WX4596 = \DFF_644.Q ;
  assign WX4597 = \DFF_645.D ;
  assign WX4598 = \DFF_645.Q ;
  assign WX4599 = \DFF_646.D ;
  assign WX4600 = \DFF_646.Q ;
  assign WX4601 = \DFF_647.D ;
  assign WX4602 = \DFF_647.Q ;
  assign WX4603 = \DFF_648.D ;
  assign WX4604 = \DFF_648.Q ;
  assign WX4605 = \DFF_649.D ;
  assign WX4606 = \DFF_649.Q ;
  assign WX4607 = \DFF_650.D ;
  assign WX4608 = \DFF_650.Q ;
  assign WX4609 = \DFF_651.D ;
  assign WX4610 = \DFF_651.Q ;
  assign WX4611 = \DFF_652.D ;
  assign WX4612 = \DFF_652.Q ;
  assign WX4613 = \DFF_653.D ;
  assign WX4614 = \DFF_653.Q ;
  assign WX4615 = \DFF_654.D ;
  assign WX4616 = \DFF_654.Q ;
  assign WX4617 = \DFF_655.D ;
  assign WX4618 = \DFF_655.Q ;
  assign WX4619 = \DFF_656.D ;
  assign WX4620 = \DFF_656.Q ;
  assign WX4621 = \DFF_657.D ;
  assign WX4622 = \DFF_657.Q ;
  assign WX4623 = \DFF_658.D ;
  assign WX4624 = \DFF_658.Q ;
  assign WX4625 = \DFF_659.D ;
  assign WX4626 = \DFF_659.Q ;
  assign WX4627 = \DFF_660.D ;
  assign WX4628 = \DFF_660.Q ;
  assign WX4629 = \DFF_661.D ;
  assign WX4630 = \DFF_661.Q ;
  assign WX4631 = \DFF_662.D ;
  assign WX4632 = \DFF_662.Q ;
  assign WX4633 = \DFF_663.D ;
  assign WX4634 = \DFF_663.Q ;
  assign WX4635 = \DFF_664.D ;
  assign WX4636 = \DFF_664.Q ;
  assign WX4637 = \DFF_665.D ;
  assign WX4638 = \DFF_665.Q ;
  assign WX4639 = \DFF_666.D ;
  assign WX4640 = \DFF_666.Q ;
  assign WX4641 = \DFF_667.D ;
  assign WX4642 = \DFF_667.Q ;
  assign WX4643 = \DFF_668.D ;
  assign WX4644 = \DFF_668.Q ;
  assign WX4645 = \DFF_669.D ;
  assign WX4646 = \DFF_669.Q ;
  assign WX4647 = \DFF_670.D ;
  assign WX4648 = \DFF_670.Q ;
  assign WX4649 = \DFF_671.D ;
  assign WX4650 = \DFF_671.Q ;
  assign WX4651 = \DFF_672.D ;
  assign WX4652 = \DFF_672.Q ;
  assign WX4653 = \DFF_673.D ;
  assign WX4654 = \DFF_673.Q ;
  assign WX4655 = \DFF_674.D ;
  assign WX4656 = \DFF_674.Q ;
  assign WX4657 = \DFF_675.D ;
  assign WX4658 = \DFF_675.Q ;
  assign WX4659 = \DFF_676.D ;
  assign WX4660 = \DFF_676.Q ;
  assign WX4661 = \DFF_677.D ;
  assign WX4662 = \DFF_677.Q ;
  assign WX4663 = \DFF_678.D ;
  assign WX4664 = \DFF_678.Q ;
  assign WX4665 = \DFF_679.D ;
  assign WX4666 = \DFF_679.Q ;
  assign WX4667 = \DFF_680.D ;
  assign WX4668 = \DFF_680.Q ;
  assign WX4669 = \DFF_681.D ;
  assign WX4670 = \DFF_681.Q ;
  assign WX4671 = \DFF_682.D ;
  assign WX4672 = \DFF_682.Q ;
  assign WX4673 = \DFF_683.D ;
  assign WX4674 = \DFF_683.Q ;
  assign WX4675 = \DFF_684.D ;
  assign WX4676 = \DFF_684.Q ;
  assign WX4677 = \DFF_685.D ;
  assign WX4678 = \DFF_685.Q ;
  assign WX4679 = \DFF_686.D ;
  assign WX4680 = \DFF_686.Q ;
  assign WX4681 = \DFF_687.D ;
  assign WX4682 = \DFF_687.Q ;
  assign WX4683 = \DFF_688.D ;
  assign WX4684 = \DFF_688.Q ;
  assign WX4685 = \DFF_689.D ;
  assign WX4686 = \DFF_689.Q ;
  assign WX4687 = \DFF_690.D ;
  assign WX4688 = \DFF_690.Q ;
  assign WX4689 = \DFF_691.D ;
  assign WX4690 = \DFF_691.Q ;
  assign WX4691 = \DFF_692.D ;
  assign WX4692 = \DFF_692.Q ;
  assign WX4693 = \DFF_693.D ;
  assign WX4694 = \DFF_693.Q ;
  assign WX4695 = \DFF_694.D ;
  assign WX4696 = \DFF_694.Q ;
  assign WX4697 = \DFF_695.D ;
  assign WX4698 = \DFF_695.Q ;
  assign WX4699 = \DFF_696.D ;
  assign WX4700 = \DFF_696.Q ;
  assign WX4701 = \DFF_697.D ;
  assign WX4702 = \DFF_697.Q ;
  assign WX4703 = \DFF_698.D ;
  assign WX4704 = \DFF_698.Q ;
  assign WX4705 = \DFF_699.D ;
  assign WX4706 = \DFF_699.Q ;
  assign WX4707 = \DFF_700.D ;
  assign WX4708 = \DFF_700.Q ;
  assign WX4709 = \DFF_701.D ;
  assign WX4710 = \DFF_701.Q ;
  assign WX4711 = \DFF_702.D ;
  assign WX4712 = \DFF_702.Q ;
  assign WX4713 = \DFF_703.D ;
  assign WX4714 = \DFF_703.Q ;
  assign WX4715 = \DFF_704.D ;
  assign WX4716 = \DFF_704.Q ;
  assign WX4717 = \DFF_705.D ;
  assign WX4718 = \DFF_705.Q ;
  assign WX4719 = \DFF_706.D ;
  assign WX4720 = \DFF_706.Q ;
  assign WX4721 = \DFF_707.D ;
  assign WX4722 = \DFF_707.Q ;
  assign WX4723 = \DFF_708.D ;
  assign WX4724 = \DFF_708.Q ;
  assign WX4725 = \DFF_709.D ;
  assign WX4726 = \DFF_709.Q ;
  assign WX4727 = \DFF_710.D ;
  assign WX4728 = \DFF_710.Q ;
  assign WX4729 = \DFF_711.D ;
  assign WX4730 = \DFF_711.Q ;
  assign WX4731 = \DFF_712.D ;
  assign WX4732 = \DFF_712.Q ;
  assign WX4733 = \DFF_713.D ;
  assign WX4734 = \DFF_713.Q ;
  assign WX4735 = \DFF_714.D ;
  assign WX4736 = \DFF_714.Q ;
  assign WX4737 = \DFF_715.D ;
  assign WX4738 = \DFF_715.Q ;
  assign WX4739 = \DFF_716.D ;
  assign WX4740 = \DFF_716.Q ;
  assign WX4741 = \DFF_717.D ;
  assign WX4742 = \DFF_717.Q ;
  assign WX4743 = \DFF_718.D ;
  assign WX4744 = \DFF_718.Q ;
  assign WX4745 = \DFF_719.D ;
  assign WX4746 = \DFF_719.Q ;
  assign WX4747 = \DFF_720.D ;
  assign WX4748 = \DFF_720.Q ;
  assign WX4749 = \DFF_721.D ;
  assign WX4750 = \DFF_721.Q ;
  assign WX4751 = \DFF_722.D ;
  assign WX4752 = \DFF_722.Q ;
  assign WX4753 = \DFF_723.D ;
  assign WX4754 = \DFF_723.Q ;
  assign WX4755 = \DFF_724.D ;
  assign WX4756 = \DFF_724.Q ;
  assign WX4757 = \DFF_725.D ;
  assign WX4758 = \DFF_725.Q ;
  assign WX4759 = \DFF_726.D ;
  assign WX4760 = \DFF_726.Q ;
  assign WX4761 = \DFF_727.D ;
  assign WX4762 = \DFF_727.Q ;
  assign WX4763 = \DFF_728.D ;
  assign WX4764 = \DFF_728.Q ;
  assign WX4765 = \DFF_729.D ;
  assign WX4766 = \DFF_729.Q ;
  assign WX4767 = \DFF_730.D ;
  assign WX4768 = \DFF_730.Q ;
  assign WX4769 = \DFF_731.D ;
  assign WX4770 = \DFF_731.Q ;
  assign WX4771 = \DFF_732.D ;
  assign WX4772 = \DFF_732.Q ;
  assign WX4773 = \DFF_733.D ;
  assign WX4774 = \DFF_733.Q ;
  assign WX4775 = \DFF_734.D ;
  assign WX4776 = \DFF_734.Q ;
  assign WX4777 = \DFF_735.D ;
  assign WX4778 = \DFF_735.Q ;
  assign WX484 = \DFF_0.D ;
  assign WX485 = \DFF_0.Q ;
  assign WX486 = \DFF_1.D ;
  assign WX487 = \DFF_1.Q ;
  assign WX488 = \DFF_2.D ;
  assign WX4880 = TM1;
  assign WX4881 = TM0;
  assign WX4882 = TM1;
  assign WX4883 = TM0;
  assign WX4884 = TM0;
  assign WX489 = \DFF_2.Q ;
  assign WX490 = \DFF_3.D ;
  assign WX491 = \DFF_3.Q ;
  assign WX492 = \DFF_4.D ;
  assign WX493 = \DFF_4.Q ;
  assign WX494 = \DFF_5.D ;
  assign WX495 = \DFF_5.Q ;
  assign WX496 = \DFF_6.D ;
  assign WX497 = \DFF_6.Q ;
  assign WX498 = \DFF_7.D ;
  assign WX499 = \DFF_7.Q ;
  assign WX500 = \DFF_8.D ;
  assign WX501 = \DFF_8.Q ;
  assign WX502 = \DFF_9.D ;
  assign WX503 = \DFF_9.Q ;
  assign WX504 = \DFF_10.D ;
  assign WX505 = \DFF_10.Q ;
  assign WX506 = \DFF_11.D ;
  assign WX507 = \DFF_11.Q ;
  assign WX508 = \DFF_12.D ;
  assign WX509 = \DFF_12.Q ;
  assign WX510 = \DFF_13.D ;
  assign WX511 = \DFF_13.Q ;
  assign WX512 = \DFF_14.D ;
  assign WX513 = \DFF_14.Q ;
  assign WX514 = \DFF_15.D ;
  assign WX5142 = RESET;
  assign WX5143 = \DFF_736.D ;
  assign WX5145 = \DFF_737.D ;
  assign WX5147 = \DFF_738.D ;
  assign WX5149 = \DFF_739.D ;
  assign WX515 = \DFF_15.Q ;
  assign WX5151 = \DFF_740.D ;
  assign WX5153 = \DFF_741.D ;
  assign WX5155 = \DFF_742.D ;
  assign WX5157 = \DFF_743.D ;
  assign WX5159 = \DFF_744.D ;
  assign WX516 = \DFF_16.D ;
  assign WX5161 = \DFF_745.D ;
  assign WX5163 = \DFF_746.D ;
  assign WX5165 = \DFF_747.D ;
  assign WX5167 = \DFF_748.D ;
  assign WX5169 = \DFF_749.D ;
  assign WX517 = \DFF_16.Q ;
  assign WX5171 = \DFF_750.D ;
  assign WX5173 = \DFF_751.D ;
  assign WX5175 = \DFF_752.D ;
  assign WX5177 = \DFF_753.D ;
  assign WX5179 = \DFF_754.D ;
  assign WX518 = \DFF_17.D ;
  assign WX5181 = \DFF_755.D ;
  assign WX5183 = \DFF_756.D ;
  assign WX5185 = \DFF_757.D ;
  assign WX5187 = \DFF_758.D ;
  assign WX5189 = \DFF_759.D ;
  assign WX519 = \DFF_17.Q ;
  assign WX5191 = \DFF_760.D ;
  assign WX5193 = \DFF_761.D ;
  assign WX5195 = \DFF_762.D ;
  assign WX5197 = \DFF_763.D ;
  assign WX5199 = \DFF_764.D ;
  assign WX520 = \DFF_18.D ;
  assign WX5201 = \DFF_765.D ;
  assign WX5203 = \DFF_766.D ;
  assign WX5205 = \DFF_767.D ;
  assign WX521 = \DFF_18.Q ;
  assign WX522 = \DFF_19.D ;
  assign WX523 = \DFF_19.Q ;
  assign WX524 = \DFF_20.D ;
  assign WX525 = \DFF_20.Q ;
  assign WX526 = \DFF_21.D ;
  assign WX527 = \DFF_21.Q ;
  assign WX528 = \DFF_22.D ;
  assign WX529 = \DFF_22.Q ;
  assign WX530 = \DFF_23.D ;
  assign WX531 = \DFF_23.Q ;
  assign WX532 = \DFF_24.D ;
  assign WX533 = \DFF_24.Q ;
  assign WX534 = \DFF_25.D ;
  assign WX535 = \DFF_25.Q ;
  assign WX536 = \DFF_26.D ;
  assign WX537 = \DFF_26.Q ;
  assign WX538 = \DFF_27.D ;
  assign WX539 = \DFF_27.Q ;
  assign WX540 = \DFF_28.D ;
  assign WX541 = \DFF_28.Q ;
  assign WX542 = \DFF_29.D ;
  assign WX543 = \DFF_29.Q ;
  assign WX544 = \DFF_30.D ;
  assign WX545 = \DFF_30.Q ;
  assign WX546 = \DFF_31.D ;
  assign WX547 = \DFF_31.Q ;
  assign WX5656 = \DFF_768.D ;
  assign WX5657 = \DFF_768.Q ;
  assign WX5658 = \DFF_769.D ;
  assign WX5659 = \DFF_769.Q ;
  assign WX5660 = \DFF_770.D ;
  assign WX5661 = \DFF_770.Q ;
  assign WX5662 = \DFF_771.D ;
  assign WX5663 = \DFF_771.Q ;
  assign WX5664 = \DFF_772.D ;
  assign WX5665 = \DFF_772.Q ;
  assign WX5666 = \DFF_773.D ;
  assign WX5667 = \DFF_773.Q ;
  assign WX5668 = \DFF_774.D ;
  assign WX5669 = \DFF_774.Q ;
  assign WX5670 = \DFF_775.D ;
  assign WX5671 = \DFF_775.Q ;
  assign WX5672 = \DFF_776.D ;
  assign WX5673 = \DFF_776.Q ;
  assign WX5674 = \DFF_777.D ;
  assign WX5675 = \DFF_777.Q ;
  assign WX5676 = \DFF_778.D ;
  assign WX5677 = \DFF_778.Q ;
  assign WX5678 = \DFF_779.D ;
  assign WX5679 = \DFF_779.Q ;
  assign WX5680 = \DFF_780.D ;
  assign WX5681 = \DFF_780.Q ;
  assign WX5682 = \DFF_781.D ;
  assign WX5683 = \DFF_781.Q ;
  assign WX5684 = \DFF_782.D ;
  assign WX5685 = \DFF_782.Q ;
  assign WX5686 = \DFF_783.D ;
  assign WX5687 = \DFF_783.Q ;
  assign WX5688 = \DFF_784.D ;
  assign WX5689 = \DFF_784.Q ;
  assign WX5690 = \DFF_785.D ;
  assign WX5691 = \DFF_785.Q ;
  assign WX5692 = \DFF_786.D ;
  assign WX5693 = \DFF_786.Q ;
  assign WX5694 = \DFF_787.D ;
  assign WX5695 = \DFF_787.Q ;
  assign WX5696 = \DFF_788.D ;
  assign WX5697 = \DFF_788.Q ;
  assign WX5698 = \DFF_789.D ;
  assign WX5699 = \DFF_789.Q ;
  assign WX5700 = \DFF_790.D ;
  assign WX5701 = \DFF_790.Q ;
  assign WX5702 = \DFF_791.D ;
  assign WX5703 = \DFF_791.Q ;
  assign WX5704 = \DFF_792.D ;
  assign WX5705 = \DFF_792.Q ;
  assign WX5706 = \DFF_793.D ;
  assign WX5707 = \DFF_793.Q ;
  assign WX5708 = \DFF_794.D ;
  assign WX5709 = \DFF_794.Q ;
  assign WX5710 = \DFF_795.D ;
  assign WX5711 = \DFF_795.Q ;
  assign WX5712 = \DFF_796.D ;
  assign WX5713 = \DFF_796.Q ;
  assign WX5714 = \DFF_797.D ;
  assign WX5715 = \DFF_797.Q ;
  assign WX5716 = \DFF_798.D ;
  assign WX5717 = \DFF_798.Q ;
  assign WX5718 = \DFF_799.D ;
  assign WX5719 = \DFF_799.Q ;
  assign WX5816 = \DFF_800.D ;
  assign WX5817 = \DFF_800.Q ;
  assign WX5818 = \DFF_801.D ;
  assign WX5819 = \DFF_801.Q ;
  assign WX5820 = \DFF_802.D ;
  assign WX5821 = \DFF_802.Q ;
  assign WX5822 = \DFF_803.D ;
  assign WX5823 = \DFF_803.Q ;
  assign WX5824 = \DFF_804.D ;
  assign WX5825 = \DFF_804.Q ;
  assign WX5826 = \DFF_805.D ;
  assign WX5827 = \DFF_805.Q ;
  assign WX5828 = \DFF_806.D ;
  assign WX5829 = \DFF_806.Q ;
  assign WX5830 = \DFF_807.D ;
  assign WX5831 = \DFF_807.Q ;
  assign WX5832 = \DFF_808.D ;
  assign WX5833 = \DFF_808.Q ;
  assign WX5834 = \DFF_809.D ;
  assign WX5835 = \DFF_809.Q ;
  assign WX5836 = \DFF_810.D ;
  assign WX5837 = \DFF_810.Q ;
  assign WX5838 = \DFF_811.D ;
  assign WX5839 = \DFF_811.Q ;
  assign WX5840 = \DFF_812.D ;
  assign WX5841 = \DFF_812.Q ;
  assign WX5842 = \DFF_813.D ;
  assign WX5843 = \DFF_813.Q ;
  assign WX5844 = \DFF_814.D ;
  assign WX5845 = \DFF_814.Q ;
  assign WX5846 = \DFF_815.D ;
  assign WX5847 = \DFF_815.Q ;
  assign WX5848 = \DFF_816.D ;
  assign WX5849 = \DFF_816.Q ;
  assign WX5850 = \DFF_817.D ;
  assign WX5851 = \DFF_817.Q ;
  assign WX5852 = \DFF_818.D ;
  assign WX5853 = \DFF_818.Q ;
  assign WX5854 = \DFF_819.D ;
  assign WX5855 = \DFF_819.Q ;
  assign WX5856 = \DFF_820.D ;
  assign WX5857 = \DFF_820.Q ;
  assign WX5858 = \DFF_821.D ;
  assign WX5859 = \DFF_821.Q ;
  assign WX5860 = \DFF_822.D ;
  assign WX5861 = \DFF_822.Q ;
  assign WX5862 = \DFF_823.D ;
  assign WX5863 = \DFF_823.Q ;
  assign WX5864 = \DFF_824.D ;
  assign WX5865 = \DFF_824.Q ;
  assign WX5866 = \DFF_825.D ;
  assign WX5867 = \DFF_825.Q ;
  assign WX5868 = \DFF_826.D ;
  assign WX5869 = \DFF_826.Q ;
  assign WX5870 = \DFF_827.D ;
  assign WX5871 = \DFF_827.Q ;
  assign WX5872 = \DFF_828.D ;
  assign WX5873 = \DFF_828.Q ;
  assign WX5874 = \DFF_829.D ;
  assign WX5875 = \DFF_829.Q ;
  assign WX5876 = \DFF_830.D ;
  assign WX5877 = \DFF_830.Q ;
  assign WX5878 = \DFF_831.D ;
  assign WX5879 = \DFF_831.Q ;
  assign WX5880 = \DFF_832.D ;
  assign WX5881 = \DFF_832.Q ;
  assign WX5882 = \DFF_833.D ;
  assign WX5883 = \DFF_833.Q ;
  assign WX5884 = \DFF_834.D ;
  assign WX5885 = \DFF_834.Q ;
  assign WX5886 = \DFF_835.D ;
  assign WX5887 = \DFF_835.Q ;
  assign WX5888 = \DFF_836.D ;
  assign WX5889 = \DFF_836.Q ;
  assign WX5890 = \DFF_837.D ;
  assign WX5891 = \DFF_837.Q ;
  assign WX5892 = \DFF_838.D ;
  assign WX5893 = \DFF_838.Q ;
  assign WX5894 = \DFF_839.D ;
  assign WX5895 = \DFF_839.Q ;
  assign WX5896 = \DFF_840.D ;
  assign WX5897 = \DFF_840.Q ;
  assign WX5898 = \DFF_841.D ;
  assign WX5899 = \DFF_841.Q ;
  assign WX5900 = \DFF_842.D ;
  assign WX5901 = \DFF_842.Q ;
  assign WX5902 = \DFF_843.D ;
  assign WX5903 = \DFF_843.Q ;
  assign WX5904 = \DFF_844.D ;
  assign WX5905 = \DFF_844.Q ;
  assign WX5906 = \DFF_845.D ;
  assign WX5907 = \DFF_845.Q ;
  assign WX5908 = \DFF_846.D ;
  assign WX5909 = \DFF_846.Q ;
  assign WX5910 = \DFF_847.D ;
  assign WX5911 = \DFF_847.Q ;
  assign WX5912 = \DFF_848.D ;
  assign WX5913 = \DFF_848.Q ;
  assign WX5914 = \DFF_849.D ;
  assign WX5915 = \DFF_849.Q ;
  assign WX5916 = \DFF_850.D ;
  assign WX5917 = \DFF_850.Q ;
  assign WX5918 = \DFF_851.D ;
  assign WX5919 = \DFF_851.Q ;
  assign WX5920 = \DFF_852.D ;
  assign WX5921 = \DFF_852.Q ;
  assign WX5922 = \DFF_853.D ;
  assign WX5923 = \DFF_853.Q ;
  assign WX5924 = \DFF_854.D ;
  assign WX5925 = \DFF_854.Q ;
  assign WX5926 = \DFF_855.D ;
  assign WX5927 = \DFF_855.Q ;
  assign WX5928 = \DFF_856.D ;
  assign WX5929 = \DFF_856.Q ;
  assign WX5930 = \DFF_857.D ;
  assign WX5931 = \DFF_857.Q ;
  assign WX5932 = \DFF_858.D ;
  assign WX5933 = \DFF_858.Q ;
  assign WX5934 = \DFF_859.D ;
  assign WX5935 = \DFF_859.Q ;
  assign WX5936 = \DFF_860.D ;
  assign WX5937 = \DFF_860.Q ;
  assign WX5938 = \DFF_861.D ;
  assign WX5939 = \DFF_861.Q ;
  assign WX5940 = \DFF_862.D ;
  assign WX5941 = \DFF_862.Q ;
  assign WX5942 = \DFF_863.D ;
  assign WX5943 = \DFF_863.Q ;
  assign WX5944 = \DFF_864.D ;
  assign WX5945 = \DFF_864.Q ;
  assign WX5946 = \DFF_865.D ;
  assign WX5947 = \DFF_865.Q ;
  assign WX5948 = \DFF_866.D ;
  assign WX5949 = \DFF_866.Q ;
  assign WX5950 = \DFF_867.D ;
  assign WX5951 = \DFF_867.Q ;
  assign WX5952 = \DFF_868.D ;
  assign WX5953 = \DFF_868.Q ;
  assign WX5954 = \DFF_869.D ;
  assign WX5955 = \DFF_869.Q ;
  assign WX5956 = \DFF_870.D ;
  assign WX5957 = \DFF_870.Q ;
  assign WX5958 = \DFF_871.D ;
  assign WX5959 = \DFF_871.Q ;
  assign WX5960 = \DFF_872.D ;
  assign WX5961 = \DFF_872.Q ;
  assign WX5962 = \DFF_873.D ;
  assign WX5963 = \DFF_873.Q ;
  assign WX5964 = \DFF_874.D ;
  assign WX5965 = \DFF_874.Q ;
  assign WX5966 = \DFF_875.D ;
  assign WX5967 = \DFF_875.Q ;
  assign WX5968 = \DFF_876.D ;
  assign WX5969 = \DFF_876.Q ;
  assign WX5970 = \DFF_877.D ;
  assign WX5971 = \DFF_877.Q ;
  assign WX5972 = \DFF_878.D ;
  assign WX5973 = \DFF_878.Q ;
  assign WX5974 = \DFF_879.D ;
  assign WX5975 = \DFF_879.Q ;
  assign WX5976 = \DFF_880.D ;
  assign WX5977 = \DFF_880.Q ;
  assign WX5978 = \DFF_881.D ;
  assign WX5979 = \DFF_881.Q ;
  assign WX5980 = \DFF_882.D ;
  assign WX5981 = \DFF_882.Q ;
  assign WX5982 = \DFF_883.D ;
  assign WX5983 = \DFF_883.Q ;
  assign WX5984 = \DFF_884.D ;
  assign WX5985 = \DFF_884.Q ;
  assign WX5986 = \DFF_885.D ;
  assign WX5987 = \DFF_885.Q ;
  assign WX5988 = \DFF_886.D ;
  assign WX5989 = \DFF_886.Q ;
  assign WX5990 = \DFF_887.D ;
  assign WX5991 = \DFF_887.Q ;
  assign WX5992 = \DFF_888.D ;
  assign WX5993 = \DFF_888.Q ;
  assign WX5994 = \DFF_889.D ;
  assign WX5995 = \DFF_889.Q ;
  assign WX5996 = \DFF_890.D ;
  assign WX5997 = \DFF_890.Q ;
  assign WX5998 = \DFF_891.D ;
  assign WX5999 = \DFF_891.Q ;
  assign WX6000 = \DFF_892.D ;
  assign WX6001 = \DFF_892.Q ;
  assign WX6002 = \DFF_893.D ;
  assign WX6003 = \DFF_893.Q ;
  assign WX6004 = \DFF_894.D ;
  assign WX6005 = \DFF_894.Q ;
  assign WX6006 = \DFF_895.D ;
  assign WX6007 = \DFF_895.Q ;
  assign WX6008 = \DFF_896.D ;
  assign WX6009 = \DFF_896.Q ;
  assign WX6010 = \DFF_897.D ;
  assign WX6011 = \DFF_897.Q ;
  assign WX6012 = \DFF_898.D ;
  assign WX6013 = \DFF_898.Q ;
  assign WX6014 = \DFF_899.D ;
  assign WX6015 = \DFF_899.Q ;
  assign WX6016 = \DFF_900.D ;
  assign WX6017 = \DFF_900.Q ;
  assign WX6018 = \DFF_901.D ;
  assign WX6019 = \DFF_901.Q ;
  assign WX6020 = \DFF_902.D ;
  assign WX6021 = \DFF_902.Q ;
  assign WX6022 = \DFF_903.D ;
  assign WX6023 = \DFF_903.Q ;
  assign WX6024 = \DFF_904.D ;
  assign WX6025 = \DFF_904.Q ;
  assign WX6026 = \DFF_905.D ;
  assign WX6027 = \DFF_905.Q ;
  assign WX6028 = \DFF_906.D ;
  assign WX6029 = \DFF_906.Q ;
  assign WX6030 = \DFF_907.D ;
  assign WX6031 = \DFF_907.Q ;
  assign WX6032 = \DFF_908.D ;
  assign WX6033 = \DFF_908.Q ;
  assign WX6034 = \DFF_909.D ;
  assign WX6035 = \DFF_909.Q ;
  assign WX6036 = \DFF_910.D ;
  assign WX6037 = \DFF_910.Q ;
  assign WX6038 = \DFF_911.D ;
  assign WX6039 = \DFF_911.Q ;
  assign WX6040 = \DFF_912.D ;
  assign WX6041 = \DFF_912.Q ;
  assign WX6042 = \DFF_913.D ;
  assign WX6043 = \DFF_913.Q ;
  assign WX6044 = \DFF_914.D ;
  assign WX6045 = \DFF_914.Q ;
  assign WX6046 = \DFF_915.D ;
  assign WX6047 = \DFF_915.Q ;
  assign WX6048 = \DFF_916.D ;
  assign WX6049 = \DFF_916.Q ;
  assign WX6050 = \DFF_917.D ;
  assign WX6051 = \DFF_917.Q ;
  assign WX6052 = \DFF_918.D ;
  assign WX6053 = \DFF_918.Q ;
  assign WX6054 = \DFF_919.D ;
  assign WX6055 = \DFF_919.Q ;
  assign WX6056 = \DFF_920.D ;
  assign WX6057 = \DFF_920.Q ;
  assign WX6058 = \DFF_921.D ;
  assign WX6059 = \DFF_921.Q ;
  assign WX6060 = \DFF_922.D ;
  assign WX6061 = \DFF_922.Q ;
  assign WX6062 = \DFF_923.D ;
  assign WX6063 = \DFF_923.Q ;
  assign WX6064 = \DFF_924.D ;
  assign WX6065 = \DFF_924.Q ;
  assign WX6066 = \DFF_925.D ;
  assign WX6067 = \DFF_925.Q ;
  assign WX6068 = \DFF_926.D ;
  assign WX6069 = \DFF_926.Q ;
  assign WX6070 = \DFF_927.D ;
  assign WX6071 = \DFF_927.Q ;
  assign WX6173 = TM1;
  assign WX6174 = TM0;
  assign WX6175 = TM1;
  assign WX6176 = TM0;
  assign WX6177 = TM0;
  assign WX6435 = RESET;
  assign WX6436 = \DFF_928.D ;
  assign WX6438 = \DFF_929.D ;
  assign WX644 = \DFF_32.D ;
  assign WX6440 = \DFF_930.D ;
  assign WX6442 = \DFF_931.D ;
  assign WX6444 = \DFF_932.D ;
  assign WX6446 = \DFF_933.D ;
  assign WX6448 = \DFF_934.D ;
  assign WX645 = \DFF_32.Q ;
  assign WX6450 = \DFF_935.D ;
  assign WX6452 = \DFF_936.D ;
  assign WX6454 = \DFF_937.D ;
  assign WX6456 = \DFF_938.D ;
  assign WX6458 = \DFF_939.D ;
  assign WX646 = \DFF_33.D ;
  assign WX6460 = \DFF_940.D ;
  assign WX6462 = \DFF_941.D ;
  assign WX6464 = \DFF_942.D ;
  assign WX6466 = \DFF_943.D ;
  assign WX6468 = \DFF_944.D ;
  assign WX647 = \DFF_33.Q ;
  assign WX6470 = \DFF_945.D ;
  assign WX6472 = \DFF_946.D ;
  assign WX6474 = \DFF_947.D ;
  assign WX6476 = \DFF_948.D ;
  assign WX6478 = \DFF_949.D ;
  assign WX648 = \DFF_34.D ;
  assign WX6480 = \DFF_950.D ;
  assign WX6482 = \DFF_951.D ;
  assign WX6484 = \DFF_952.D ;
  assign WX6486 = \DFF_953.D ;
  assign WX6488 = \DFF_954.D ;
  assign WX649 = \DFF_34.Q ;
  assign WX6490 = \DFF_955.D ;
  assign WX6492 = \DFF_956.D ;
  assign WX6494 = \DFF_957.D ;
  assign WX6496 = \DFF_958.D ;
  assign WX6498 = \DFF_959.D ;
  assign WX650 = \DFF_35.D ;
  assign WX651 = \DFF_35.Q ;
  assign WX652 = \DFF_36.D ;
  assign WX653 = \DFF_36.Q ;
  assign WX654 = \DFF_37.D ;
  assign WX655 = \DFF_37.Q ;
  assign WX656 = \DFF_38.D ;
  assign WX657 = \DFF_38.Q ;
  assign WX658 = \DFF_39.D ;
  assign WX659 = \DFF_39.Q ;
  assign WX660 = \DFF_40.D ;
  assign WX661 = \DFF_40.Q ;
  assign WX662 = \DFF_41.D ;
  assign WX663 = \DFF_41.Q ;
  assign WX664 = \DFF_42.D ;
  assign WX665 = \DFF_42.Q ;
  assign WX666 = \DFF_43.D ;
  assign WX667 = \DFF_43.Q ;
  assign WX668 = \DFF_44.D ;
  assign WX669 = \DFF_44.Q ;
  assign WX670 = \DFF_45.D ;
  assign WX671 = \DFF_45.Q ;
  assign WX672 = \DFF_46.D ;
  assign WX673 = \DFF_46.Q ;
  assign WX674 = \DFF_47.D ;
  assign WX675 = \DFF_47.Q ;
  assign WX676 = \DFF_48.D ;
  assign WX677 = \DFF_48.Q ;
  assign WX678 = \DFF_49.D ;
  assign WX679 = \DFF_49.Q ;
  assign WX680 = \DFF_50.D ;
  assign WX681 = \DFF_50.Q ;
  assign WX682 = \DFF_51.D ;
  assign WX683 = \DFF_51.Q ;
  assign WX684 = \DFF_52.D ;
  assign WX685 = \DFF_52.Q ;
  assign WX686 = \DFF_53.D ;
  assign WX687 = \DFF_53.Q ;
  assign WX688 = \DFF_54.D ;
  assign WX689 = \DFF_54.Q ;
  assign WX690 = \DFF_55.D ;
  assign WX691 = \DFF_55.Q ;
  assign WX692 = \DFF_56.D ;
  assign WX693 = \DFF_56.Q ;
  assign WX694 = \DFF_57.D ;
  assign WX6949 = \DFF_960.D ;
  assign WX695 = \DFF_57.Q ;
  assign WX6950 = \DFF_960.Q ;
  assign WX6951 = \DFF_961.D ;
  assign WX6952 = \DFF_961.Q ;
  assign WX6953 = \DFF_962.D ;
  assign WX6954 = \DFF_962.Q ;
  assign WX6955 = \DFF_963.D ;
  assign WX6956 = \DFF_963.Q ;
  assign WX6957 = \DFF_964.D ;
  assign WX6958 = \DFF_964.Q ;
  assign WX6959 = \DFF_965.D ;
  assign WX696 = \DFF_58.D ;
  assign WX6960 = \DFF_965.Q ;
  assign WX6961 = \DFF_966.D ;
  assign WX6962 = \DFF_966.Q ;
  assign WX6963 = \DFF_967.D ;
  assign WX6964 = \DFF_967.Q ;
  assign WX6965 = \DFF_968.D ;
  assign WX6966 = \DFF_968.Q ;
  assign WX6967 = \DFF_969.D ;
  assign WX6968 = \DFF_969.Q ;
  assign WX6969 = \DFF_970.D ;
  assign WX697 = \DFF_58.Q ;
  assign WX6970 = \DFF_970.Q ;
  assign WX6971 = \DFF_971.D ;
  assign WX6972 = \DFF_971.Q ;
  assign WX6973 = \DFF_972.D ;
  assign WX6974 = \DFF_972.Q ;
  assign WX6975 = \DFF_973.D ;
  assign WX6976 = \DFF_973.Q ;
  assign WX6977 = \DFF_974.D ;
  assign WX6978 = \DFF_974.Q ;
  assign WX6979 = \DFF_975.D ;
  assign WX698 = \DFF_59.D ;
  assign WX6980 = \DFF_975.Q ;
  assign WX6981 = \DFF_976.D ;
  assign WX6982 = \DFF_976.Q ;
  assign WX6983 = \DFF_977.D ;
  assign WX6984 = \DFF_977.Q ;
  assign WX6985 = \DFF_978.D ;
  assign WX6986 = \DFF_978.Q ;
  assign WX6987 = \DFF_979.D ;
  assign WX6988 = \DFF_979.Q ;
  assign WX6989 = \DFF_980.D ;
  assign WX699 = \DFF_59.Q ;
  assign WX6990 = \DFF_980.Q ;
  assign WX6991 = \DFF_981.D ;
  assign WX6992 = \DFF_981.Q ;
  assign WX6993 = \DFF_982.D ;
  assign WX6994 = \DFF_982.Q ;
  assign WX6995 = \DFF_983.D ;
  assign WX6996 = \DFF_983.Q ;
  assign WX6997 = \DFF_984.D ;
  assign WX6998 = \DFF_984.Q ;
  assign WX6999 = \DFF_985.D ;
  assign WX700 = \DFF_60.D ;
  assign WX7000 = \DFF_985.Q ;
  assign WX7001 = \DFF_986.D ;
  assign WX7002 = \DFF_986.Q ;
  assign WX7003 = \DFF_987.D ;
  assign WX7004 = \DFF_987.Q ;
  assign WX7005 = \DFF_988.D ;
  assign WX7006 = \DFF_988.Q ;
  assign WX7007 = \DFF_989.D ;
  assign WX7008 = \DFF_989.Q ;
  assign WX7009 = \DFF_990.D ;
  assign WX701 = \DFF_60.Q ;
  assign WX7010 = \DFF_990.Q ;
  assign WX7011 = \DFF_991.D ;
  assign WX7012 = \DFF_991.Q ;
  assign WX702 = \DFF_61.D ;
  assign WX703 = \DFF_61.Q ;
  assign WX704 = \DFF_62.D ;
  assign WX705 = \DFF_62.Q ;
  assign WX706 = \DFF_63.D ;
  assign WX707 = \DFF_63.Q ;
  assign WX708 = \DFF_64.D ;
  assign WX709 = \DFF_64.Q ;
  assign WX710 = \DFF_65.D ;
  assign WX7109 = \DFF_992.D ;
  assign WX711 = \DFF_65.Q ;
  assign WX7110 = \DFF_992.Q ;
  assign WX7111 = \DFF_993.D ;
  assign WX7112 = \DFF_993.Q ;
  assign WX7113 = \DFF_994.D ;
  assign WX7114 = \DFF_994.Q ;
  assign WX7115 = \DFF_995.D ;
  assign WX7116 = \DFF_995.Q ;
  assign WX7117 = \DFF_996.D ;
  assign WX7118 = \DFF_996.Q ;
  assign WX7119 = \DFF_997.D ;
  assign WX712 = \DFF_66.D ;
  assign WX7120 = \DFF_997.Q ;
  assign WX7121 = \DFF_998.D ;
  assign WX7122 = \DFF_998.Q ;
  assign WX7123 = \DFF_999.D ;
  assign WX7124 = \DFF_999.Q ;
  assign WX7125 = \DFF_1000.D ;
  assign WX7126 = \DFF_1000.Q ;
  assign WX7127 = \DFF_1001.D ;
  assign WX7128 = \DFF_1001.Q ;
  assign WX7129 = \DFF_1002.D ;
  assign WX713 = \DFF_66.Q ;
  assign WX7130 = \DFF_1002.Q ;
  assign WX7131 = \DFF_1003.D ;
  assign WX7132 = \DFF_1003.Q ;
  assign WX7133 = \DFF_1004.D ;
  assign WX7134 = \DFF_1004.Q ;
  assign WX7135 = \DFF_1005.D ;
  assign WX7136 = \DFF_1005.Q ;
  assign WX7137 = \DFF_1006.D ;
  assign WX7138 = \DFF_1006.Q ;
  assign WX7139 = \DFF_1007.D ;
  assign WX714 = \DFF_67.D ;
  assign WX7140 = \DFF_1007.Q ;
  assign WX7141 = \DFF_1008.D ;
  assign WX7142 = \DFF_1008.Q ;
  assign WX7143 = \DFF_1009.D ;
  assign WX7144 = \DFF_1009.Q ;
  assign WX7145 = \DFF_1010.D ;
  assign WX7146 = \DFF_1010.Q ;
  assign WX7147 = \DFF_1011.D ;
  assign WX7148 = \DFF_1011.Q ;
  assign WX7149 = \DFF_1012.D ;
  assign WX715 = \DFF_67.Q ;
  assign WX7150 = \DFF_1012.Q ;
  assign WX7151 = \DFF_1013.D ;
  assign WX7152 = \DFF_1013.Q ;
  assign WX7153 = \DFF_1014.D ;
  assign WX7154 = \DFF_1014.Q ;
  assign WX7155 = \DFF_1015.D ;
  assign WX7156 = \DFF_1015.Q ;
  assign WX7157 = \DFF_1016.D ;
  assign WX7158 = \DFF_1016.Q ;
  assign WX7159 = \DFF_1017.D ;
  assign WX716 = \DFF_68.D ;
  assign WX7160 = \DFF_1017.Q ;
  assign WX7161 = \DFF_1018.D ;
  assign WX7162 = \DFF_1018.Q ;
  assign WX7163 = \DFF_1019.D ;
  assign WX7164 = \DFF_1019.Q ;
  assign WX7165 = \DFF_1020.D ;
  assign WX7166 = \DFF_1020.Q ;
  assign WX7167 = \DFF_1021.D ;
  assign WX7168 = \DFF_1021.Q ;
  assign WX7169 = \DFF_1022.D ;
  assign WX717 = \DFF_68.Q ;
  assign WX7170 = \DFF_1022.Q ;
  assign WX7171 = \DFF_1023.D ;
  assign WX7172 = \DFF_1023.Q ;
  assign WX7173 = \DFF_1024.D ;
  assign WX7174 = \DFF_1024.Q ;
  assign WX7175 = \DFF_1025.D ;
  assign WX7176 = \DFF_1025.Q ;
  assign WX7177 = \DFF_1026.D ;
  assign WX7178 = \DFF_1026.Q ;
  assign WX7179 = \DFF_1027.D ;
  assign WX718 = \DFF_69.D ;
  assign WX7180 = \DFF_1027.Q ;
  assign WX7181 = \DFF_1028.D ;
  assign WX7182 = \DFF_1028.Q ;
  assign WX7183 = \DFF_1029.D ;
  assign WX7184 = \DFF_1029.Q ;
  assign WX7185 = \DFF_1030.D ;
  assign WX7186 = \DFF_1030.Q ;
  assign WX7187 = \DFF_1031.D ;
  assign WX7188 = \DFF_1031.Q ;
  assign WX7189 = \DFF_1032.D ;
  assign WX719 = \DFF_69.Q ;
  assign WX7190 = \DFF_1032.Q ;
  assign WX7191 = \DFF_1033.D ;
  assign WX7192 = \DFF_1033.Q ;
  assign WX7193 = \DFF_1034.D ;
  assign WX7194 = \DFF_1034.Q ;
  assign WX7195 = \DFF_1035.D ;
  assign WX7196 = \DFF_1035.Q ;
  assign WX7197 = \DFF_1036.D ;
  assign WX7198 = \DFF_1036.Q ;
  assign WX7199 = \DFF_1037.D ;
  assign WX720 = \DFF_70.D ;
  assign WX7200 = \DFF_1037.Q ;
  assign WX7201 = \DFF_1038.D ;
  assign WX7202 = \DFF_1038.Q ;
  assign WX7203 = \DFF_1039.D ;
  assign WX7204 = \DFF_1039.Q ;
  assign WX7205 = \DFF_1040.D ;
  assign WX7206 = \DFF_1040.Q ;
  assign WX7207 = \DFF_1041.D ;
  assign WX7208 = \DFF_1041.Q ;
  assign WX7209 = \DFF_1042.D ;
  assign WX721 = \DFF_70.Q ;
  assign WX7210 = \DFF_1042.Q ;
  assign WX7211 = \DFF_1043.D ;
  assign WX7212 = \DFF_1043.Q ;
  assign WX7213 = \DFF_1044.D ;
  assign WX7214 = \DFF_1044.Q ;
  assign WX7215 = \DFF_1045.D ;
  assign WX7216 = \DFF_1045.Q ;
  assign WX7217 = \DFF_1046.D ;
  assign WX7218 = \DFF_1046.Q ;
  assign WX7219 = \DFF_1047.D ;
  assign WX722 = \DFF_71.D ;
  assign WX7220 = \DFF_1047.Q ;
  assign WX7221 = \DFF_1048.D ;
  assign WX7222 = \DFF_1048.Q ;
  assign WX7223 = \DFF_1049.D ;
  assign WX7224 = \DFF_1049.Q ;
  assign WX7225 = \DFF_1050.D ;
  assign WX7226 = \DFF_1050.Q ;
  assign WX7227 = \DFF_1051.D ;
  assign WX7228 = \DFF_1051.Q ;
  assign WX7229 = \DFF_1052.D ;
  assign WX723 = \DFF_71.Q ;
  assign WX7230 = \DFF_1052.Q ;
  assign WX7231 = \DFF_1053.D ;
  assign WX7232 = \DFF_1053.Q ;
  assign WX7233 = \DFF_1054.D ;
  assign WX7234 = \DFF_1054.Q ;
  assign WX7235 = \DFF_1055.D ;
  assign WX7236 = \DFF_1055.Q ;
  assign WX7237 = \DFF_1056.D ;
  assign WX7238 = \DFF_1056.Q ;
  assign WX7239 = \DFF_1057.D ;
  assign WX724 = \DFF_72.D ;
  assign WX7240 = \DFF_1057.Q ;
  assign WX7241 = \DFF_1058.D ;
  assign WX7242 = \DFF_1058.Q ;
  assign WX7243 = \DFF_1059.D ;
  assign WX7244 = \DFF_1059.Q ;
  assign WX7245 = \DFF_1060.D ;
  assign WX7246 = \DFF_1060.Q ;
  assign WX7247 = \DFF_1061.D ;
  assign WX7248 = \DFF_1061.Q ;
  assign WX7249 = \DFF_1062.D ;
  assign WX725 = \DFF_72.Q ;
  assign WX7250 = \DFF_1062.Q ;
  assign WX7251 = \DFF_1063.D ;
  assign WX7252 = \DFF_1063.Q ;
  assign WX7253 = \DFF_1064.D ;
  assign WX7254 = \DFF_1064.Q ;
  assign WX7255 = \DFF_1065.D ;
  assign WX7256 = \DFF_1065.Q ;
  assign WX7257 = \DFF_1066.D ;
  assign WX7258 = \DFF_1066.Q ;
  assign WX7259 = \DFF_1067.D ;
  assign WX726 = \DFF_73.D ;
  assign WX7260 = \DFF_1067.Q ;
  assign WX7261 = \DFF_1068.D ;
  assign WX7262 = \DFF_1068.Q ;
  assign WX7263 = \DFF_1069.D ;
  assign WX7264 = \DFF_1069.Q ;
  assign WX7265 = \DFF_1070.D ;
  assign WX7266 = \DFF_1070.Q ;
  assign WX7267 = \DFF_1071.D ;
  assign WX7268 = \DFF_1071.Q ;
  assign WX7269 = \DFF_1072.D ;
  assign WX727 = \DFF_73.Q ;
  assign WX7270 = \DFF_1072.Q ;
  assign WX7271 = \DFF_1073.D ;
  assign WX7272 = \DFF_1073.Q ;
  assign WX7273 = \DFF_1074.D ;
  assign WX7274 = \DFF_1074.Q ;
  assign WX7275 = \DFF_1075.D ;
  assign WX7276 = \DFF_1075.Q ;
  assign WX7277 = \DFF_1076.D ;
  assign WX7278 = \DFF_1076.Q ;
  assign WX7279 = \DFF_1077.D ;
  assign WX728 = \DFF_74.D ;
  assign WX7280 = \DFF_1077.Q ;
  assign WX7281 = \DFF_1078.D ;
  assign WX7282 = \DFF_1078.Q ;
  assign WX7283 = \DFF_1079.D ;
  assign WX7284 = \DFF_1079.Q ;
  assign WX7285 = \DFF_1080.D ;
  assign WX7286 = \DFF_1080.Q ;
  assign WX7287 = \DFF_1081.D ;
  assign WX7288 = \DFF_1081.Q ;
  assign WX7289 = \DFF_1082.D ;
  assign WX729 = \DFF_74.Q ;
  assign WX7290 = \DFF_1082.Q ;
  assign WX7291 = \DFF_1083.D ;
  assign WX7292 = \DFF_1083.Q ;
  assign WX7293 = \DFF_1084.D ;
  assign WX7294 = \DFF_1084.Q ;
  assign WX7295 = \DFF_1085.D ;
  assign WX7296 = \DFF_1085.Q ;
  assign WX7297 = \DFF_1086.D ;
  assign WX7298 = \DFF_1086.Q ;
  assign WX7299 = \DFF_1087.D ;
  assign WX730 = \DFF_75.D ;
  assign WX7300 = \DFF_1087.Q ;
  assign WX7301 = \DFF_1088.D ;
  assign WX7302 = \DFF_1088.Q ;
  assign WX7303 = \DFF_1089.D ;
  assign WX7304 = \DFF_1089.Q ;
  assign WX7305 = \DFF_1090.D ;
  assign WX7306 = \DFF_1090.Q ;
  assign WX7307 = \DFF_1091.D ;
  assign WX7308 = \DFF_1091.Q ;
  assign WX7309 = \DFF_1092.D ;
  assign WX731 = \DFF_75.Q ;
  assign WX7310 = \DFF_1092.Q ;
  assign WX7311 = \DFF_1093.D ;
  assign WX7312 = \DFF_1093.Q ;
  assign WX7313 = \DFF_1094.D ;
  assign WX7314 = \DFF_1094.Q ;
  assign WX7315 = \DFF_1095.D ;
  assign WX7316 = \DFF_1095.Q ;
  assign WX7317 = \DFF_1096.D ;
  assign WX7318 = \DFF_1096.Q ;
  assign WX7319 = \DFF_1097.D ;
  assign WX732 = \DFF_76.D ;
  assign WX7320 = \DFF_1097.Q ;
  assign WX7321 = \DFF_1098.D ;
  assign WX7322 = \DFF_1098.Q ;
  assign WX7323 = \DFF_1099.D ;
  assign WX7324 = \DFF_1099.Q ;
  assign WX7325 = \DFF_1100.D ;
  assign WX7326 = \DFF_1100.Q ;
  assign WX7327 = \DFF_1101.D ;
  assign WX7328 = \DFF_1101.Q ;
  assign WX7329 = \DFF_1102.D ;
  assign WX733 = \DFF_76.Q ;
  assign WX7330 = \DFF_1102.Q ;
  assign WX7331 = \DFF_1103.D ;
  assign WX7332 = \DFF_1103.Q ;
  assign WX7333 = \DFF_1104.D ;
  assign WX7334 = \DFF_1104.Q ;
  assign WX7335 = \DFF_1105.D ;
  assign WX7336 = \DFF_1105.Q ;
  assign WX7337 = \DFF_1106.D ;
  assign WX7338 = \DFF_1106.Q ;
  assign WX7339 = \DFF_1107.D ;
  assign WX734 = \DFF_77.D ;
  assign WX7340 = \DFF_1107.Q ;
  assign WX7341 = \DFF_1108.D ;
  assign WX7342 = \DFF_1108.Q ;
  assign WX7343 = \DFF_1109.D ;
  assign WX7344 = \DFF_1109.Q ;
  assign WX7345 = \DFF_1110.D ;
  assign WX7346 = \DFF_1110.Q ;
  assign WX7347 = \DFF_1111.D ;
  assign WX7348 = \DFF_1111.Q ;
  assign WX7349 = \DFF_1112.D ;
  assign WX735 = \DFF_77.Q ;
  assign WX7350 = \DFF_1112.Q ;
  assign WX7351 = \DFF_1113.D ;
  assign WX7352 = \DFF_1113.Q ;
  assign WX7353 = \DFF_1114.D ;
  assign WX7354 = \DFF_1114.Q ;
  assign WX7355 = \DFF_1115.D ;
  assign WX7356 = \DFF_1115.Q ;
  assign WX7357 = \DFF_1116.D ;
  assign WX7358 = \DFF_1116.Q ;
  assign WX7359 = \DFF_1117.D ;
  assign WX736 = \DFF_78.D ;
  assign WX7360 = \DFF_1117.Q ;
  assign WX7361 = \DFF_1118.D ;
  assign WX7362 = \DFF_1118.Q ;
  assign WX7363 = \DFF_1119.D ;
  assign WX7364 = \DFF_1119.Q ;
  assign WX737 = \DFF_78.Q ;
  assign WX738 = \DFF_79.D ;
  assign WX739 = \DFF_79.Q ;
  assign WX740 = \DFF_80.D ;
  assign WX741 = \DFF_80.Q ;
  assign WX742 = \DFF_81.D ;
  assign WX743 = \DFF_81.Q ;
  assign WX744 = \DFF_82.D ;
  assign WX745 = \DFF_82.Q ;
  assign WX746 = \DFF_83.D ;
  assign WX7466 = TM1;
  assign WX7467 = TM0;
  assign WX7468 = TM1;
  assign WX7469 = TM0;
  assign WX747 = \DFF_83.Q ;
  assign WX7470 = TM0;
  assign WX748 = \DFF_84.D ;
  assign WX749 = \DFF_84.Q ;
  assign WX750 = \DFF_85.D ;
  assign WX751 = \DFF_85.Q ;
  assign WX752 = \DFF_86.D ;
  assign WX753 = \DFF_86.Q ;
  assign WX754 = \DFF_87.D ;
  assign WX755 = \DFF_87.Q ;
  assign WX756 = \DFF_88.D ;
  assign WX757 = \DFF_88.Q ;
  assign WX758 = \DFF_89.D ;
  assign WX759 = \DFF_89.Q ;
  assign WX760 = \DFF_90.D ;
  assign WX761 = \DFF_90.Q ;
  assign WX762 = \DFF_91.D ;
  assign WX763 = \DFF_91.Q ;
  assign WX764 = \DFF_92.D ;
  assign WX765 = \DFF_92.Q ;
  assign WX766 = \DFF_93.D ;
  assign WX767 = \DFF_93.Q ;
  assign WX768 = \DFF_94.D ;
  assign WX769 = \DFF_94.Q ;
  assign WX770 = \DFF_95.D ;
  assign WX771 = \DFF_95.Q ;
  assign WX772 = \DFF_96.D ;
  assign WX7728 = RESET;
  assign WX7729 = \DFF_1120.D ;
  assign WX773 = \DFF_96.Q ;
  assign WX7731 = \DFF_1121.D ;
  assign WX7733 = \DFF_1122.D ;
  assign WX7735 = \DFF_1123.D ;
  assign WX7737 = \DFF_1124.D ;
  assign WX7739 = \DFF_1125.D ;
  assign WX774 = \DFF_97.D ;
  assign WX7741 = \DFF_1126.D ;
  assign WX7743 = \DFF_1127.D ;
  assign WX7745 = \DFF_1128.D ;
  assign WX7747 = \DFF_1129.D ;
  assign WX7749 = \DFF_1130.D ;
  assign WX775 = \DFF_97.Q ;
  assign WX7751 = \DFF_1131.D ;
  assign WX7753 = \DFF_1132.D ;
  assign WX7755 = \DFF_1133.D ;
  assign WX7757 = \DFF_1134.D ;
  assign WX7759 = \DFF_1135.D ;
  assign WX776 = \DFF_98.D ;
  assign WX7761 = \DFF_1136.D ;
  assign WX7763 = \DFF_1137.D ;
  assign WX7765 = \DFF_1138.D ;
  assign WX7767 = \DFF_1139.D ;
  assign WX7769 = \DFF_1140.D ;
  assign WX777 = \DFF_98.Q ;
  assign WX7771 = \DFF_1141.D ;
  assign WX7773 = \DFF_1142.D ;
  assign WX7775 = \DFF_1143.D ;
  assign WX7777 = \DFF_1144.D ;
  assign WX7779 = \DFF_1145.D ;
  assign WX778 = \DFF_99.D ;
  assign WX7781 = \DFF_1146.D ;
  assign WX7783 = \DFF_1147.D ;
  assign WX7785 = \DFF_1148.D ;
  assign WX7787 = \DFF_1149.D ;
  assign WX7789 = \DFF_1150.D ;
  assign WX779 = \DFF_99.Q ;
  assign WX7791 = \DFF_1151.D ;
  assign WX780 = \DFF_100.D ;
  assign WX781 = \DFF_100.Q ;
  assign WX782 = \DFF_101.D ;
  assign WX783 = \DFF_101.Q ;
  assign WX784 = \DFF_102.D ;
  assign WX785 = \DFF_102.Q ;
  assign WX786 = \DFF_103.D ;
  assign WX787 = \DFF_103.Q ;
  assign WX788 = \DFF_104.D ;
  assign WX789 = \DFF_104.Q ;
  assign WX790 = \DFF_105.D ;
  assign WX791 = \DFF_105.Q ;
  assign WX792 = \DFF_106.D ;
  assign WX793 = \DFF_106.Q ;
  assign WX794 = \DFF_107.D ;
  assign WX795 = \DFF_107.Q ;
  assign WX796 = \DFF_108.D ;
  assign WX797 = \DFF_108.Q ;
  assign WX798 = \DFF_109.D ;
  assign WX799 = \DFF_109.Q ;
  assign WX800 = \DFF_110.D ;
  assign WX801 = \DFF_110.Q ;
  assign WX802 = \DFF_111.D ;
  assign WX803 = \DFF_111.Q ;
  assign WX804 = \DFF_112.D ;
  assign WX805 = \DFF_112.Q ;
  assign WX806 = \DFF_113.D ;
  assign WX807 = \DFF_113.Q ;
  assign WX808 = \DFF_114.D ;
  assign WX809 = \DFF_114.Q ;
  assign WX810 = \DFF_115.D ;
  assign WX811 = \DFF_115.Q ;
  assign WX812 = \DFF_116.D ;
  assign WX813 = \DFF_116.Q ;
  assign WX814 = \DFF_117.D ;
  assign WX815 = \DFF_117.Q ;
  assign WX816 = \DFF_118.D ;
  assign WX817 = \DFF_118.Q ;
  assign WX818 = \DFF_119.D ;
  assign WX819 = \DFF_119.Q ;
  assign WX820 = \DFF_120.D ;
  assign WX821 = \DFF_120.Q ;
  assign WX822 = \DFF_121.D ;
  assign WX823 = \DFF_121.Q ;
  assign WX824 = \DFF_122.D ;
  assign WX8242 = \DFF_1152.D ;
  assign WX8243 = \DFF_1152.Q ;
  assign WX8244 = \DFF_1153.D ;
  assign WX8245 = \DFF_1153.Q ;
  assign WX8246 = \DFF_1154.D ;
  assign WX8247 = \DFF_1154.Q ;
  assign WX8248 = \DFF_1155.D ;
  assign WX8249 = \DFF_1155.Q ;
  assign WX825 = \DFF_122.Q ;
  assign WX8250 = \DFF_1156.D ;
  assign WX8251 = \DFF_1156.Q ;
  assign WX8252 = \DFF_1157.D ;
  assign WX8253 = \DFF_1157.Q ;
  assign WX8254 = \DFF_1158.D ;
  assign WX8255 = \DFF_1158.Q ;
  assign WX8256 = \DFF_1159.D ;
  assign WX8257 = \DFF_1159.Q ;
  assign WX8258 = \DFF_1160.D ;
  assign WX8259 = \DFF_1160.Q ;
  assign WX826 = \DFF_123.D ;
  assign WX8260 = \DFF_1161.D ;
  assign WX8261 = \DFF_1161.Q ;
  assign WX8262 = \DFF_1162.D ;
  assign WX8263 = \DFF_1162.Q ;
  assign WX8264 = \DFF_1163.D ;
  assign WX8265 = \DFF_1163.Q ;
  assign WX8266 = \DFF_1164.D ;
  assign WX8267 = \DFF_1164.Q ;
  assign WX8268 = \DFF_1165.D ;
  assign WX8269 = \DFF_1165.Q ;
  assign WX827 = \DFF_123.Q ;
  assign WX8270 = \DFF_1166.D ;
  assign WX8271 = \DFF_1166.Q ;
  assign WX8272 = \DFF_1167.D ;
  assign WX8273 = \DFF_1167.Q ;
  assign WX8274 = \DFF_1168.D ;
  assign WX8275 = \DFF_1168.Q ;
  assign WX8276 = \DFF_1169.D ;
  assign WX8277 = \DFF_1169.Q ;
  assign WX8278 = \DFF_1170.D ;
  assign WX8279 = \DFF_1170.Q ;
  assign WX828 = \DFF_124.D ;
  assign WX8280 = \DFF_1171.D ;
  assign WX8281 = \DFF_1171.Q ;
  assign WX8282 = \DFF_1172.D ;
  assign WX8283 = \DFF_1172.Q ;
  assign WX8284 = \DFF_1173.D ;
  assign WX8285 = \DFF_1173.Q ;
  assign WX8286 = \DFF_1174.D ;
  assign WX8287 = \DFF_1174.Q ;
  assign WX8288 = \DFF_1175.D ;
  assign WX8289 = \DFF_1175.Q ;
  assign WX829 = \DFF_124.Q ;
  assign WX8290 = \DFF_1176.D ;
  assign WX8291 = \DFF_1176.Q ;
  assign WX8292 = \DFF_1177.D ;
  assign WX8293 = \DFF_1177.Q ;
  assign WX8294 = \DFF_1178.D ;
  assign WX8295 = \DFF_1178.Q ;
  assign WX8296 = \DFF_1179.D ;
  assign WX8297 = \DFF_1179.Q ;
  assign WX8298 = \DFF_1180.D ;
  assign WX8299 = \DFF_1180.Q ;
  assign WX830 = \DFF_125.D ;
  assign WX8300 = \DFF_1181.D ;
  assign WX8301 = \DFF_1181.Q ;
  assign WX8302 = \DFF_1182.D ;
  assign WX8303 = \DFF_1182.Q ;
  assign WX8304 = \DFF_1183.D ;
  assign WX8305 = \DFF_1183.Q ;
  assign WX831 = \DFF_125.Q ;
  assign WX832 = \DFF_126.D ;
  assign WX833 = \DFF_126.Q ;
  assign WX834 = \DFF_127.D ;
  assign WX835 = \DFF_127.Q ;
  assign WX836 = \DFF_128.D ;
  assign WX837 = \DFF_128.Q ;
  assign WX838 = \DFF_129.D ;
  assign WX839 = \DFF_129.Q ;
  assign WX840 = \DFF_130.D ;
  assign WX8402 = \DFF_1184.D ;
  assign WX8403 = \DFF_1184.Q ;
  assign WX8404 = \DFF_1185.D ;
  assign WX8405 = \DFF_1185.Q ;
  assign WX8406 = \DFF_1186.D ;
  assign WX8407 = \DFF_1186.Q ;
  assign WX8408 = \DFF_1187.D ;
  assign WX8409 = \DFF_1187.Q ;
  assign WX841 = \DFF_130.Q ;
  assign WX8410 = \DFF_1188.D ;
  assign WX8411 = \DFF_1188.Q ;
  assign WX8412 = \DFF_1189.D ;
  assign WX8413 = \DFF_1189.Q ;
  assign WX8414 = \DFF_1190.D ;
  assign WX8415 = \DFF_1190.Q ;
  assign WX8416 = \DFF_1191.D ;
  assign WX8417 = \DFF_1191.Q ;
  assign WX8418 = \DFF_1192.D ;
  assign WX8419 = \DFF_1192.Q ;
  assign WX842 = \DFF_131.D ;
  assign WX8420 = \DFF_1193.D ;
  assign WX8421 = \DFF_1193.Q ;
  assign WX8422 = \DFF_1194.D ;
  assign WX8423 = \DFF_1194.Q ;
  assign WX8424 = \DFF_1195.D ;
  assign WX8425 = \DFF_1195.Q ;
  assign WX8426 = \DFF_1196.D ;
  assign WX8427 = \DFF_1196.Q ;
  assign WX8428 = \DFF_1197.D ;
  assign WX8429 = \DFF_1197.Q ;
  assign WX843 = \DFF_131.Q ;
  assign WX8430 = \DFF_1198.D ;
  assign WX8431 = \DFF_1198.Q ;
  assign WX8432 = \DFF_1199.D ;
  assign WX8433 = \DFF_1199.Q ;
  assign WX8434 = \DFF_1200.D ;
  assign WX8435 = \DFF_1200.Q ;
  assign WX8436 = \DFF_1201.D ;
  assign WX8437 = \DFF_1201.Q ;
  assign WX8438 = \DFF_1202.D ;
  assign WX8439 = \DFF_1202.Q ;
  assign WX844 = \DFF_132.D ;
  assign WX8440 = \DFF_1203.D ;
  assign WX8441 = \DFF_1203.Q ;
  assign WX8442 = \DFF_1204.D ;
  assign WX8443 = \DFF_1204.Q ;
  assign WX8444 = \DFF_1205.D ;
  assign WX8445 = \DFF_1205.Q ;
  assign WX8446 = \DFF_1206.D ;
  assign WX8447 = \DFF_1206.Q ;
  assign WX8448 = \DFF_1207.D ;
  assign WX8449 = \DFF_1207.Q ;
  assign WX845 = \DFF_132.Q ;
  assign WX8450 = \DFF_1208.D ;
  assign WX8451 = \DFF_1208.Q ;
  assign WX8452 = \DFF_1209.D ;
  assign WX8453 = \DFF_1209.Q ;
  assign WX8454 = \DFF_1210.D ;
  assign WX8455 = \DFF_1210.Q ;
  assign WX8456 = \DFF_1211.D ;
  assign WX8457 = \DFF_1211.Q ;
  assign WX8458 = \DFF_1212.D ;
  assign WX8459 = \DFF_1212.Q ;
  assign WX846 = \DFF_133.D ;
  assign WX8460 = \DFF_1213.D ;
  assign WX8461 = \DFF_1213.Q ;
  assign WX8462 = \DFF_1214.D ;
  assign WX8463 = \DFF_1214.Q ;
  assign WX8464 = \DFF_1215.D ;
  assign WX8465 = \DFF_1215.Q ;
  assign WX8466 = \DFF_1216.D ;
  assign WX8467 = \DFF_1216.Q ;
  assign WX8468 = \DFF_1217.D ;
  assign WX8469 = \DFF_1217.Q ;
  assign WX847 = \DFF_133.Q ;
  assign WX8470 = \DFF_1218.D ;
  assign WX8471 = \DFF_1218.Q ;
  assign WX8472 = \DFF_1219.D ;
  assign WX8473 = \DFF_1219.Q ;
  assign WX8474 = \DFF_1220.D ;
  assign WX8475 = \DFF_1220.Q ;
  assign WX8476 = \DFF_1221.D ;
  assign WX8477 = \DFF_1221.Q ;
  assign WX8478 = \DFF_1222.D ;
  assign WX8479 = \DFF_1222.Q ;
  assign WX848 = \DFF_134.D ;
  assign WX8480 = \DFF_1223.D ;
  assign WX8481 = \DFF_1223.Q ;
  assign WX8482 = \DFF_1224.D ;
  assign WX8483 = \DFF_1224.Q ;
  assign WX8484 = \DFF_1225.D ;
  assign WX8485 = \DFF_1225.Q ;
  assign WX8486 = \DFF_1226.D ;
  assign WX8487 = \DFF_1226.Q ;
  assign WX8488 = \DFF_1227.D ;
  assign WX8489 = \DFF_1227.Q ;
  assign WX849 = \DFF_134.Q ;
  assign WX8490 = \DFF_1228.D ;
  assign WX8491 = \DFF_1228.Q ;
  assign WX8492 = \DFF_1229.D ;
  assign WX8493 = \DFF_1229.Q ;
  assign WX8494 = \DFF_1230.D ;
  assign WX8495 = \DFF_1230.Q ;
  assign WX8496 = \DFF_1231.D ;
  assign WX8497 = \DFF_1231.Q ;
  assign WX8498 = \DFF_1232.D ;
  assign WX8499 = \DFF_1232.Q ;
  assign WX850 = \DFF_135.D ;
  assign WX8500 = \DFF_1233.D ;
  assign WX8501 = \DFF_1233.Q ;
  assign WX8502 = \DFF_1234.D ;
  assign WX8503 = \DFF_1234.Q ;
  assign WX8504 = \DFF_1235.D ;
  assign WX8505 = \DFF_1235.Q ;
  assign WX8506 = \DFF_1236.D ;
  assign WX8507 = \DFF_1236.Q ;
  assign WX8508 = \DFF_1237.D ;
  assign WX8509 = \DFF_1237.Q ;
  assign WX851 = \DFF_135.Q ;
  assign WX8510 = \DFF_1238.D ;
  assign WX8511 = \DFF_1238.Q ;
  assign WX8512 = \DFF_1239.D ;
  assign WX8513 = \DFF_1239.Q ;
  assign WX8514 = \DFF_1240.D ;
  assign WX8515 = \DFF_1240.Q ;
  assign WX8516 = \DFF_1241.D ;
  assign WX8517 = \DFF_1241.Q ;
  assign WX8518 = \DFF_1242.D ;
  assign WX8519 = \DFF_1242.Q ;
  assign WX852 = \DFF_136.D ;
  assign WX8520 = \DFF_1243.D ;
  assign WX8521 = \DFF_1243.Q ;
  assign WX8522 = \DFF_1244.D ;
  assign WX8523 = \DFF_1244.Q ;
  assign WX8524 = \DFF_1245.D ;
  assign WX8525 = \DFF_1245.Q ;
  assign WX8526 = \DFF_1246.D ;
  assign WX8527 = \DFF_1246.Q ;
  assign WX8528 = \DFF_1247.D ;
  assign WX8529 = \DFF_1247.Q ;
  assign WX853 = \DFF_136.Q ;
  assign WX8530 = \DFF_1248.D ;
  assign WX8531 = \DFF_1248.Q ;
  assign WX8532 = \DFF_1249.D ;
  assign WX8533 = \DFF_1249.Q ;
  assign WX8534 = \DFF_1250.D ;
  assign WX8535 = \DFF_1250.Q ;
  assign WX8536 = \DFF_1251.D ;
  assign WX8537 = \DFF_1251.Q ;
  assign WX8538 = \DFF_1252.D ;
  assign WX8539 = \DFF_1252.Q ;
  assign WX854 = \DFF_137.D ;
  assign WX8540 = \DFF_1253.D ;
  assign WX8541 = \DFF_1253.Q ;
  assign WX8542 = \DFF_1254.D ;
  assign WX8543 = \DFF_1254.Q ;
  assign WX8544 = \DFF_1255.D ;
  assign WX8545 = \DFF_1255.Q ;
  assign WX8546 = \DFF_1256.D ;
  assign WX8547 = \DFF_1256.Q ;
  assign WX8548 = \DFF_1257.D ;
  assign WX8549 = \DFF_1257.Q ;
  assign WX855 = \DFF_137.Q ;
  assign WX8550 = \DFF_1258.D ;
  assign WX8551 = \DFF_1258.Q ;
  assign WX8552 = \DFF_1259.D ;
  assign WX8553 = \DFF_1259.Q ;
  assign WX8554 = \DFF_1260.D ;
  assign WX8555 = \DFF_1260.Q ;
  assign WX8556 = \DFF_1261.D ;
  assign WX8557 = \DFF_1261.Q ;
  assign WX8558 = \DFF_1262.D ;
  assign WX8559 = \DFF_1262.Q ;
  assign WX856 = \DFF_138.D ;
  assign WX8560 = \DFF_1263.D ;
  assign WX8561 = \DFF_1263.Q ;
  assign WX8562 = \DFF_1264.D ;
  assign WX8563 = \DFF_1264.Q ;
  assign WX8564 = \DFF_1265.D ;
  assign WX8565 = \DFF_1265.Q ;
  assign WX8566 = \DFF_1266.D ;
  assign WX8567 = \DFF_1266.Q ;
  assign WX8568 = \DFF_1267.D ;
  assign WX8569 = \DFF_1267.Q ;
  assign WX857 = \DFF_138.Q ;
  assign WX8570 = \DFF_1268.D ;
  assign WX8571 = \DFF_1268.Q ;
  assign WX8572 = \DFF_1269.D ;
  assign WX8573 = \DFF_1269.Q ;
  assign WX8574 = \DFF_1270.D ;
  assign WX8575 = \DFF_1270.Q ;
  assign WX8576 = \DFF_1271.D ;
  assign WX8577 = \DFF_1271.Q ;
  assign WX8578 = \DFF_1272.D ;
  assign WX8579 = \DFF_1272.Q ;
  assign WX858 = \DFF_139.D ;
  assign WX8580 = \DFF_1273.D ;
  assign WX8581 = \DFF_1273.Q ;
  assign WX8582 = \DFF_1274.D ;
  assign WX8583 = \DFF_1274.Q ;
  assign WX8584 = \DFF_1275.D ;
  assign WX8585 = \DFF_1275.Q ;
  assign WX8586 = \DFF_1276.D ;
  assign WX8587 = \DFF_1276.Q ;
  assign WX8588 = \DFF_1277.D ;
  assign WX8589 = \DFF_1277.Q ;
  assign WX859 = \DFF_139.Q ;
  assign WX8590 = \DFF_1278.D ;
  assign WX8591 = \DFF_1278.Q ;
  assign WX8592 = \DFF_1279.D ;
  assign WX8593 = \DFF_1279.Q ;
  assign WX8594 = \DFF_1280.D ;
  assign WX8595 = \DFF_1280.Q ;
  assign WX8596 = \DFF_1281.D ;
  assign WX8597 = \DFF_1281.Q ;
  assign WX8598 = \DFF_1282.D ;
  assign WX8599 = \DFF_1282.Q ;
  assign WX860 = \DFF_140.D ;
  assign WX8600 = \DFF_1283.D ;
  assign WX8601 = \DFF_1283.Q ;
  assign WX8602 = \DFF_1284.D ;
  assign WX8603 = \DFF_1284.Q ;
  assign WX8604 = \DFF_1285.D ;
  assign WX8605 = \DFF_1285.Q ;
  assign WX8606 = \DFF_1286.D ;
  assign WX8607 = \DFF_1286.Q ;
  assign WX8608 = \DFF_1287.D ;
  assign WX8609 = \DFF_1287.Q ;
  assign WX861 = \DFF_140.Q ;
  assign WX8610 = \DFF_1288.D ;
  assign WX8611 = \DFF_1288.Q ;
  assign WX8612 = \DFF_1289.D ;
  assign WX8613 = \DFF_1289.Q ;
  assign WX8614 = \DFF_1290.D ;
  assign WX8615 = \DFF_1290.Q ;
  assign WX8616 = \DFF_1291.D ;
  assign WX8617 = \DFF_1291.Q ;
  assign WX8618 = \DFF_1292.D ;
  assign WX8619 = \DFF_1292.Q ;
  assign WX862 = \DFF_141.D ;
  assign WX8620 = \DFF_1293.D ;
  assign WX8621 = \DFF_1293.Q ;
  assign WX8622 = \DFF_1294.D ;
  assign WX8623 = \DFF_1294.Q ;
  assign WX8624 = \DFF_1295.D ;
  assign WX8625 = \DFF_1295.Q ;
  assign WX8626 = \DFF_1296.D ;
  assign WX8627 = \DFF_1296.Q ;
  assign WX8628 = \DFF_1297.D ;
  assign WX8629 = \DFF_1297.Q ;
  assign WX863 = \DFF_141.Q ;
  assign WX8630 = \DFF_1298.D ;
  assign WX8631 = \DFF_1298.Q ;
  assign WX8632 = \DFF_1299.D ;
  assign WX8633 = \DFF_1299.Q ;
  assign WX8634 = \DFF_1300.D ;
  assign WX8635 = \DFF_1300.Q ;
  assign WX8636 = \DFF_1301.D ;
  assign WX8637 = \DFF_1301.Q ;
  assign WX8638 = \DFF_1302.D ;
  assign WX8639 = \DFF_1302.Q ;
  assign WX864 = \DFF_142.D ;
  assign WX8640 = \DFF_1303.D ;
  assign WX8641 = \DFF_1303.Q ;
  assign WX8642 = \DFF_1304.D ;
  assign WX8643 = \DFF_1304.Q ;
  assign WX8644 = \DFF_1305.D ;
  assign WX8645 = \DFF_1305.Q ;
  assign WX8646 = \DFF_1306.D ;
  assign WX8647 = \DFF_1306.Q ;
  assign WX8648 = \DFF_1307.D ;
  assign WX8649 = \DFF_1307.Q ;
  assign WX865 = \DFF_142.Q ;
  assign WX8650 = \DFF_1308.D ;
  assign WX8651 = \DFF_1308.Q ;
  assign WX8652 = \DFF_1309.D ;
  assign WX8653 = \DFF_1309.Q ;
  assign WX8654 = \DFF_1310.D ;
  assign WX8655 = \DFF_1310.Q ;
  assign WX8656 = \DFF_1311.D ;
  assign WX8657 = \DFF_1311.Q ;
  assign WX866 = \DFF_143.D ;
  assign WX867 = \DFF_143.Q ;
  assign WX868 = \DFF_144.D ;
  assign WX869 = \DFF_144.Q ;
  assign WX870 = \DFF_145.D ;
  assign WX871 = \DFF_145.Q ;
  assign WX872 = \DFF_146.D ;
  assign WX873 = \DFF_146.Q ;
  assign WX874 = \DFF_147.D ;
  assign WX875 = \DFF_147.Q ;
  assign WX8759 = TM1;
  assign WX876 = \DFF_148.D ;
  assign WX8760 = TM0;
  assign WX8761 = TM1;
  assign WX8762 = TM0;
  assign WX8763 = TM0;
  assign WX877 = \DFF_148.Q ;
  assign WX878 = \DFF_149.D ;
  assign WX879 = \DFF_149.Q ;
  assign WX880 = \DFF_150.D ;
  assign WX881 = \DFF_150.Q ;
  assign WX882 = \DFF_151.D ;
  assign WX883 = \DFF_151.Q ;
  assign WX884 = \DFF_152.D ;
  assign WX885 = \DFF_152.Q ;
  assign WX886 = \DFF_153.D ;
  assign WX887 = \DFF_153.Q ;
  assign WX888 = \DFF_154.D ;
  assign WX889 = \DFF_154.Q ;
  assign WX890 = \DFF_155.D ;
  assign WX891 = \DFF_155.Q ;
  assign WX892 = \DFF_156.D ;
  assign WX893 = \DFF_156.Q ;
  assign WX894 = \DFF_157.D ;
  assign WX895 = \DFF_157.Q ;
  assign WX896 = \DFF_158.D ;
  assign WX897 = \DFF_158.Q ;
  assign WX898 = \DFF_159.D ;
  assign WX899 = \DFF_159.Q ;
  assign WX9021 = RESET;
  assign WX9022 = \DFF_1312.D ;
  assign WX9024 = \DFF_1313.D ;
  assign WX9026 = \DFF_1314.D ;
  assign WX9028 = \DFF_1315.D ;
  assign WX9030 = \DFF_1316.D ;
  assign WX9032 = \DFF_1317.D ;
  assign WX9034 = \DFF_1318.D ;
  assign WX9036 = \DFF_1319.D ;
  assign WX9038 = \DFF_1320.D ;
  assign WX9040 = \DFF_1321.D ;
  assign WX9042 = \DFF_1322.D ;
  assign WX9044 = \DFF_1323.D ;
  assign WX9046 = \DFF_1324.D ;
  assign WX9048 = \DFF_1325.D ;
  assign WX9050 = \DFF_1326.D ;
  assign WX9052 = \DFF_1327.D ;
  assign WX9054 = \DFF_1328.D ;
  assign WX9056 = \DFF_1329.D ;
  assign WX9058 = \DFF_1330.D ;
  assign WX9060 = \DFF_1331.D ;
  assign WX9062 = \DFF_1332.D ;
  assign WX9064 = \DFF_1333.D ;
  assign WX9066 = \DFF_1334.D ;
  assign WX9068 = \DFF_1335.D ;
  assign WX9070 = \DFF_1336.D ;
  assign WX9072 = \DFF_1337.D ;
  assign WX9074 = \DFF_1338.D ;
  assign WX9076 = \DFF_1339.D ;
  assign WX9078 = \DFF_1340.D ;
  assign WX9080 = \DFF_1341.D ;
  assign WX9082 = \DFF_1342.D ;
  assign WX9084 = \DFF_1343.D ;
  assign WX9535 = \DFF_1344.D ;
  assign WX9536 = \DFF_1344.Q ;
  assign WX9537 = \DFF_1345.D ;
  assign WX9538 = \DFF_1345.Q ;
  assign WX9539 = \DFF_1346.D ;
  assign WX9540 = \DFF_1346.Q ;
  assign WX9541 = \DFF_1347.D ;
  assign WX9542 = \DFF_1347.Q ;
  assign WX9543 = \DFF_1348.D ;
  assign WX9544 = \DFF_1348.Q ;
  assign WX9545 = \DFF_1349.D ;
  assign WX9546 = \DFF_1349.Q ;
  assign WX9547 = \DFF_1350.D ;
  assign WX9548 = \DFF_1350.Q ;
  assign WX9549 = \DFF_1351.D ;
  assign WX9550 = \DFF_1351.Q ;
  assign WX9551 = \DFF_1352.D ;
  assign WX9552 = \DFF_1352.Q ;
  assign WX9553 = \DFF_1353.D ;
  assign WX9554 = \DFF_1353.Q ;
  assign WX9555 = \DFF_1354.D ;
  assign WX9556 = \DFF_1354.Q ;
  assign WX9557 = \DFF_1355.D ;
  assign WX9558 = \DFF_1355.Q ;
  assign WX9559 = \DFF_1356.D ;
  assign WX9560 = \DFF_1356.Q ;
  assign WX9561 = \DFF_1357.D ;
  assign WX9562 = \DFF_1357.Q ;
  assign WX9563 = \DFF_1358.D ;
  assign WX9564 = \DFF_1358.Q ;
  assign WX9565 = \DFF_1359.D ;
  assign WX9566 = \DFF_1359.Q ;
  assign WX9567 = \DFF_1360.D ;
  assign WX9568 = \DFF_1360.Q ;
  assign WX9569 = \DFF_1361.D ;
  assign WX9570 = \DFF_1361.Q ;
  assign WX9571 = \DFF_1362.D ;
  assign WX9572 = \DFF_1362.Q ;
  assign WX9573 = \DFF_1363.D ;
  assign WX9574 = \DFF_1363.Q ;
  assign WX9575 = \DFF_1364.D ;
  assign WX9576 = \DFF_1364.Q ;
  assign WX9577 = \DFF_1365.D ;
  assign WX9578 = \DFF_1365.Q ;
  assign WX9579 = \DFF_1366.D ;
  assign WX9580 = \DFF_1366.Q ;
  assign WX9581 = \DFF_1367.D ;
  assign WX9582 = \DFF_1367.Q ;
  assign WX9583 = \DFF_1368.D ;
  assign WX9584 = \DFF_1368.Q ;
  assign WX9585 = \DFF_1369.D ;
  assign WX9586 = \DFF_1369.Q ;
  assign WX9587 = \DFF_1370.D ;
  assign WX9588 = \DFF_1370.Q ;
  assign WX9589 = \DFF_1371.D ;
  assign WX9590 = \DFF_1371.Q ;
  assign WX9591 = \DFF_1372.D ;
  assign WX9592 = \DFF_1372.Q ;
  assign WX9593 = \DFF_1373.D ;
  assign WX9594 = \DFF_1373.Q ;
  assign WX9595 = \DFF_1374.D ;
  assign WX9596 = \DFF_1374.Q ;
  assign WX9597 = \DFF_1375.D ;
  assign WX9598 = \DFF_1375.Q ;
  assign WX9695 = \DFF_1376.D ;
  assign WX9696 = \DFF_1376.Q ;
  assign WX9697 = \DFF_1377.D ;
  assign WX9698 = \DFF_1377.Q ;
  assign WX9699 = \DFF_1378.D ;
  assign WX9700 = \DFF_1378.Q ;
  assign WX9701 = \DFF_1379.D ;
  assign WX9702 = \DFF_1379.Q ;
  assign WX9703 = \DFF_1380.D ;
  assign WX9704 = \DFF_1380.Q ;
  assign WX9705 = \DFF_1381.D ;
  assign WX9706 = \DFF_1381.Q ;
  assign WX9707 = \DFF_1382.D ;
  assign WX9708 = \DFF_1382.Q ;
  assign WX9709 = \DFF_1383.D ;
  assign WX9710 = \DFF_1383.Q ;
  assign WX9711 = \DFF_1384.D ;
  assign WX9712 = \DFF_1384.Q ;
  assign WX9713 = \DFF_1385.D ;
  assign WX9714 = \DFF_1385.Q ;
  assign WX9715 = \DFF_1386.D ;
  assign WX9716 = \DFF_1386.Q ;
  assign WX9717 = \DFF_1387.D ;
  assign WX9718 = \DFF_1387.Q ;
  assign WX9719 = \DFF_1388.D ;
  assign WX9720 = \DFF_1388.Q ;
  assign WX9721 = \DFF_1389.D ;
  assign WX9722 = \DFF_1389.Q ;
  assign WX9723 = \DFF_1390.D ;
  assign WX9724 = \DFF_1390.Q ;
  assign WX9725 = \DFF_1391.D ;
  assign WX9726 = \DFF_1391.Q ;
  assign WX9727 = \DFF_1392.D ;
  assign WX9728 = \DFF_1392.Q ;
  assign WX9729 = \DFF_1393.D ;
  assign WX9730 = \DFF_1393.Q ;
  assign WX9731 = \DFF_1394.D ;
  assign WX9732 = \DFF_1394.Q ;
  assign WX9733 = \DFF_1395.D ;
  assign WX9734 = \DFF_1395.Q ;
  assign WX9735 = \DFF_1396.D ;
  assign WX9736 = \DFF_1396.Q ;
  assign WX9737 = \DFF_1397.D ;
  assign WX9738 = \DFF_1397.Q ;
  assign WX9739 = \DFF_1398.D ;
  assign WX9740 = \DFF_1398.Q ;
  assign WX9741 = \DFF_1399.D ;
  assign WX9742 = \DFF_1399.Q ;
  assign WX9743 = \DFF_1400.D ;
  assign WX9744 = \DFF_1400.Q ;
  assign WX9745 = \DFF_1401.D ;
  assign WX9746 = \DFF_1401.Q ;
  assign WX9747 = \DFF_1402.D ;
  assign WX9748 = \DFF_1402.Q ;
  assign WX9749 = \DFF_1403.D ;
  assign WX9750 = \DFF_1403.Q ;
  assign WX9751 = \DFF_1404.D ;
  assign WX9752 = \DFF_1404.Q ;
  assign WX9753 = \DFF_1405.D ;
  assign WX9754 = \DFF_1405.Q ;
  assign WX9755 = \DFF_1406.D ;
  assign WX9756 = \DFF_1406.Q ;
  assign WX9757 = \DFF_1407.D ;
  assign WX9758 = \DFF_1407.Q ;
  assign WX9759 = \DFF_1408.D ;
  assign WX9760 = \DFF_1408.Q ;
  assign WX9761 = \DFF_1409.D ;
  assign WX9762 = \DFF_1409.Q ;
  assign WX9763 = \DFF_1410.D ;
  assign WX9764 = \DFF_1410.Q ;
  assign WX9765 = \DFF_1411.D ;
  assign WX9766 = \DFF_1411.Q ;
  assign WX9767 = \DFF_1412.D ;
  assign WX9768 = \DFF_1412.Q ;
  assign WX9769 = \DFF_1413.D ;
  assign WX9770 = \DFF_1413.Q ;
  assign WX9771 = \DFF_1414.D ;
  assign WX9772 = \DFF_1414.Q ;
  assign WX9773 = \DFF_1415.D ;
  assign WX9774 = \DFF_1415.Q ;
  assign WX9775 = \DFF_1416.D ;
  assign WX9776 = \DFF_1416.Q ;
  assign WX9777 = \DFF_1417.D ;
  assign WX9778 = \DFF_1417.Q ;
  assign WX9779 = \DFF_1418.D ;
  assign WX9780 = \DFF_1418.Q ;
  assign WX9781 = \DFF_1419.D ;
  assign WX9782 = \DFF_1419.Q ;
  assign WX9783 = \DFF_1420.D ;
  assign WX9784 = \DFF_1420.Q ;
  assign WX9785 = \DFF_1421.D ;
  assign WX9786 = \DFF_1421.Q ;
  assign WX9787 = \DFF_1422.D ;
  assign WX9788 = \DFF_1422.Q ;
  assign WX9789 = \DFF_1423.D ;
  assign WX9790 = \DFF_1423.Q ;
  assign WX9791 = \DFF_1424.D ;
  assign WX9792 = \DFF_1424.Q ;
  assign WX9793 = \DFF_1425.D ;
  assign WX9794 = \DFF_1425.Q ;
  assign WX9795 = \DFF_1426.D ;
  assign WX9796 = \DFF_1426.Q ;
  assign WX9797 = \DFF_1427.D ;
  assign WX9798 = \DFF_1427.Q ;
  assign WX9799 = \DFF_1428.D ;
  assign WX9800 = \DFF_1428.Q ;
  assign WX9801 = \DFF_1429.D ;
  assign WX9802 = \DFF_1429.Q ;
  assign WX9803 = \DFF_1430.D ;
  assign WX9804 = \DFF_1430.Q ;
  assign WX9805 = \DFF_1431.D ;
  assign WX9806 = \DFF_1431.Q ;
  assign WX9807 = \DFF_1432.D ;
  assign WX9808 = \DFF_1432.Q ;
  assign WX9809 = \DFF_1433.D ;
  assign WX9810 = \DFF_1433.Q ;
  assign WX9811 = \DFF_1434.D ;
  assign WX9812 = \DFF_1434.Q ;
  assign WX9813 = \DFF_1435.D ;
  assign WX9814 = \DFF_1435.Q ;
  assign WX9815 = \DFF_1436.D ;
  assign WX9816 = \DFF_1436.Q ;
  assign WX9817 = \DFF_1437.D ;
  assign WX9818 = \DFF_1437.Q ;
  assign WX9819 = \DFF_1438.D ;
  assign WX9820 = \DFF_1438.Q ;
  assign WX9821 = \DFF_1439.D ;
  assign WX9822 = \DFF_1439.Q ;
  assign WX9823 = \DFF_1440.D ;
  assign WX9824 = \DFF_1440.Q ;
  assign WX9825 = \DFF_1441.D ;
  assign WX9826 = \DFF_1441.Q ;
  assign WX9827 = \DFF_1442.D ;
  assign WX9828 = \DFF_1442.Q ;
  assign WX9829 = \DFF_1443.D ;
  assign WX9830 = \DFF_1443.Q ;
  assign WX9831 = \DFF_1444.D ;
  assign WX9832 = \DFF_1444.Q ;
  assign WX9833 = \DFF_1445.D ;
  assign WX9834 = \DFF_1445.Q ;
  assign WX9835 = \DFF_1446.D ;
  assign WX9836 = \DFF_1446.Q ;
  assign WX9837 = \DFF_1447.D ;
  assign WX9838 = \DFF_1447.Q ;
  assign WX9839 = \DFF_1448.D ;
  assign WX9840 = \DFF_1448.Q ;
  assign WX9841 = \DFF_1449.D ;
  assign WX9842 = \DFF_1449.Q ;
  assign WX9843 = \DFF_1450.D ;
  assign WX9844 = \DFF_1450.Q ;
  assign WX9845 = \DFF_1451.D ;
  assign WX9846 = \DFF_1451.Q ;
  assign WX9847 = \DFF_1452.D ;
  assign WX9848 = \DFF_1452.Q ;
  assign WX9849 = \DFF_1453.D ;
  assign WX9850 = \DFF_1453.Q ;
  assign WX9851 = \DFF_1454.D ;
  assign WX9852 = \DFF_1454.Q ;
  assign WX9853 = \DFF_1455.D ;
  assign WX9854 = \DFF_1455.Q ;
  assign WX9855 = \DFF_1456.D ;
  assign WX9856 = \DFF_1456.Q ;
  assign WX9857 = \DFF_1457.D ;
  assign WX9858 = \DFF_1457.Q ;
  assign WX9859 = \DFF_1458.D ;
  assign WX9860 = \DFF_1458.Q ;
  assign WX9861 = \DFF_1459.D ;
  assign WX9862 = \DFF_1459.Q ;
  assign WX9863 = \DFF_1460.D ;
  assign WX9864 = \DFF_1460.Q ;
  assign WX9865 = \DFF_1461.D ;
  assign WX9866 = \DFF_1461.Q ;
  assign WX9867 = \DFF_1462.D ;
  assign WX9868 = \DFF_1462.Q ;
  assign WX9869 = \DFF_1463.D ;
  assign WX9870 = \DFF_1463.Q ;
  assign WX9871 = \DFF_1464.D ;
  assign WX9872 = \DFF_1464.Q ;
  assign WX9873 = \DFF_1465.D ;
  assign WX9874 = \DFF_1465.Q ;
  assign WX9875 = \DFF_1466.D ;
  assign WX9876 = \DFF_1466.Q ;
  assign WX9877 = \DFF_1467.D ;
  assign WX9878 = \DFF_1467.Q ;
  assign WX9879 = \DFF_1468.D ;
  assign WX9880 = \DFF_1468.Q ;
  assign WX9881 = \DFF_1469.D ;
  assign WX9882 = \DFF_1469.Q ;
  assign WX9883 = \DFF_1470.D ;
  assign WX9884 = \DFF_1470.Q ;
  assign WX9885 = \DFF_1471.D ;
  assign WX9886 = \DFF_1471.Q ;
  assign WX9887 = \DFF_1472.D ;
  assign WX9888 = \DFF_1472.Q ;
  assign WX9889 = \DFF_1473.D ;
  assign WX9890 = \DFF_1473.Q ;
  assign WX9891 = \DFF_1474.D ;
  assign WX9892 = \DFF_1474.Q ;
  assign WX9893 = \DFF_1475.D ;
  assign WX9894 = \DFF_1475.Q ;
  assign WX9895 = \DFF_1476.D ;
  assign WX9896 = \DFF_1476.Q ;
  assign WX9897 = \DFF_1477.D ;
  assign WX9898 = \DFF_1477.Q ;
  assign WX9899 = \DFF_1478.D ;
  assign WX9900 = \DFF_1478.Q ;
  assign WX9901 = \DFF_1479.D ;
  assign WX9902 = \DFF_1479.Q ;
  assign WX9903 = \DFF_1480.D ;
  assign WX9904 = \DFF_1480.Q ;
  assign WX9905 = \DFF_1481.D ;
  assign WX9906 = \DFF_1481.Q ;
  assign WX9907 = \DFF_1482.D ;
  assign WX9908 = \DFF_1482.Q ;
  assign WX9909 = \DFF_1483.D ;
  assign WX9910 = \DFF_1483.Q ;
  assign WX9911 = \DFF_1484.D ;
  assign WX9912 = \DFF_1484.Q ;
  assign WX9913 = \DFF_1485.D ;
  assign WX9914 = \DFF_1485.Q ;
  assign WX9915 = \DFF_1486.D ;
  assign WX9916 = \DFF_1486.Q ;
  assign WX9917 = \DFF_1487.D ;
  assign WX9918 = \DFF_1487.Q ;
  assign WX9919 = \DFF_1488.D ;
  assign WX9920 = \DFF_1488.Q ;
  assign WX9921 = \DFF_1489.D ;
  assign WX9922 = \DFF_1489.Q ;
  assign WX9923 = \DFF_1490.D ;
  assign WX9924 = \DFF_1490.Q ;
  assign WX9925 = \DFF_1491.D ;
  assign WX9926 = \DFF_1491.Q ;
  assign WX9927 = \DFF_1492.D ;
  assign WX9928 = \DFF_1492.Q ;
  assign WX9929 = \DFF_1493.D ;
  assign WX9930 = \DFF_1493.Q ;
  assign WX9931 = \DFF_1494.D ;
  assign WX9932 = \DFF_1494.Q ;
  assign WX9933 = \DFF_1495.D ;
  assign WX9934 = \DFF_1495.Q ;
  assign WX9935 = \DFF_1496.D ;
  assign WX9936 = \DFF_1496.Q ;
  assign WX9937 = \DFF_1497.D ;
  assign WX9938 = \DFF_1497.Q ;
  assign WX9939 = \DFF_1498.D ;
  assign WX9940 = \DFF_1498.Q ;
  assign WX9941 = \DFF_1499.D ;
  assign WX9942 = \DFF_1499.Q ;
  assign WX9943 = \DFF_1500.D ;
  assign WX9944 = \DFF_1500.Q ;
  assign WX9945 = \DFF_1501.D ;
  assign WX9946 = \DFF_1501.Q ;
  assign WX9947 = \DFF_1502.D ;
  assign WX9948 = \DFF_1502.Q ;
  assign WX9949 = \DFF_1503.D ;
  assign WX9950 = \DFF_1503.Q ;
endmodule
