
module s1238(GND, VDD, CK, G0, G1, G10, G11, G12, G13, G2, G3, G4, G45, G5, G530, G532, G535, G537, G539, G542, G546, G547, G548, G549, G550, G551, G552, G6, G7, G8, G9);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  input CK;
  wire \DFF_0.CK ;
  wire \DFF_0.D ;
  wire \DFF_0.Q ;
  wire \DFF_1.CK ;
  wire \DFF_1.D ;
  wire \DFF_1.Q ;
  wire \DFF_10.CK ;
  wire \DFF_10.D ;
  wire \DFF_10.Q ;
  wire \DFF_11.CK ;
  wire \DFF_11.D ;
  wire \DFF_11.Q ;
  wire \DFF_12.CK ;
  wire \DFF_12.D ;
  wire \DFF_12.Q ;
  wire \DFF_13.CK ;
  wire \DFF_13.D ;
  wire \DFF_13.Q ;
  wire \DFF_14.CK ;
  wire \DFF_14.D ;
  wire \DFF_14.Q ;
  wire \DFF_15.CK ;
  wire \DFF_15.D ;
  wire \DFF_15.Q ;
  wire \DFF_16.CK ;
  wire \DFF_16.D ;
  wire \DFF_16.Q ;
  wire \DFF_17.CK ;
  wire \DFF_17.D ;
  wire \DFF_17.Q ;
  wire \DFF_2.CK ;
  wire \DFF_2.D ;
  wire \DFF_2.Q ;
  wire \DFF_3.CK ;
  wire \DFF_3.D ;
  wire \DFF_3.Q ;
  wire \DFF_4.CK ;
  wire \DFF_4.D ;
  wire \DFF_4.Q ;
  wire \DFF_5.CK ;
  wire \DFF_5.D ;
  wire \DFF_5.Q ;
  wire \DFF_6.CK ;
  wire \DFF_6.D ;
  wire \DFF_6.Q ;
  wire \DFF_7.CK ;
  wire \DFF_7.D ;
  wire \DFF_7.Q ;
  wire \DFF_8.CK ;
  wire \DFF_8.D ;
  wire \DFF_8.Q ;
  wire \DFF_9.CK ;
  wire \DFF_9.D ;
  wire \DFF_9.Q ;
  input G0;
  input G1;
  input G10;
  input G11;
  input G12;
  input G13;
  input G2;
  wire G29;
  input G3;
  wire G30;
  wire G31;
  wire G32;
  wire G33;
  wire G34;
  wire G35;
  wire G36;
  wire G37;
  wire G38;
  wire G39;
  input G4;
  wire G40;
  wire G41;
  wire G42;
  wire G43;
  wire G44;
  output G45;
  wire G46;
  input G5;
  wire G502;
  wire G503;
  wire G504;
  wire G505;
  wire G506;
  wire G507;
  wire G508;
  wire G509;
  wire G510;
  wire G511;
  wire G512;
  wire G513;
  wire G514;
  wire G515;
  wire G516;
  wire G517;
  wire G518;
  wire G519;
  output G530;
  output G532;
  output G535;
  output G537;
  output G539;
  output G542;
  output G546;
  output G547;
  output G548;
  output G549;
  output G550;
  output G551;
  output G552;
  input G6;
  input G7;
  input G8;
  input G9;
  input GND;
  input VDD;
  al_oai21ftf _296_ (
    .a(G11),
    .b(G9),
    .c(G10),
    .y(\DFF_1.D )
  );
  al_ao21ttf _297_ (
    .a(G9),
    .b(G11),
    .c(G10),
    .y(_265_)
  );
  al_ao21ftf _298_ (
    .a(G7),
    .b(G11),
    .c(_265_),
    .y(\DFF_2.D )
  );
  al_oai21ftf _299_ (
    .a(G6),
    .b(G4),
    .c(G5),
    .y(_266_)
  );
  al_nand3ftt _300_ (
    .a(G2),
    .b(G3),
    .c(_266_),
    .y(_267_)
  );
  al_and3 _301_ (
    .a(G3),
    .b(G4),
    .c(G6),
    .y(_268_)
  );
  al_nand2 _302_ (
    .a(G5),
    .b(_268_),
    .y(_269_)
  );
  al_oai21 _303_ (
    .a(G4),
    .b(G5),
    .c(G2),
    .y(_270_)
  );
  al_ao21ftf _304_ (
    .a(_270_),
    .b(_269_),
    .c(_267_),
    .y(\DFF_3.D )
  );
  al_and3fft _305_ (
    .a(G9),
    .b(G10),
    .c(G7),
    .y(_271_)
  );
  al_and2ft _306_ (
    .a(G8),
    .b(_271_),
    .y(_272_)
  );
  al_nor2 _307_ (
    .a(G7),
    .b(G8),
    .y(_273_)
  );
  al_nand2 _308_ (
    .a(G9),
    .b(G10),
    .y(_274_)
  );
  al_nand2 _309_ (
    .a(G8),
    .b(_271_),
    .y(_275_)
  );
  al_ao21ftf _310_ (
    .a(_274_),
    .b(_273_),
    .c(_275_),
    .y(_276_)
  );
  al_mux2h _311_ (
    .a(_272_),
    .b(_276_),
    .s(G6),
    .y(\DFF_6.D )
  );
  al_and2ft _312_ (
    .a(G6),
    .b(G9),
    .y(_277_)
  );
  al_nand2ft _313_ (
    .a(G9),
    .b(G6),
    .y(_278_)
  );
  al_nand2ft _314_ (
    .a(_277_),
    .b(_278_),
    .y(\DFF_8.D )
  );
  al_nand2ft _315_ (
    .a(G5),
    .b(G2),
    .y(_279_)
  );
  al_nand3ftt _316_ (
    .a(G2),
    .b(G3),
    .c(G5),
    .y(_280_)
  );
  al_nand2ft _317_ (
    .a(G3),
    .b(G2),
    .y(_281_)
  );
  al_nand3 _318_ (
    .a(_280_),
    .b(_279_),
    .c(_281_),
    .y(\DFF_10.D )
  );
  al_inv _319_ (
    .a(G12),
    .y(_282_)
  );
  al_and2 _320_ (
    .a(G1),
    .b(G2),
    .y(_283_)
  );
  al_inv _321_ (
    .a(G0),
    .y(_284_)
  );
  al_and3 _322_ (
    .a(G8),
    .b(G9),
    .c(G11),
    .y(_285_)
  );
  al_and3 _323_ (
    .a(G7),
    .b(G10),
    .c(_285_),
    .y(_286_)
  );
  al_nand3fft _324_ (
    .a(_284_),
    .b(_269_),
    .c(_286_),
    .y(_287_)
  );
  al_nand3fft _325_ (
    .a(G3),
    .b(G8),
    .c(G10),
    .y(_288_)
  );
  al_nor2 _326_ (
    .a(G5),
    .b(G7),
    .y(_289_)
  );
  al_nand3fft _327_ (
    .a(_288_),
    .b(_278_),
    .c(_289_),
    .y(_290_)
  );
  al_and2ft _328_ (
    .a(G10),
    .b(G7),
    .y(_291_)
  );
  al_and3 _329_ (
    .a(G3),
    .b(G5),
    .c(G8),
    .y(_292_)
  );
  al_nand3 _330_ (
    .a(\DFF_8.Q ),
    .b(_291_),
    .c(_292_),
    .y(_293_)
  );
  al_nand3fft _331_ (
    .a(G0),
    .b(G4),
    .c(G11),
    .y(_294_)
  );
  al_ao21 _332_ (
    .a(_293_),
    .b(_290_),
    .c(_294_),
    .y(_295_)
  );
  al_aoi21ttf _333_ (
    .a(_287_),
    .b(_295_),
    .c(_283_),
    .y(_000_)
  );
  al_inv _334_ (
    .a(G11),
    .y(_001_)
  );
  al_or2 _335_ (
    .a(\DFF_1.Q ),
    .b(G6),
    .y(_002_)
  );
  al_aoi21ttf _336_ (
    .a(G8),
    .b(G10),
    .c(G9),
    .y(_003_)
  );
  al_and3ftt _337_ (
    .a(G6),
    .b(\DFF_1.Q ),
    .c(G7),
    .y(_004_)
  );
  al_and3fft _338_ (
    .a(\DFF_2.Q ),
    .b(_004_),
    .c(G8),
    .y(_005_)
  );
  al_oai21ttf _339_ (
    .a(_273_),
    .b(_005_),
    .c(_003_),
    .y(_006_)
  );
  al_ao21 _340_ (
    .a(_002_),
    .b(_006_),
    .c(_001_),
    .y(_007_)
  );
  al_oai21ftf _341_ (
    .a(G5),
    .b(G1),
    .c(G4),
    .y(_008_)
  );
  al_ao21 _342_ (
    .a(G2),
    .b(_008_),
    .c(G3),
    .y(_009_)
  );
  al_oai21ftf _343_ (
    .a(G5),
    .b(G3),
    .c(G4),
    .y(_010_)
  );
  al_ao21 _344_ (
    .a(G0),
    .b(_009_),
    .c(_010_),
    .y(_011_)
  );
  al_or3 _345_ (
    .a(G9),
    .b(G10),
    .c(G11),
    .y(_012_)
  );
  al_nand2 _346_ (
    .a(G8),
    .b(\DFF_2.Q ),
    .y(_013_)
  );
  al_nand3fft _347_ (
    .a(_012_),
    .b(_004_),
    .c(_013_),
    .y(_014_)
  );
  al_inv _348_ (
    .a(G7),
    .y(_015_)
  );
  al_and2ft _349_ (
    .a(G8),
    .b(G10),
    .y(_016_)
  );
  al_ao21ftt _350_ (
    .a(\DFF_2.Q ),
    .b(G8),
    .c(_016_),
    .y(_017_)
  );
  al_and2ft _351_ (
    .a(G11),
    .b(G9),
    .y(_018_)
  );
  al_nand3 _352_ (
    .a(_015_),
    .b(_018_),
    .c(_017_),
    .y(_019_)
  );
  al_and3 _353_ (
    .a(\DFF_17.Q ),
    .b(_014_),
    .c(_019_),
    .y(_020_)
  );
  al_nand3 _354_ (
    .a(_011_),
    .b(_020_),
    .c(_007_),
    .y(_021_)
  );
  al_and2ft _355_ (
    .a(G13),
    .b(G12),
    .y(_022_)
  );
  al_and3 _356_ (
    .a(_022_),
    .b(_000_),
    .c(_021_),
    .y(_023_)
  );
  al_and2ft _357_ (
    .a(G10),
    .b(G9),
    .y(_024_)
  );
  al_nand2ft _358_ (
    .a(G7),
    .b(G8),
    .y(_025_)
  );
  al_aoi21ftf _359_ (
    .a(_025_),
    .b(_024_),
    .c(_275_),
    .y(_026_)
  );
  al_ao21ftf _360_ (
    .a(_274_),
    .b(_273_),
    .c(_026_),
    .y(_027_)
  );
  al_nand2 _361_ (
    .a(G2),
    .b(G5),
    .y(_028_)
  );
  al_nor2 _362_ (
    .a(G10),
    .b(G11),
    .y(_029_)
  );
  al_nand3 _363_ (
    .a(G9),
    .b(_029_),
    .c(_273_),
    .y(_030_)
  );
  al_and3fft _364_ (
    .a(_028_),
    .b(_030_),
    .c(_268_),
    .y(_031_)
  );
  al_and2ft _365_ (
    .a(G5),
    .b(G11),
    .y(_032_)
  );
  al_and3ftt _366_ (
    .a(G2),
    .b(_032_),
    .c(_268_),
    .y(_033_)
  );
  al_aoi21 _367_ (
    .a(_033_),
    .b(_027_),
    .c(_031_),
    .y(_034_)
  );
  al_nor2 _368_ (
    .a(G2),
    .b(G3),
    .y(_035_)
  );
  al_and2ft _369_ (
    .a(G6),
    .b(\DFF_7.Q ),
    .y(_036_)
  );
  al_and2 _370_ (
    .a(G4),
    .b(G6),
    .y(_037_)
  );
  al_and3 _371_ (
    .a(G5),
    .b(G11),
    .c(_037_),
    .y(_038_)
  );
  al_ao21 _372_ (
    .a(_038_),
    .b(_276_),
    .c(_036_),
    .y(_039_)
  );
  al_inv _373_ (
    .a(G2),
    .y(_040_)
  );
  al_and2 _374_ (
    .a(G5),
    .b(_268_),
    .y(_041_)
  );
  al_and2 _375_ (
    .a(G7),
    .b(G10),
    .y(_042_)
  );
  al_nand3 _376_ (
    .a(_285_),
    .b(_042_),
    .c(_041_),
    .y(_043_)
  );
  al_and2ft _377_ (
    .a(G4),
    .b(G3),
    .y(_044_)
  );
  al_nand3 _378_ (
    .a(\DFF_6.Q ),
    .b(_044_),
    .c(_032_),
    .y(_045_)
  );
  al_ao21 _379_ (
    .a(_045_),
    .b(_043_),
    .c(_040_),
    .y(_046_)
  );
  al_aoi21ttf _380_ (
    .a(_035_),
    .b(_039_),
    .c(_046_),
    .y(_047_)
  );
  al_or3fft _381_ (
    .a(G7),
    .b(G10),
    .c(_285_),
    .y(_048_)
  );
  al_nand3ftt _382_ (
    .a(G10),
    .b(G7),
    .c(G9),
    .y(_049_)
  );
  al_nand3ftt _383_ (
    .a(G7),
    .b(\DFF_1.Q ),
    .c(G8),
    .y(_050_)
  );
  al_nand3 _384_ (
    .a(_049_),
    .b(_050_),
    .c(_048_),
    .y(_051_)
  );
  al_ao21 _385_ (
    .a(\DFF_3.Q ),
    .b(_051_),
    .c(G13),
    .y(_052_)
  );
  al_ao21 _386_ (
    .a(_034_),
    .b(_047_),
    .c(_052_),
    .y(_053_)
  );
  al_inv _387_ (
    .a(G13),
    .y(_054_)
  );
  al_and2ft _388_ (
    .a(G2),
    .b(G3),
    .y(_055_)
  );
  al_ao21ttf _389_ (
    .a(G3),
    .b(G5),
    .c(G4),
    .y(_056_)
  );
  al_nand3ftt _390_ (
    .a(_055_),
    .b(_281_),
    .c(_056_),
    .y(_057_)
  );
  al_aoi21ttf _391_ (
    .a(G4),
    .b(G6),
    .c(G5),
    .y(_058_)
  );
  al_oai21ttf _392_ (
    .a(G4),
    .b(G6),
    .c(G3),
    .y(_059_)
  );
  al_and3fft _393_ (
    .a(G3),
    .b(G5),
    .c(G4),
    .y(_060_)
  );
  al_aoi21 _394_ (
    .a(_058_),
    .b(_059_),
    .c(_060_),
    .y(_061_)
  );
  al_ao21ttf _395_ (
    .a(G6),
    .b(_057_),
    .c(_061_),
    .y(_062_)
  );
  al_inv _396_ (
    .a(G6),
    .y(_063_)
  );
  al_and2 _397_ (
    .a(G1),
    .b(G4),
    .y(_064_)
  );
  al_ao21ttf _398_ (
    .a(G2),
    .b(_064_),
    .c(_028_),
    .y(_065_)
  );
  al_and3ftt _399_ (
    .a(G1),
    .b(G2),
    .c(_266_),
    .y(_066_)
  );
  al_ao21 _400_ (
    .a(_063_),
    .b(_065_),
    .c(_066_),
    .y(_067_)
  );
  al_ao21 _401_ (
    .a(G1),
    .b(_062_),
    .c(_067_),
    .y(_068_)
  );
  al_aoi21 _402_ (
    .a(_051_),
    .b(_068_),
    .c(_054_),
    .y(_069_)
  );
  al_nand3fft _403_ (
    .a(G1),
    .b(G6),
    .c(_044_),
    .y(_070_)
  );
  al_nand2 _404_ (
    .a(G11),
    .b(_271_),
    .y(_071_)
  );
  al_aoi21ftt _405_ (
    .a(G8),
    .b(_070_),
    .c(_071_),
    .y(_072_)
  );
  al_and3 _406_ (
    .a(G9),
    .b(G11),
    .c(_016_),
    .y(_073_)
  );
  al_and2ft _407_ (
    .a(G1),
    .b(_268_),
    .y(_074_)
  );
  al_and2ft _408_ (
    .a(G10),
    .b(_285_),
    .y(_075_)
  );
  al_ao21 _409_ (
    .a(_074_),
    .b(_075_),
    .c(_073_),
    .y(_076_)
  );
  al_ao21 _410_ (
    .a(_015_),
    .b(_076_),
    .c(_072_),
    .y(_077_)
  );
  al_or3 _411_ (
    .a(G8),
    .b(_071_),
    .c(_070_),
    .y(_078_)
  );
  al_and3ftt _412_ (
    .a(G4),
    .b(G1),
    .c(G3),
    .y(_079_)
  );
  al_aoi21ftt _413_ (
    .a(_063_),
    .b(_079_),
    .c(_074_),
    .y(_080_)
  );
  al_aoi21 _414_ (
    .a(_078_),
    .b(_080_),
    .c(_279_),
    .y(_081_)
  );
  al_ao21ttf _415_ (
    .a(_285_),
    .b(_042_),
    .c(_030_),
    .y(_082_)
  );
  al_and3 _416_ (
    .a(_041_),
    .b(_283_),
    .c(_082_),
    .y(_083_)
  );
  al_ao21 _417_ (
    .a(_081_),
    .b(_077_),
    .c(_083_),
    .y(_084_)
  );
  al_ao21ttf _418_ (
    .a(_069_),
    .b(_084_),
    .c(_053_),
    .y(_085_)
  );
  al_ao21 _419_ (
    .a(_282_),
    .b(_085_),
    .c(_023_),
    .y(\DFF_16.D )
  );
  al_and3fft _420_ (
    .a(G13),
    .b(_021_),
    .c(G12),
    .y(_086_)
  );
  al_nand2 _421_ (
    .a(G6),
    .b(_086_),
    .y(_087_)
  );
  al_nand2 _422_ (
    .a(G8),
    .b(\DFF_5.Q ),
    .y(_088_)
  );
  al_ao21 _423_ (
    .a(_088_),
    .b(_087_),
    .c(_049_),
    .y(_089_)
  );
  al_oai21ftt _424_ (
    .a(G7),
    .b(G8),
    .c(G11),
    .y(_090_)
  );
  al_nand3fft _425_ (
    .a(G9),
    .b(_029_),
    .c(_090_),
    .y(_091_)
  );
  al_nand2 _426_ (
    .a(G7),
    .b(G9),
    .y(_092_)
  );
  al_nand3 _427_ (
    .a(G8),
    .b(G10),
    .c(_092_),
    .y(_093_)
  );
  al_nand3ftt _428_ (
    .a(_073_),
    .b(_091_),
    .c(_093_),
    .y(_094_)
  );
  al_nand3 _429_ (
    .a(G6),
    .b(_094_),
    .c(_086_),
    .y(_095_)
  );
  al_and3 _430_ (
    .a(G7),
    .b(G10),
    .c(\DFF_5.Q ),
    .y(_096_)
  );
  al_ao21ttf _431_ (
    .a(G8),
    .b(G9),
    .c(_096_),
    .y(_097_)
  );
  al_nand3 _432_ (
    .a(_095_),
    .b(_097_),
    .c(_089_),
    .y(G542)
  );
  al_nand2ft _433_ (
    .a(G5),
    .b(G4),
    .y(_098_)
  );
  al_nand3ftt _434_ (
    .a(G2),
    .b(G3),
    .c(_098_),
    .y(_099_)
  );
  al_nand2ft _435_ (
    .a(G1),
    .b(G2),
    .y(_100_)
  );
  al_mux2l _436_ (
    .a(G3),
    .b(G5),
    .s(G4),
    .y(_101_)
  );
  al_aoi21ftf _437_ (
    .a(_100_),
    .b(_101_),
    .c(_099_),
    .y(\DFF_0.D )
  );
  al_nand3ftt _438_ (
    .a(G5),
    .b(G2),
    .c(G4),
    .y(_102_)
  );
  al_and3 _439_ (
    .a(_282_),
    .b(\DFF_3.Q ),
    .c(_051_),
    .y(_103_)
  );
  al_and3ftt _440_ (
    .a(G4),
    .b(G0),
    .c(G1),
    .y(_104_)
  );
  al_or3fft _441_ (
    .a(G12),
    .b(_104_),
    .c(_021_),
    .y(_105_)
  );
  al_aoi21ftf _442_ (
    .a(_102_),
    .b(_103_),
    .c(_105_),
    .y(\DFF_4.D )
  );
  al_nand2ft _443_ (
    .a(G12),
    .b(G13),
    .y(_106_)
  );
  al_ao21ftt _444_ (
    .a(_106_),
    .b(_051_),
    .c(_103_),
    .y(_107_)
  );
  al_oa21ftt _445_ (
    .a(G13),
    .b(_068_),
    .c(_107_),
    .y(\DFF_5.D )
  );
  al_nand3fft _446_ (
    .a(G7),
    .b(G8),
    .c(_029_),
    .y(_108_)
  );
  al_oa21ftf _447_ (
    .a(_108_),
    .b(_286_),
    .c(G5),
    .y(\DFF_7.D )
  );
  al_ao21ftf _448_ (
    .a(G10),
    .b(_285_),
    .c(_013_),
    .y(_109_)
  );
  al_and3 _449_ (
    .a(G7),
    .b(G8),
    .c(_002_),
    .y(_110_)
  );
  al_ao21ftf _450_ (
    .a(_018_),
    .b(G6),
    .c(_110_),
    .y(_111_)
  );
  al_aoi21ftf _451_ (
    .a(_063_),
    .b(_109_),
    .c(_111_),
    .y(\DFF_11.D )
  );
  al_and2 _452_ (
    .a(G6),
    .b(G9),
    .y(_112_)
  );
  al_nand3ftt _453_ (
    .a(_112_),
    .b(_042_),
    .c(_086_),
    .y(_113_)
  );
  al_inv _454_ (
    .a(\DFF_5.Q ),
    .y(_114_)
  );
  al_or2 _455_ (
    .a(_114_),
    .b(_093_),
    .y(_115_)
  );
  al_and3 _456_ (
    .a(_113_),
    .b(_115_),
    .c(_089_),
    .y(\DFF_12.D )
  );
  al_or3fft _457_ (
    .a(G8),
    .b(G10),
    .c(_278_),
    .y(_116_)
  );
  al_aoi21ftf _458_ (
    .a(_042_),
    .b(_112_),
    .c(_116_),
    .y(_117_)
  );
  al_oai21 _459_ (
    .a(G8),
    .b(G9),
    .c(G6),
    .y(_118_)
  );
  al_or3fft _460_ (
    .a(G7),
    .b(_118_),
    .c(_024_),
    .y(_119_)
  );
  al_ao21 _461_ (
    .a(_119_),
    .b(_117_),
    .c(_001_),
    .y(\DFF_13.D )
  );
  al_and2 _462_ (
    .a(G1),
    .b(G3),
    .y(_120_)
  );
  al_oai21ttf _463_ (
    .a(G2),
    .b(G6),
    .c(_098_),
    .y(_121_)
  );
  al_ao21ftf _464_ (
    .a(_058_),
    .b(_121_),
    .c(_120_),
    .y(_122_)
  );
  al_or3fft _465_ (
    .a(G3),
    .b(_266_),
    .c(_100_),
    .y(_123_)
  );
  al_nand3 _466_ (
    .a(G1),
    .b(G6),
    .c(_055_),
    .y(_124_)
  );
  al_and3 _467_ (
    .a(_124_),
    .b(_123_),
    .c(_122_),
    .y(\DFF_14.D )
  );
  al_or3 _468_ (
    .a(G4),
    .b(G5),
    .c(G6),
    .y(_125_)
  );
  al_inv _469_ (
    .a(_273_),
    .y(_126_)
  );
  al_or3 _470_ (
    .a(G5),
    .b(G6),
    .c(_012_),
    .y(_127_)
  );
  al_nand2ft _471_ (
    .a(_274_),
    .b(_038_),
    .y(_128_)
  );
  al_ao21 _472_ (
    .a(_127_),
    .b(_128_),
    .c(_126_),
    .y(_129_)
  );
  al_aoi21ftf _473_ (
    .a(_125_),
    .b(_286_),
    .c(_129_),
    .y(\DFF_15.D )
  );
  al_ao21ftt _474_ (
    .a(G2),
    .b(G3),
    .c(_098_),
    .y(_130_)
  );
  al_ao21ttf _475_ (
    .a(_098_),
    .b(_009_),
    .c(_130_),
    .y(_131_)
  );
  al_ao21 _476_ (
    .a(G0),
    .b(_131_),
    .c(G1),
    .y(_132_)
  );
  al_aoi21 _477_ (
    .a(G7),
    .b(G10),
    .c(G6),
    .y(_133_)
  );
  al_ao21ttf _478_ (
    .a(\DFF_1.Q ),
    .b(G7),
    .c(_133_),
    .y(_134_)
  );
  al_ao21 _479_ (
    .a(G0),
    .b(_056_),
    .c(_044_),
    .y(_135_)
  );
  al_aoi21ftt _480_ (
    .a(G1),
    .b(G5),
    .c(_079_),
    .y(_136_)
  );
  al_nand3 _481_ (
    .a(G2),
    .b(_136_),
    .c(_135_),
    .y(_137_)
  );
  al_and3 _482_ (
    .a(_134_),
    .b(_137_),
    .c(_132_),
    .y(\DFF_17.D )
  );
  al_inv _483_ (
    .a(\DFF_12.Q ),
    .y(G546)
  );
  al_and3fft _484_ (
    .a(G0),
    .b(G4),
    .c(_291_),
    .y(\DFF_9.D )
  );
  al_inv _485_ (
    .a(G3),
    .y(_138_)
  );
  al_and2 _486_ (
    .a(_138_),
    .b(_039_),
    .y(_139_)
  );
  al_aoi21 _487_ (
    .a(_034_),
    .b(_047_),
    .c(_052_),
    .y(_140_)
  );
  al_and3 _488_ (
    .a(_040_),
    .b(_282_),
    .c(_140_),
    .y(_141_)
  );
  al_nand3 _489_ (
    .a(G0),
    .b(_056_),
    .c(_136_),
    .y(_142_)
  );
  al_and2 _490_ (
    .a(G0),
    .b(G2),
    .y(_143_)
  );
  al_ao21 _491_ (
    .a(_010_),
    .b(_283_),
    .c(_143_),
    .y(_144_)
  );
  al_and3 _492_ (
    .a(_142_),
    .b(_144_),
    .c(_086_),
    .y(_145_)
  );
  al_ao21 _493_ (
    .a(_139_),
    .b(_141_),
    .c(_145_),
    .y(G530)
  );
  al_inv _494_ (
    .a(_268_),
    .y(_146_)
  );
  al_nand3fft _495_ (
    .a(G2),
    .b(_146_),
    .c(_140_),
    .y(_147_)
  );
  al_nand3 _496_ (
    .a(_074_),
    .b(_084_),
    .c(_069_),
    .y(_148_)
  );
  al_nand3ftt _497_ (
    .a(G8),
    .b(G9),
    .c(G11),
    .y(_149_)
  );
  al_or3fft _498_ (
    .a(G10),
    .b(_289_),
    .c(_149_),
    .y(_150_)
  );
  al_ao21 _499_ (
    .a(_148_),
    .b(_147_),
    .c(_150_),
    .y(_151_)
  );
  al_nand2 _500_ (
    .a(G3),
    .b(G5),
    .y(_152_)
  );
  al_nor3fft _501_ (
    .a(G2),
    .b(_064_),
    .c(_152_),
    .y(_153_)
  );
  al_and3 _502_ (
    .a(G6),
    .b(_153_),
    .c(_082_),
    .y(_154_)
  );
  al_aoi21 _503_ (
    .a(_081_),
    .b(_077_),
    .c(_154_),
    .y(_155_)
  );
  al_or3fft _504_ (
    .a(G1),
    .b(_069_),
    .c(_155_),
    .y(_156_)
  );
  al_nor2 _505_ (
    .a(G4),
    .b(G5),
    .y(_157_)
  );
  al_and3 _506_ (
    .a(G3),
    .b(G6),
    .c(_157_),
    .y(_158_)
  );
  al_and3 _507_ (
    .a(G2),
    .b(G11),
    .c(_158_),
    .y(_159_)
  );
  al_aoi21 _508_ (
    .a(_276_),
    .b(_159_),
    .c(_031_),
    .y(_160_)
  );
  al_ao21 _509_ (
    .a(_053_),
    .b(_156_),
    .c(_160_),
    .y(_161_)
  );
  al_and2ft _510_ (
    .a(\DFF_14.Q ),
    .b(G13),
    .y(_162_)
  );
  al_and3 _511_ (
    .a(_051_),
    .b(_162_),
    .c(_068_),
    .y(_163_)
  );
  al_nand3 _512_ (
    .a(G8),
    .b(_271_),
    .c(_038_),
    .y(_164_)
  );
  al_nand3fft _513_ (
    .a(G4),
    .b(G6),
    .c(\DFF_7.Q ),
    .y(_165_)
  );
  al_aoi21ttf _514_ (
    .a(_165_),
    .b(_164_),
    .c(_035_),
    .y(_166_)
  );
  al_aoi21 _515_ (
    .a(_166_),
    .b(_140_),
    .c(_163_),
    .y(_167_)
  );
  al_nand3 _516_ (
    .a(_167_),
    .b(_161_),
    .c(_151_),
    .y(_168_)
  );
  al_ao21ttf _517_ (
    .a(G1),
    .b(G3),
    .c(G2),
    .y(_169_)
  );
  al_aoi21ttf _518_ (
    .a(_280_),
    .b(_169_),
    .c(G4),
    .y(_170_)
  );
  al_and3fft _519_ (
    .a(G2),
    .b(G3),
    .c(G5),
    .y(_171_)
  );
  al_ao21 _520_ (
    .a(G1),
    .b(_171_),
    .c(_060_),
    .y(_172_)
  );
  al_or3 _521_ (
    .a(_079_),
    .b(_172_),
    .c(_170_),
    .y(_173_)
  );
  al_and3 _522_ (
    .a(G0),
    .b(_173_),
    .c(_086_),
    .y(_174_)
  );
  al_ao21 _523_ (
    .a(_282_),
    .b(_168_),
    .c(_174_),
    .y(G532)
  );
  al_or3fft _524_ (
    .a(_268_),
    .b(_032_),
    .c(_026_),
    .y(_175_)
  );
  al_aoi21ftf _525_ (
    .a(\DFF_15.Q ),
    .b(_138_),
    .c(_175_),
    .y(_176_)
  );
  al_nand3 _526_ (
    .a(G1),
    .b(_292_),
    .c(_023_),
    .y(_177_)
  );
  al_or3fft _527_ (
    .a(\DFF_9.Q ),
    .b(\DFF_8.Q ),
    .c(_177_),
    .y(_178_)
  );
  al_aoi21ftf _528_ (
    .a(_176_),
    .b(_141_),
    .c(_178_),
    .y(_179_)
  );
  al_and3ftt _529_ (
    .a(G12),
    .b(G3),
    .c(G6),
    .y(_180_)
  );
  al_nand3fft _530_ (
    .a(G4),
    .b(G5),
    .c(_276_),
    .y(_181_)
  );
  al_ao21 _531_ (
    .a(_053_),
    .b(_156_),
    .c(_181_),
    .y(_182_)
  );
  al_or3 _532_ (
    .a(G1),
    .b(_098_),
    .c(_026_),
    .y(_183_)
  );
  al_nand3ftt _533_ (
    .a(_183_),
    .b(_084_),
    .c(_069_),
    .y(_184_)
  );
  al_nand2 _534_ (
    .a(_184_),
    .b(_182_),
    .y(_185_)
  );
  al_ao21ttf _535_ (
    .a(_180_),
    .b(_185_),
    .c(_179_),
    .y(G535)
  );
  al_nand2 _536_ (
    .a(_053_),
    .b(_156_),
    .y(_186_)
  );
  al_and3 _537_ (
    .a(G7),
    .b(G9),
    .c(G10),
    .y(_187_)
  );
  al_nand3 _538_ (
    .a(_292_),
    .b(_037_),
    .c(_187_),
    .y(_188_)
  );
  al_aoi21ftf _539_ (
    .a(_275_),
    .b(_158_),
    .c(_188_),
    .y(_189_)
  );
  al_inv _540_ (
    .a(G5),
    .y(_190_)
  );
  al_or3fft _541_ (
    .a(_190_),
    .b(_276_),
    .c(_148_),
    .y(_191_)
  );
  al_ao21ftf _542_ (
    .a(_189_),
    .b(_186_),
    .c(_191_),
    .y(_192_)
  );
  al_nand3 _543_ (
    .a(_268_),
    .b(_032_),
    .c(_276_),
    .y(_193_)
  );
  al_ao21ftf _544_ (
    .a(_125_),
    .b(_029_),
    .c(_128_),
    .y(_194_)
  );
  al_nand3fft _545_ (
    .a(G3),
    .b(_126_),
    .c(_194_),
    .y(_195_)
  );
  al_nand3 _546_ (
    .a(_063_),
    .b(_060_),
    .c(_286_),
    .y(_196_)
  );
  al_nand3 _547_ (
    .a(_196_),
    .b(_193_),
    .c(_195_),
    .y(_197_)
  );
  al_oai21ftf _548_ (
    .a(\DFF_9.Q ),
    .b(_278_),
    .c(G0),
    .y(_198_)
  );
  al_or2ft _549_ (
    .a(_198_),
    .b(_177_),
    .y(_199_)
  );
  al_ao21ttf _550_ (
    .a(_141_),
    .b(_197_),
    .c(_199_),
    .y(_200_)
  );
  al_ao21 _551_ (
    .a(_282_),
    .b(_192_),
    .c(_200_),
    .y(G537)
  );
  al_or2 _552_ (
    .a(G12),
    .b(_052_),
    .y(_201_)
  );
  al_nand3ftt _553_ (
    .a(_201_),
    .b(_034_),
    .c(_047_),
    .y(_202_)
  );
  al_nand2 _554_ (
    .a(_051_),
    .b(_068_),
    .y(_203_)
  );
  al_inv _555_ (
    .a(_106_),
    .y(_204_)
  );
  al_nand3 _556_ (
    .a(_204_),
    .b(_203_),
    .c(_155_),
    .y(_205_)
  );
  al_nand3ftt _557_ (
    .a(_000_),
    .b(_022_),
    .c(_021_),
    .y(_206_)
  );
  al_nand3 _558_ (
    .a(_206_),
    .b(_202_),
    .c(_205_),
    .y(G539)
  );
  al_ao21ttf _559_ (
    .a(G8),
    .b(G10),
    .c(G7),
    .y(_207_)
  );
  al_oai21ftt _560_ (
    .a(G10),
    .b(_025_),
    .c(_207_),
    .y(_208_)
  );
  al_nand3 _561_ (
    .a(G9),
    .b(\DFF_5.Q ),
    .c(_208_),
    .y(_209_)
  );
  al_nand2ft _562_ (
    .a(G9),
    .b(G10),
    .y(_210_)
  );
  al_nand3fft _563_ (
    .a(_025_),
    .b(_029_),
    .c(_210_),
    .y(_211_)
  );
  al_nand3ftt _564_ (
    .a(G10),
    .b(G9),
    .c(_025_),
    .y(_212_)
  );
  al_nand3 _565_ (
    .a(_149_),
    .b(_212_),
    .c(_211_),
    .y(_213_)
  );
  al_mux2h _566_ (
    .a(_187_),
    .b(_213_),
    .s(G6),
    .y(_214_)
  );
  al_ao21ttf _567_ (
    .a(_214_),
    .b(_086_),
    .c(_209_),
    .y(G547)
  );
  al_or3fft _568_ (
    .a(G9),
    .b(G11),
    .c(_207_),
    .y(_215_)
  );
  al_ao21ftf _569_ (
    .a(G9),
    .b(_042_),
    .c(_025_),
    .y(_216_)
  );
  al_nand3fft _570_ (
    .a(_001_),
    .b(_024_),
    .c(_216_),
    .y(_217_)
  );
  al_ao21 _571_ (
    .a(_215_),
    .b(_217_),
    .c(_114_),
    .y(_218_)
  );
  al_ao21ftf _572_ (
    .a(\DFF_13.Q ),
    .b(_086_),
    .c(_218_),
    .y(G548)
  );
  al_nand2 _573_ (
    .a(G0),
    .b(G3),
    .y(_219_)
  );
  al_nand3 _574_ (
    .a(_064_),
    .b(_219_),
    .c(_086_),
    .y(_220_)
  );
  al_and3 _575_ (
    .a(G1),
    .b(_051_),
    .c(_068_),
    .y(_221_)
  );
  al_nand3 _576_ (
    .a(G6),
    .b(_281_),
    .c(_152_),
    .y(_222_)
  );
  al_oai21ttf _577_ (
    .a(G5),
    .b(G6),
    .c(G4),
    .y(_223_)
  );
  al_and3ftt _578_ (
    .a(G3),
    .b(G4),
    .c(G6),
    .y(_224_)
  );
  al_nand2 _579_ (
    .a(G5),
    .b(_224_),
    .y(_225_)
  );
  al_and3 _580_ (
    .a(_102_),
    .b(_280_),
    .c(_225_),
    .y(_226_)
  );
  al_ao21ftf _581_ (
    .a(_223_),
    .b(_222_),
    .c(_226_),
    .y(_227_)
  );
  al_nand3 _582_ (
    .a(_204_),
    .b(_227_),
    .c(_221_),
    .y(_228_)
  );
  al_or3ftt _583_ (
    .a(G3),
    .b(\DFF_4.Q ),
    .c(G13),
    .y(_229_)
  );
  al_and2 _584_ (
    .a(_054_),
    .b(_103_),
    .y(_230_)
  );
  al_aoi21 _585_ (
    .a(G3),
    .b(G4),
    .c(_028_),
    .y(_231_)
  );
  al_aoi21ttf _586_ (
    .a(_231_),
    .b(_230_),
    .c(_229_),
    .y(_232_)
  );
  al_nand3 _587_ (
    .a(_228_),
    .b(_232_),
    .c(_220_),
    .y(G549)
  );
  al_and3ftt _588_ (
    .a(\DFF_0.Q ),
    .b(G0),
    .c(_086_),
    .y(_233_)
  );
  al_nand2 _589_ (
    .a(G4),
    .b(G5),
    .y(_234_)
  );
  al_oa21ftf _590_ (
    .a(G1),
    .b(_234_),
    .c(_106_),
    .y(_235_)
  );
  al_nor3fft _591_ (
    .a(_065_),
    .b(_235_),
    .c(_203_),
    .y(_236_)
  );
  al_and2 _592_ (
    .a(G2),
    .b(G4),
    .y(_237_)
  );
  al_nand3fft _593_ (
    .a(_152_),
    .b(_237_),
    .c(_230_),
    .y(_238_)
  );
  al_and3ftt _594_ (
    .a(G0),
    .b(G1),
    .c(G4),
    .y(_239_)
  );
  al_nand3 _595_ (
    .a(G3),
    .b(_239_),
    .c(_086_),
    .y(_240_)
  );
  al_and3 _596_ (
    .a(_229_),
    .b(_238_),
    .c(_240_),
    .y(_241_)
  );
  al_nand3fft _597_ (
    .a(_233_),
    .b(_236_),
    .c(_241_),
    .y(G550)
  );
  al_nand3ftt _598_ (
    .a(G5),
    .b(G6),
    .c(_055_),
    .y(_242_)
  );
  al_and3ftt _599_ (
    .a(_224_),
    .b(_242_),
    .c(_130_),
    .y(_243_)
  );
  al_and3ftt _600_ (
    .a(G1),
    .b(G2),
    .c(G4),
    .y(_244_)
  );
  al_ao21 _601_ (
    .a(_055_),
    .b(_064_),
    .c(_244_),
    .y(_245_)
  );
  al_or3fft _602_ (
    .a(G5),
    .b(_245_),
    .c(_203_),
    .y(_246_)
  );
  al_ao21ftf _603_ (
    .a(_243_),
    .b(_221_),
    .c(_246_),
    .y(_247_)
  );
  al_ao21ttf _604_ (
    .a(G0),
    .b(G2),
    .c(G1),
    .y(_248_)
  );
  al_nand3 _605_ (
    .a(G0),
    .b(G2),
    .c(G4),
    .y(_249_)
  );
  al_ao21 _606_ (
    .a(_248_),
    .b(_249_),
    .c(G3),
    .y(_250_)
  );
  al_mux2l _607_ (
    .a(G0),
    .b(_219_),
    .s(_064_),
    .y(_251_)
  );
  al_aoi21 _608_ (
    .a(_250_),
    .b(_251_),
    .c(_190_),
    .y(_252_)
  );
  al_and3 _609_ (
    .a(G4),
    .b(\DFF_10.Q ),
    .c(_230_),
    .y(_253_)
  );
  al_aoi21 _610_ (
    .a(_252_),
    .b(_086_),
    .c(_253_),
    .y(_254_)
  );
  al_ao21ttf _611_ (
    .a(_204_),
    .b(_247_),
    .c(_254_),
    .y(G551)
  );
  al_oai21ftt _612_ (
    .a(G5),
    .b(G1),
    .c(G4),
    .y(_255_)
  );
  al_nand3ftt _613_ (
    .a(G4),
    .b(G5),
    .c(_120_),
    .y(_256_)
  );
  al_aoi21ttf _614_ (
    .a(_028_),
    .b(_064_),
    .c(_256_),
    .y(_257_)
  );
  al_ao21ftf _615_ (
    .a(_169_),
    .b(_255_),
    .c(_257_),
    .y(_258_)
  );
  al_or3fft _616_ (
    .a(_204_),
    .b(_258_),
    .c(_203_),
    .y(_259_)
  );
  al_ao21ftf _617_ (
    .a(_270_),
    .b(_234_),
    .c(_099_),
    .y(_260_)
  );
  al_and2 _618_ (
    .a(G2),
    .b(_224_),
    .y(_261_)
  );
  al_ao21 _619_ (
    .a(G6),
    .b(_260_),
    .c(_261_),
    .y(_262_)
  );
  al_nand3 _620_ (
    .a(_054_),
    .b(_262_),
    .c(_103_),
    .y(_263_)
  );
  al_aoi21ftf _621_ (
    .a(\DFF_11.Q ),
    .b(_086_),
    .c(_263_),
    .y(_264_)
  );
  al_ao21ftf _622_ (
    .a(_259_),
    .b(G6),
    .c(_264_),
    .y(G552)
  );
  al_dffl _623_ (
    .clk(CK),
    .d(\DFF_0.D ),
    .q(\DFF_0.Q )
  );
  al_dffl _624_ (
    .clk(CK),
    .d(\DFF_1.D ),
    .q(\DFF_1.Q )
  );
  al_dffl _625_ (
    .clk(CK),
    .d(\DFF_2.D ),
    .q(\DFF_2.Q )
  );
  al_dffl _626_ (
    .clk(CK),
    .d(\DFF_3.D ),
    .q(\DFF_3.Q )
  );
  al_dffl _627_ (
    .clk(CK),
    .d(\DFF_4.D ),
    .q(\DFF_4.Q )
  );
  al_dffl _628_ (
    .clk(CK),
    .d(\DFF_5.D ),
    .q(\DFF_5.Q )
  );
  al_dffl _629_ (
    .clk(CK),
    .d(\DFF_6.D ),
    .q(\DFF_6.Q )
  );
  al_dffl _630_ (
    .clk(CK),
    .d(\DFF_7.D ),
    .q(\DFF_7.Q )
  );
  al_dffl _631_ (
    .clk(CK),
    .d(\DFF_8.D ),
    .q(\DFF_8.Q )
  );
  al_dffl _632_ (
    .clk(CK),
    .d(\DFF_9.D ),
    .q(\DFF_9.Q )
  );
  al_dffl _633_ (
    .clk(CK),
    .d(\DFF_10.D ),
    .q(\DFF_10.Q )
  );
  al_dffl _634_ (
    .clk(CK),
    .d(\DFF_11.D ),
    .q(\DFF_11.Q )
  );
  al_dffl _635_ (
    .clk(CK),
    .d(\DFF_12.D ),
    .q(\DFF_12.Q )
  );
  al_dffl _636_ (
    .clk(CK),
    .d(\DFF_13.D ),
    .q(\DFF_13.Q )
  );
  al_dffl _637_ (
    .clk(CK),
    .d(\DFF_14.D ),
    .q(\DFF_14.Q )
  );
  al_dffl _638_ (
    .clk(CK),
    .d(\DFF_15.D ),
    .q(\DFF_15.Q )
  );
  al_dffl _639_ (
    .clk(CK),
    .d(\DFF_16.D ),
    .q(\DFF_16.Q )
  );
  al_dffl _640_ (
    .clk(CK),
    .d(\DFF_17.D ),
    .q(\DFF_17.Q )
  );
  assign \DFF_0.CK  = CK;
  assign \DFF_1.CK  = CK;
  assign \DFF_10.CK  = CK;
  assign \DFF_11.CK  = CK;
  assign \DFF_12.CK  = CK;
  assign \DFF_13.CK  = CK;
  assign \DFF_14.CK  = CK;
  assign \DFF_15.CK  = CK;
  assign \DFF_16.CK  = CK;
  assign \DFF_17.CK  = CK;
  assign \DFF_2.CK  = CK;
  assign \DFF_3.CK  = CK;
  assign \DFF_4.CK  = CK;
  assign \DFF_5.CK  = CK;
  assign \DFF_6.CK  = CK;
  assign \DFF_7.CK  = CK;
  assign \DFF_8.CK  = CK;
  assign \DFF_9.CK  = CK;
  assign G29 = \DFF_0.Q ;
  assign G30 = \DFF_1.Q ;
  assign G31 = \DFF_2.Q ;
  assign G32 = \DFF_3.Q ;
  assign G33 = \DFF_4.Q ;
  assign G34 = \DFF_5.Q ;
  assign G35 = \DFF_6.Q ;
  assign G36 = \DFF_7.Q ;
  assign G37 = \DFF_8.Q ;
  assign G38 = \DFF_9.Q ;
  assign G39 = \DFF_10.Q ;
  assign G40 = \DFF_11.Q ;
  assign G41 = \DFF_12.Q ;
  assign G42 = \DFF_13.Q ;
  assign G43 = \DFF_14.Q ;
  assign G44 = \DFF_15.Q ;
  assign G45 = \DFF_16.Q ;
  assign G46 = \DFF_17.Q ;
  assign G502 = \DFF_0.D ;
  assign G503 = \DFF_1.D ;
  assign G504 = \DFF_2.D ;
  assign G505 = \DFF_3.D ;
  assign G506 = \DFF_4.D ;
  assign G507 = \DFF_5.D ;
  assign G508 = \DFF_6.D ;
  assign G509 = \DFF_7.D ;
  assign G510 = \DFF_8.D ;
  assign G511 = \DFF_9.D ;
  assign G512 = \DFF_10.D ;
  assign G513 = \DFF_11.D ;
  assign G514 = \DFF_12.D ;
  assign G515 = \DFF_13.D ;
  assign G516 = \DFF_14.D ;
  assign G517 = \DFF_15.D ;
  assign G518 = \DFF_16.D ;
  assign G519 = \DFF_17.D ;
endmodule
