
module s5378(GND, VDD, CK, n3065gat, n3066gat, n3067gat, n3068gat, n3069gat, n3070gat, n3071gat, n3072gat, n3073gat, n3074gat, n3075gat, n3076gat, n3077gat, n3078gat, n3079gat, n3080gat, n3081gat, n3082gat, n3083gat, n3084gat, n3085gat, n3086gat, n3087gat, n3088gat, n3089gat, n3090gat, n3091gat, n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat, n3099gat, n3100gat, n3104gat, n3105gat, n3106gat, n3107gat, n3108gat, n3109gat, n3110gat, n3111gat, n3112gat, n3113gat, n3114gat, n3115gat, n3116gat, n3117gat, n3118gat, n3119gat, n3120gat, n3121gat, n3122gat, n3123gat, n3124gat, n3125gat, n3126gat, n3127gat, n3128gat, n3129gat, n3130gat, n3131gat, n3132gat, n3133gat, n3134gat, n3135gat, n3136gat, n3137gat, n3138gat, n3139gat, n3140gat, n3141gat, n3142gat, n3143gat, n3144gat, n3145gat, n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, n3151gat, n3152gat);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  input CK;
  wire \DFF_0.CK ;
  wire \DFF_0.D ;
  wire \DFF_0.Q ;
  wire \DFF_1.CK ;
  wire \DFF_1.D ;
  wire \DFF_1.Q ;
  wire \DFF_10.CK ;
  wire \DFF_10.D ;
  wire \DFF_10.Q ;
  wire \DFF_100.CK ;
  wire \DFF_100.D ;
  wire \DFF_100.Q ;
  wire \DFF_101.CK ;
  wire \DFF_101.D ;
  wire \DFF_101.Q ;
  wire \DFF_102.CK ;
  wire \DFF_102.D ;
  wire \DFF_102.Q ;
  wire \DFF_103.CK ;
  wire \DFF_103.D ;
  wire \DFF_103.Q ;
  wire \DFF_104.CK ;
  wire \DFF_104.D ;
  wire \DFF_104.Q ;
  wire \DFF_105.CK ;
  wire \DFF_105.D ;
  wire \DFF_105.Q ;
  wire \DFF_106.CK ;
  wire \DFF_106.D ;
  wire \DFF_106.Q ;
  wire \DFF_107.CK ;
  wire \DFF_107.D ;
  wire \DFF_107.Q ;
  wire \DFF_108.CK ;
  wire \DFF_108.D ;
  wire \DFF_108.Q ;
  wire \DFF_109.CK ;
  wire \DFF_109.D ;
  wire \DFF_109.Q ;
  wire \DFF_11.CK ;
  wire \DFF_11.D ;
  wire \DFF_11.Q ;
  wire \DFF_110.CK ;
  wire \DFF_110.D ;
  wire \DFF_110.Q ;
  wire \DFF_111.CK ;
  wire \DFF_111.D ;
  wire \DFF_111.Q ;
  wire \DFF_112.CK ;
  wire \DFF_112.D ;
  wire \DFF_112.Q ;
  wire \DFF_113.CK ;
  wire \DFF_113.D ;
  wire \DFF_113.Q ;
  wire \DFF_114.CK ;
  wire \DFF_114.D ;
  wire \DFF_114.Q ;
  wire \DFF_115.CK ;
  wire \DFF_115.D ;
  wire \DFF_115.Q ;
  wire \DFF_116.CK ;
  wire \DFF_116.D ;
  wire \DFF_116.Q ;
  wire \DFF_117.CK ;
  wire \DFF_117.D ;
  wire \DFF_117.Q ;
  wire \DFF_118.CK ;
  wire \DFF_118.D ;
  wire \DFF_118.Q ;
  wire \DFF_119.CK ;
  wire \DFF_119.D ;
  wire \DFF_119.Q ;
  wire \DFF_12.CK ;
  wire \DFF_12.D ;
  wire \DFF_12.Q ;
  wire \DFF_120.CK ;
  wire \DFF_120.D ;
  wire \DFF_120.Q ;
  wire \DFF_121.CK ;
  wire \DFF_121.D ;
  wire \DFF_121.Q ;
  wire \DFF_122.CK ;
  wire \DFF_122.D ;
  wire \DFF_122.Q ;
  wire \DFF_123.CK ;
  wire \DFF_123.D ;
  wire \DFF_123.Q ;
  wire \DFF_124.CK ;
  wire \DFF_124.D ;
  wire \DFF_124.Q ;
  wire \DFF_125.CK ;
  wire \DFF_125.D ;
  wire \DFF_125.Q ;
  wire \DFF_126.CK ;
  wire \DFF_126.D ;
  wire \DFF_126.Q ;
  wire \DFF_127.CK ;
  wire \DFF_127.D ;
  wire \DFF_127.Q ;
  wire \DFF_128.CK ;
  wire \DFF_128.D ;
  wire \DFF_128.Q ;
  wire \DFF_129.CK ;
  wire \DFF_129.D ;
  wire \DFF_129.Q ;
  wire \DFF_13.CK ;
  wire \DFF_13.D ;
  wire \DFF_13.Q ;
  wire \DFF_130.CK ;
  wire \DFF_130.D ;
  wire \DFF_130.Q ;
  wire \DFF_131.CK ;
  wire \DFF_131.D ;
  wire \DFF_131.Q ;
  wire \DFF_132.CK ;
  wire \DFF_132.D ;
  wire \DFF_132.Q ;
  wire \DFF_133.CK ;
  wire \DFF_133.D ;
  wire \DFF_133.Q ;
  wire \DFF_134.CK ;
  wire \DFF_134.D ;
  wire \DFF_134.Q ;
  wire \DFF_135.CK ;
  wire \DFF_135.D ;
  wire \DFF_135.Q ;
  wire \DFF_136.CK ;
  wire \DFF_137.CK ;
  wire \DFF_138.CK ;
  wire \DFF_139.CK ;
  wire \DFF_139.D ;
  wire \DFF_139.Q ;
  wire \DFF_14.CK ;
  wire \DFF_14.D ;
  wire \DFF_14.Q ;
  wire \DFF_140.CK ;
  wire \DFF_140.D ;
  wire \DFF_140.Q ;
  wire \DFF_141.CK ;
  wire \DFF_141.D ;
  wire \DFF_141.Q ;
  wire \DFF_142.CK ;
  wire \DFF_142.D ;
  wire \DFF_142.Q ;
  wire \DFF_143.CK ;
  wire \DFF_143.D ;
  wire \DFF_143.Q ;
  wire \DFF_144.CK ;
  wire \DFF_144.D ;
  wire \DFF_144.Q ;
  wire \DFF_145.CK ;
  wire \DFF_145.D ;
  wire \DFF_145.Q ;
  wire \DFF_146.CK ;
  wire \DFF_146.D ;
  wire \DFF_146.Q ;
  wire \DFF_147.CK ;
  wire \DFF_147.D ;
  wire \DFF_147.Q ;
  wire \DFF_148.CK ;
  wire \DFF_148.D ;
  wire \DFF_148.Q ;
  wire \DFF_149.CK ;
  wire \DFF_149.D ;
  wire \DFF_149.Q ;
  wire \DFF_15.CK ;
  wire \DFF_15.D ;
  wire \DFF_15.Q ;
  wire \DFF_150.CK ;
  wire \DFF_150.D ;
  wire \DFF_150.Q ;
  wire \DFF_151.CK ;
  wire \DFF_151.D ;
  wire \DFF_151.Q ;
  wire \DFF_152.CK ;
  wire \DFF_152.D ;
  wire \DFF_152.Q ;
  wire \DFF_153.CK ;
  wire \DFF_153.D ;
  wire \DFF_153.Q ;
  wire \DFF_154.CK ;
  wire \DFF_154.D ;
  wire \DFF_154.Q ;
  wire \DFF_155.CK ;
  wire \DFF_155.D ;
  wire \DFF_155.Q ;
  wire \DFF_156.CK ;
  wire \DFF_156.D ;
  wire \DFF_156.Q ;
  wire \DFF_157.CK ;
  wire \DFF_157.D ;
  wire \DFF_157.Q ;
  wire \DFF_158.CK ;
  wire \DFF_158.D ;
  wire \DFF_158.Q ;
  wire \DFF_159.CK ;
  wire \DFF_159.D ;
  wire \DFF_159.Q ;
  wire \DFF_16.CK ;
  wire \DFF_16.D ;
  wire \DFF_16.Q ;
  wire \DFF_160.CK ;
  wire \DFF_160.D ;
  wire \DFF_160.Q ;
  wire \DFF_161.CK ;
  wire \DFF_161.D ;
  wire \DFF_161.Q ;
  wire \DFF_162.CK ;
  wire \DFF_162.D ;
  wire \DFF_162.Q ;
  wire \DFF_163.CK ;
  wire \DFF_163.D ;
  wire \DFF_163.Q ;
  wire \DFF_164.CK ;
  wire \DFF_164.D ;
  wire \DFF_164.Q ;
  wire \DFF_165.CK ;
  wire \DFF_165.D ;
  wire \DFF_165.Q ;
  wire \DFF_166.CK ;
  wire \DFF_166.D ;
  wire \DFF_166.Q ;
  wire \DFF_167.CK ;
  wire \DFF_167.D ;
  wire \DFF_167.Q ;
  wire \DFF_168.CK ;
  wire \DFF_168.D ;
  wire \DFF_168.Q ;
  wire \DFF_169.CK ;
  wire \DFF_169.D ;
  wire \DFF_169.Q ;
  wire \DFF_17.CK ;
  wire \DFF_17.D ;
  wire \DFF_17.Q ;
  wire \DFF_170.CK ;
  wire \DFF_170.D ;
  wire \DFF_170.Q ;
  wire \DFF_171.CK ;
  wire \DFF_171.D ;
  wire \DFF_171.Q ;
  wire \DFF_172.CK ;
  wire \DFF_172.D ;
  wire \DFF_172.Q ;
  wire \DFF_173.CK ;
  wire \DFF_173.D ;
  wire \DFF_173.Q ;
  wire \DFF_174.CK ;
  wire \DFF_174.D ;
  wire \DFF_174.Q ;
  wire \DFF_175.CK ;
  wire \DFF_175.D ;
  wire \DFF_175.Q ;
  wire \DFF_176.CK ;
  wire \DFF_176.D ;
  wire \DFF_176.Q ;
  wire \DFF_177.CK ;
  wire \DFF_177.D ;
  wire \DFF_177.Q ;
  wire \DFF_178.CK ;
  wire \DFF_178.D ;
  wire \DFF_178.Q ;
  wire \DFF_18.CK ;
  wire \DFF_18.D ;
  wire \DFF_18.Q ;
  wire \DFF_19.CK ;
  wire \DFF_19.D ;
  wire \DFF_19.Q ;
  wire \DFF_2.CK ;
  wire \DFF_2.D ;
  wire \DFF_2.Q ;
  wire \DFF_20.CK ;
  wire \DFF_20.D ;
  wire \DFF_20.Q ;
  wire \DFF_21.CK ;
  wire \DFF_21.D ;
  wire \DFF_21.Q ;
  wire \DFF_22.CK ;
  wire \DFF_22.D ;
  wire \DFF_22.Q ;
  wire \DFF_23.CK ;
  wire \DFF_23.D ;
  wire \DFF_23.Q ;
  wire \DFF_24.CK ;
  wire \DFF_24.D ;
  wire \DFF_24.Q ;
  wire \DFF_25.CK ;
  wire \DFF_25.D ;
  wire \DFF_25.Q ;
  wire \DFF_26.CK ;
  wire \DFF_26.D ;
  wire \DFF_26.Q ;
  wire \DFF_27.CK ;
  wire \DFF_27.D ;
  wire \DFF_27.Q ;
  wire \DFF_28.CK ;
  wire \DFF_28.D ;
  wire \DFF_28.Q ;
  wire \DFF_29.CK ;
  wire \DFF_29.D ;
  wire \DFF_29.Q ;
  wire \DFF_3.CK ;
  wire \DFF_3.D ;
  wire \DFF_3.Q ;
  wire \DFF_30.CK ;
  wire \DFF_30.D ;
  wire \DFF_30.Q ;
  wire \DFF_31.CK ;
  wire \DFF_31.D ;
  wire \DFF_31.Q ;
  wire \DFF_32.CK ;
  wire \DFF_32.D ;
  wire \DFF_32.Q ;
  wire \DFF_33.CK ;
  wire \DFF_33.D ;
  wire \DFF_33.Q ;
  wire \DFF_34.CK ;
  wire \DFF_34.D ;
  wire \DFF_34.Q ;
  wire \DFF_35.CK ;
  wire \DFF_35.D ;
  wire \DFF_35.Q ;
  wire \DFF_36.CK ;
  wire \DFF_36.D ;
  wire \DFF_36.Q ;
  wire \DFF_37.CK ;
  wire \DFF_37.D ;
  wire \DFF_37.Q ;
  wire \DFF_38.CK ;
  wire \DFF_38.D ;
  wire \DFF_38.Q ;
  wire \DFF_39.CK ;
  wire \DFF_39.D ;
  wire \DFF_39.Q ;
  wire \DFF_4.CK ;
  wire \DFF_4.D ;
  wire \DFF_4.Q ;
  wire \DFF_40.CK ;
  wire \DFF_40.D ;
  wire \DFF_40.Q ;
  wire \DFF_41.CK ;
  wire \DFF_41.D ;
  wire \DFF_41.Q ;
  wire \DFF_42.CK ;
  wire \DFF_42.D ;
  wire \DFF_42.Q ;
  wire \DFF_43.CK ;
  wire \DFF_43.D ;
  wire \DFF_43.Q ;
  wire \DFF_44.CK ;
  wire \DFF_44.D ;
  wire \DFF_44.Q ;
  wire \DFF_45.CK ;
  wire \DFF_45.D ;
  wire \DFF_45.Q ;
  wire \DFF_46.CK ;
  wire \DFF_46.D ;
  wire \DFF_46.Q ;
  wire \DFF_47.CK ;
  wire \DFF_47.D ;
  wire \DFF_47.Q ;
  wire \DFF_48.CK ;
  wire \DFF_48.D ;
  wire \DFF_48.Q ;
  wire \DFF_49.CK ;
  wire \DFF_49.D ;
  wire \DFF_49.Q ;
  wire \DFF_5.CK ;
  wire \DFF_5.D ;
  wire \DFF_5.Q ;
  wire \DFF_50.CK ;
  wire \DFF_50.D ;
  wire \DFF_50.Q ;
  wire \DFF_51.CK ;
  wire \DFF_51.D ;
  wire \DFF_51.Q ;
  wire \DFF_52.CK ;
  wire \DFF_52.D ;
  wire \DFF_52.Q ;
  wire \DFF_53.CK ;
  wire \DFF_53.D ;
  wire \DFF_53.Q ;
  wire \DFF_54.CK ;
  wire \DFF_54.D ;
  wire \DFF_54.Q ;
  wire \DFF_55.CK ;
  wire \DFF_55.D ;
  wire \DFF_55.Q ;
  wire \DFF_56.CK ;
  wire \DFF_56.D ;
  wire \DFF_56.Q ;
  wire \DFF_57.CK ;
  wire \DFF_57.D ;
  wire \DFF_57.Q ;
  wire \DFF_58.CK ;
  wire \DFF_58.D ;
  wire \DFF_58.Q ;
  wire \DFF_59.CK ;
  wire \DFF_59.D ;
  wire \DFF_59.Q ;
  wire \DFF_6.CK ;
  wire \DFF_6.D ;
  wire \DFF_6.Q ;
  wire \DFF_60.CK ;
  wire \DFF_60.D ;
  wire \DFF_60.Q ;
  wire \DFF_61.CK ;
  wire \DFF_61.D ;
  wire \DFF_61.Q ;
  wire \DFF_62.CK ;
  wire \DFF_62.D ;
  wire \DFF_62.Q ;
  wire \DFF_63.CK ;
  wire \DFF_63.D ;
  wire \DFF_63.Q ;
  wire \DFF_64.CK ;
  wire \DFF_64.D ;
  wire \DFF_64.Q ;
  wire \DFF_65.CK ;
  wire \DFF_65.D ;
  wire \DFF_65.Q ;
  wire \DFF_66.CK ;
  wire \DFF_66.D ;
  wire \DFF_66.Q ;
  wire \DFF_67.CK ;
  wire \DFF_67.D ;
  wire \DFF_67.Q ;
  wire \DFF_68.CK ;
  wire \DFF_68.D ;
  wire \DFF_68.Q ;
  wire \DFF_69.CK ;
  wire \DFF_69.D ;
  wire \DFF_69.Q ;
  wire \DFF_7.CK ;
  wire \DFF_7.D ;
  wire \DFF_7.Q ;
  wire \DFF_70.CK ;
  wire \DFF_70.D ;
  wire \DFF_70.Q ;
  wire \DFF_71.CK ;
  wire \DFF_71.D ;
  wire \DFF_71.Q ;
  wire \DFF_72.CK ;
  wire \DFF_72.D ;
  wire \DFF_72.Q ;
  wire \DFF_73.CK ;
  wire \DFF_73.D ;
  wire \DFF_73.Q ;
  wire \DFF_74.CK ;
  wire \DFF_74.D ;
  wire \DFF_74.Q ;
  wire \DFF_75.CK ;
  wire \DFF_75.D ;
  wire \DFF_75.Q ;
  wire \DFF_76.CK ;
  wire \DFF_76.D ;
  wire \DFF_76.Q ;
  wire \DFF_77.CK ;
  wire \DFF_77.D ;
  wire \DFF_77.Q ;
  wire \DFF_78.CK ;
  wire \DFF_78.D ;
  wire \DFF_78.Q ;
  wire \DFF_79.CK ;
  wire \DFF_79.D ;
  wire \DFF_79.Q ;
  wire \DFF_8.CK ;
  wire \DFF_8.D ;
  wire \DFF_8.Q ;
  wire \DFF_80.CK ;
  wire \DFF_80.D ;
  wire \DFF_80.Q ;
  wire \DFF_81.CK ;
  wire \DFF_81.D ;
  wire \DFF_81.Q ;
  wire \DFF_82.CK ;
  wire \DFF_82.D ;
  wire \DFF_82.Q ;
  wire \DFF_83.CK ;
  wire \DFF_83.D ;
  wire \DFF_83.Q ;
  wire \DFF_84.CK ;
  wire \DFF_84.D ;
  wire \DFF_84.Q ;
  wire \DFF_85.CK ;
  wire \DFF_85.D ;
  wire \DFF_85.Q ;
  wire \DFF_86.CK ;
  wire \DFF_86.D ;
  wire \DFF_86.Q ;
  wire \DFF_87.CK ;
  wire \DFF_87.D ;
  wire \DFF_87.Q ;
  wire \DFF_88.CK ;
  wire \DFF_88.D ;
  wire \DFF_88.Q ;
  wire \DFF_89.CK ;
  wire \DFF_89.D ;
  wire \DFF_89.Q ;
  wire \DFF_9.CK ;
  wire \DFF_9.D ;
  wire \DFF_9.Q ;
  wire \DFF_90.CK ;
  wire \DFF_90.D ;
  wire \DFF_90.Q ;
  wire \DFF_91.CK ;
  wire \DFF_91.D ;
  wire \DFF_91.Q ;
  wire \DFF_92.CK ;
  wire \DFF_92.D ;
  wire \DFF_92.Q ;
  wire \DFF_93.CK ;
  wire \DFF_93.D ;
  wire \DFF_93.Q ;
  wire \DFF_94.CK ;
  wire \DFF_94.D ;
  wire \DFF_94.Q ;
  wire \DFF_95.CK ;
  wire \DFF_95.D ;
  wire \DFF_95.Q ;
  wire \DFF_96.CK ;
  wire \DFF_96.D ;
  wire \DFF_96.Q ;
  wire \DFF_97.CK ;
  wire \DFF_97.D ;
  wire \DFF_97.Q ;
  wire \DFF_98.CK ;
  wire \DFF_98.D ;
  wire \DFF_98.Q ;
  wire \DFF_99.CK ;
  wire \DFF_99.D ;
  wire \DFF_99.Q ;
  input GND;
  wire II1007;
  wire II1011;
  wire II1016;
  wire II1067;
  wire II1079;
  wire II1103;
  wire II1115;
  wire II1138;
  wire II1141;
  wire II1152;
  wire II1155;
  wire II1166;
  wire II1169;
  wire II1174;
  wire II1178;
  wire II1183;
  wire II1201;
  wire II1204;
  wire II1209;
  wire II1227;
  wire II1230;
  wire II1236;
  wire II1344;
  wire II1348;
  wire II1353;
  wire II1371;
  wire II1374;
  wire II1385;
  wire II1388;
  wire II1399;
  wire II1402;
  wire II1407;
  wire II1411;
  wire II1416;
  wire II1450;
  wire II1453;
  wire II1464;
  wire II1467;
  wire II1472;
  wire II1476;
  wire II1481;
  wire II1538;
  wire II1550;
  wire II1606;
  wire II1617;
  wire II1630;
  wire II1703;
  wire II1708;
  wire II1719;
  wire II1791;
  wire II1795;
  wire II1800;
  wire II1899;
  wire II1903;
  wire II1908;
  wire II196;
  wire II1961;
  wire II203;
  wire II2040;
  wire II2044;
  wire II2049;
  wire II210;
  wire II2153;
  wire II2157;
  wire II2162;
  wire II2213;
  wire II2225;
  wire II2228;
  wire II2232;
  wire II2235;
  wire II2238;
  wire II2242;
  wire II2251;
  wire II2254;
  wire II2257;
  wire II2260;
  wire II2263;
  wire II2268;
  wire II2271;
  wire II2275;
  wire II2316;
  wire II2319;
  wire II2344;
  wire II2349;
  wire II2372;
  wire II2376;
  wire II2380;
  wire II2385;
  wire II2389;
  wire II2394;
  wire II2403;
  wire II2414;
  wire II2417;
  wire II2420;
  wire II2425;
  wire II2428;
  wire II2433;
  wire II2813;
  wire II3143;
  wire II3168;
  wire II3315;
  wire II3318;
  wire II3339;
  wire II3342;
  wire II3394;
  wire II3461;
  wire II3509;
  wire II3587;
  wire II359;
  wire II363;
  wire II368;
  wire II406;
  wire II409;
  wire II4117;
  wire II4122;
  wire II414;
  wire II4222;
  wire II4227;
  wire II4482;
  wire II4485;
  wire II4489;
  wire II4492;
  wire II4496;
  wire II4499;
  wire II453;
  wire II4558;
  wire II456;
  wire II461;
  wire II4626;
  wire II4630;
  wire II4633;
  wire II4660;
  wire II4720;
  wire II4723;
  wire II4726;
  wire II642;
  wire II646;
  wire II651;
  wire II683;
  wire II687;
  wire II692;
  wire II726;
  wire II729;
  wire II734;
  wire II842;
  wire II846;
  wire II851;
  wire II921;
  wire II925;
  wire II930;
  input VDD;
  wire n1018gat;
  wire n1019gat;
  wire n1020gat;
  wire n1025gat;
  wire n1026gat;
  wire n1034gat;
  wire n1035gat;
  wire n1044gat;
  wire n1045gat;
  wire n1055gat;
  wire n1056gat;
  wire n1057gat;
  wire n1067gat;
  wire n1068gat;
  wire n1071gat;
  wire n1072gat;
  wire n1079gat;
  wire n1080gat;
  wire n1084gat;
  wire n1085gat;
  wire n1086gat;
  wire n1118gat;
  wire n1120gat;
  wire n1121gat;
  wire n1134gat;
  wire n1135gat;
  wire n1147gat;
  wire n1148gat;
  wire n1150gat;
  wire n1189gat;
  wire n1190gat;
  wire n1191gat;
  wire n1196gat;
  wire n1197gat;
  wire n1206gat;
  wire n1207gat;
  wire n1208gat;
  wire n1221gat;
  wire n1222gat;
  wire n1223gat;
  wire n1225gat;
  wire n1226gat;
  wire n1233gat;
  wire n1234gat;
  wire n1235gat;
  wire n1240gat;
  wire n1241gat;
  wire n1269gat;
  wire n1281gat;
  wire n1282gat;
  wire n1293gat;
  wire n1294gat;
  wire n1297gat;
  wire n1298gat;
  wire n1311gat;
  wire n1312gat;
  wire n1314gat;
  wire n1315gat;
  wire n1316gat;
  wire n1328gat;
  wire n1330gat;
  wire n1332gat;
  wire n1336gat;
  wire n1339gat;
  wire n1340gat;
  wire n1350gat;
  wire n1361gat;
  wire n1363gat;
  wire n1382gat;
  wire n1389gat;
  wire n1391gat;
  wire n1392gat;
  wire n1393gat;
  wire n1394gat;
  wire n1431gat;
  wire n1433gat;
  wire n1442gat;
  wire n1455gat;
  wire n1456gat;
  wire n1461gat;
  wire n1462gat;
  wire n147gat;
  wire n148gat;
  wire n1495gat;
  wire n1496gat;
  wire n1507gat;
  wire n1508gat;
  wire n1516gat;
  wire n1518gat;
  wire n151gat;
  wire n1524gat;
  wire n1525gat;
  wire n152gat;
  wire n155gat;
  wire n1564gat;
  wire n1565gat;
  wire n1567gat;
  wire n156gat;
  wire n1587gat;
  wire n1588gat;
  wire n1593gat;
  wire n1595gat;
  wire n1596gat;
  wire n159gat;
  wire n1603gat;
  wire n1606gat;
  wire n160gat;
  wire n1610gat;
  wire n1613gat;
  wire n1620gat;
  wire n1625gat;
  wire n1626gat;
  wire n1631gat;
  wire n1632gat;
  wire n1633gat;
  wire n1636gat;
  wire n164gat;
  wire n1658gat;
  wire n165gat;
  wire n1674gat;
  wire n1675gat;
  wire n1677gat;
  wire n1678gat;
  wire n1685gat;
  wire n1691gat;
  wire n1696gat;
  wire n1699gat;
  wire n1708gat;
  wire n1712gat;
  wire n1713gat;
  wire n1717gat;
  wire n1721gat;
  wire n172gat;
  wire n1739gat;
  wire n173gat;
  wire n1740gat;
  wire n1742gat;
  wire n1745gat;
  wire n1747gat;
  wire n1748gat;
  wire n174gat;
  wire n1762gat;
  wire n1763gat;
  wire n1767gat;
  wire n1771gat;
  wire n1773gat;
  wire n1774gat;
  wire n1775gat;
  wire n1777gat;
  wire n1781gat;
  wire n1783gat;
  wire n1785gat;
  wire n1787gat;
  wire n1793gat;
  wire n1800gat;
  wire n1806gat;
  wire n1807gat;
  wire n1816gat;
  wire n1821gat;
  wire n1825gat;
  wire n1827gat;
  wire n1828gat;
  wire n1829gat;
  wire n1834gat;
  wire n1836gat;
  wire n1845gat;
  wire n1849gat;
  wire n1850gat;
  wire n1858gat;
  wire n1869gat;
  wire n1870gat;
  wire n1871gat;
  wire n1879gat;
  wire n1880gat;
  wire n1882gat;
  wire n1884gat;
  wire n1886gat;
  wire n1891gat;
  wire n1898gat;
  wire n1899gat;
  wire n1915gat;
  wire n1918gat;
  wire n1927gat;
  wire n1945gat;
  wire n1954gat;
  wire n1955gat;
  wire n1963gat;
  wire n1974gat;
  wire n1975gat;
  wire n1988gat;
  wire n1989gat;
  wire n2009gat;
  wire n2015gat;
  wire n2017gat;
  wire n2021gat;
  wire n2023gat;
  wire n2025gat;
  wire n2027gat;
  wire n2029gat;
  wire n2031gat;
  wire n2033gat;
  wire n2035gat;
  wire n2037gat;
  wire n2039gat;
  wire n2040gat;
  wire n2042gat;
  wire n2044gat;
  wire n2046gat;
  wire n2057gat;
  wire n2060gat;
  wire n2061gat;
  wire n2084gat;
  wire n2090gat;
  wire n2091gat;
  wire n2093gat;
  wire n2095gat;
  wire n2099gat;
  wire n2101gat;
  wire n2102gat;
  wire n2108gat;
  wire n2110gat;
  wire n2117gat;
  wire n2119gat;
  wire n2121gat;
  wire n2123gat;
  wire n2124gat;
  wire n2125gat;
  wire n2127gat;
  wire n2134gat;
  wire n2135gat;
  wire n2138gat;
  wire n2139gat;
  wire n2142gat;
  wire n2143gat;
  wire n2154gat;
  wire n2155gat;
  wire n2163gat;
  wire n2168gat;
  wire n2169gat;
  wire n2174gat;
  wire n2176gat;
  wire n2178gat;
  wire n2179gat;
  wire n2181gat;
  wire n2182gat;
  wire n2189gat;
  wire n2190gat;
  wire n2192gat;
  wire n2194gat;
  wire n2196gat;
  wire n2197gat;
  wire n2198gat;
  wire n2201gat;
  wire n2202gat;
  wire n2203gat;
  wire n2205gat;
  wire n2206gat;
  wire n2207gat;
  wire n2214gat;
  wire n2217gat;
  wire n2251gat;
  wire n2252gat;
  wire n2261gat;
  wire n2262gat;
  wire n2265gat;
  wire n2266gat;
  wire n2268gat;
  wire n2269gat;
  wire n226gat;
  wire n2270gat;
  wire n227gat;
  wire n2283gat;
  wire n2284gat;
  wire n2285gat;
  wire n228gat;
  wire n2290gat;
  wire n2319gat;
  wire n2330gat;
  wire n2332gat;
  wire n2333gat;
  wire n2337gat;
  wire n2338gat;
  wire n2339gat;
  wire n2341gat;
  wire n2342gat;
  wire n2343gat;
  wire n2346gat;
  wire n2347gat;
  wire n2351gat;
  wire n2353gat;
  wire n2354gat;
  wire n2355gat;
  wire n2356gat;
  wire n2387gat;
  wire n2388gat;
  wire n2389gat;
  wire n2390gat;
  wire n2393gat;
  wire n2394gat;
  wire n2396gat;
  wire n2397gat;
  wire n2398gat;
  wire n2399gat;
  wire n2402gat;
  wire n2403gat;
  wire n2406gat;
  wire n2407gat;
  wire n2414gat;
  wire n2415gat;
  wire n2416gat;
  wire n2417gat;
  wire n2418gat;
  wire n2419gat;
  wire n2429gat;
  wire n2436gat;
  wire n2439gat;
  wire n2440gat;
  wire n2443gat;
  wire n2454gat;
  wire n2456gat;
  wire n2458gat;
  wire n2464gat;
  wire n2468gat;
  wire n2470gat;
  wire n2472gat;
  wire n2476gat;
  wire n2482gat;
  wire n2486gat;
  wire n2487gat;
  wire n2488gat;
  wire n2489gat;
  wire n2490gat;
  wire n2492gat;
  wire n2493gat;
  wire n2494gat;
  wire n2495gat;
  wire n2498gat;
  wire n2502gat;
  wire n2506gat;
  wire n2510gat;
  wire n2514gat;
  wire n2518gat;
  wire n2522gat;
  wire n2526gat;
  wire n2532gat;
  wire n2536gat;
  wire n2539gat;
  wire n2540gat;
  wire n2541gat;
  wire n2542gat;
  wire n2543gat;
  wire n2550gat;
  wire n2551gat;
  wire n2552gat;
  wire n2553gat;
  wire n2554gat;
  wire n2555gat;
  wire n2556gat;
  wire n2557gat;
  wire n2558gat;
  wire n255gat;
  wire n2560gat;
  wire n2561gat;
  wire n2562gat;
  wire n256gat;
  wire n2573gat;
  wire n2574gat;
  wire n2575gat;
  wire n2576gat;
  wire n2577gat;
  wire n2578gat;
  wire n2579gat;
  wire n2588gat;
  wire n2590gat;
  wire n2591gat;
  wire n2592gat;
  wire n2599gat;
  wire n2606gat;
  wire n2607gat;
  wire n2608gat;
  wire n2609gat;
  wire n2610gat;
  wire n2611gat;
  wire n2612gat;
  wire n2613gat;
  wire n2620gat;
  wire n2621gat;
  wire n2622gat;
  wire n2624gat;
  wire n2625gat;
  wire n2626gat;
  wire n2628gat;
  wire n2629gat;
  wire n2630gat;
  wire n2632gat;
  wire n2633gat;
  wire n2634gat;
  wire n2636gat;
  wire n2638gat;
  wire n2639gat;
  wire n263gat;
  wire n2640gat;
  wire n2643gat;
  wire n2644gat;
  wire n2646gat;
  wire n264gat;
  wire n2658gat;
  wire n265gat;
  wire n2667gat;
  wire n2668gat;
  wire n2670gat;
  wire n2671gat;
  wire n2673gat;
  wire n2674gat;
  wire n2677gat;
  wire n2678gat;
  wire n2680gat;
  wire n2681gat;
  wire n2682gat;
  wire n2684gat;
  wire n2685gat;
  wire n2686gat;
  wire n2688gat;
  wire n2689gat;
  wire n2691gat;
  wire n2692gat;
  wire n2693gat;
  wire n2696gat;
  wire n2698gat;
  wire n2699gat;
  wire n2700gat;
  wire n2702gat;
  wire n2704gat;
  wire n2705gat;
  wire n2706gat;
  wire n2708gat;
  wire n2709gat;
  wire n270gat;
  wire n2712gat;
  wire n2716gat;
  wire n2717gat;
  wire n2719gat;
  wire n271gat;
  wire n2721gat;
  wire n2722gat;
  wire n2724gat;
  wire n2725gat;
  wire n2727gat;
  wire n2728gat;
  wire n2729gat;
  wire n2730gat;
  wire n2732gat;
  wire n2733gat;
  wire n2735gat;
  wire n2736gat;
  wire n2737gat;
  wire n2738gat;
  wire n2739gat;
  wire n2740gat;
  wire n2741gat;
  wire n2742gat;
  wire n2744gat;
  wire n2745gat;
  wire n2746gat;
  wire n2747gat;
  wire n2748gat;
  wire n2749gat;
  wire n274gat;
  wire n2750gat;
  wire n2753gat;
  wire n2754gat;
  wire n2755gat;
  wire n2756gat;
  wire n2757gat;
  wire n2759gat;
  wire n275gat;
  wire n2760gat;
  wire n2761gat;
  wire n2762gat;
  wire n2763gat;
  wire n2764gat;
  wire n2765gat;
  wire n2766gat;
  wire n2767gat;
  wire n2768gat;
  wire n2776gat;
  wire n2777gat;
  wire n2779gat;
  wire n2780gat;
  wire n2782gat;
  wire n2783gat;
  wire n278gat;
  wire n2790gat;
  wire n2791gat;
  wire n2793gat;
  wire n2794gat;
  wire n2795gat;
  wire n2796gat;
  wire n2797gat;
  wire n2798gat;
  wire n2799gat;
  wire n279gat;
  wire n2800gat;
  wire n2801gat;
  wire n2802gat;
  wire n2803gat;
  wire n2804gat;
  wire n2805gat;
  wire n2806gat;
  wire n2807gat;
  wire n2808gat;
  wire n2809gat;
  wire n2810gat;
  wire n2811gat;
  wire n2812gat;
  wire n2813gat;
  wire n2814gat;
  wire n2815gat;
  wire n2816gat;
  wire n2817gat;
  wire n2818gat;
  wire n2819gat;
  wire n2820gat;
  wire n2821gat;
  wire n2822gat;
  wire n2823gat;
  wire n2824gat;
  wire n2825gat;
  wire n2826gat;
  wire n2828gat;
  wire n2829gat;
  wire n282gat;
  wire n2831gat;
  wire n2832gat;
  wire n2837gat;
  wire n2839gat;
  wire n283gat;
  wire n2841gat;
  wire n2843gat;
  wire n2845gat;
  wire n2847gat;
  wire n2850gat;
  wire n2851gat;
  wire n2853gat;
  wire n2855gat;
  wire n2856gat;
  wire n2858gat;
  wire n2860gat;
  wire n2861gat;
  wire n2863gat;
  wire n2864gat;
  wire n2868gat;
  wire n2869gat;
  wire n2886gat;
  wire n2887gat;
  wire n2888gat;
  wire n2890gat;
  wire n2891gat;
  wire n2892gat;
  wire n2894gat;
  wire n2895gat;
  wire n2896gat;
  wire n2897gat;
  wire n2898gat;
  wire n2899gat;
  wire n2900gat;
  wire n2901gat;
  wire n2903gat;
  wire n2904gat;
  wire n2905gat;
  wire n2907gat;
  wire n2908gat;
  wire n2909gat;
  wire n2910gat;
  wire n2911gat;
  wire n2912gat;
  wire n2913gat;
  wire n2914gat;
  wire n2915gat;
  wire n2916gat;
  wire n2917gat;
  wire n2918gat;
  wire n2919gat;
  wire n2920gat;
  wire n2921gat;
  wire n2922gat;
  wire n2923gat;
  wire n2924gat;
  wire n2925gat;
  wire n2926gat;
  wire n2927gat;
  wire n2928gat;
  wire n2929gat;
  wire n2935gat;
  wire n2936gat;
  wire n2937gat;
  wire n2938gat;
  wire n2941gat;
  wire n2950gat;
  wire n2951gat;
  wire n2952gat;
  wire n2955gat;
  wire n2956gat;
  wire n2971gat;
  wire n2980gat;
  wire n2983gat;
  wire n2989gat;
  wire n3010gat;
  wire n3016gat;
  wire n3020gat;
  wire n3021gat;
  wire n3022gat;
  wire n3023gat;
  wire n3024gat;
  wire n3025gat;
  wire n3026gat;
  wire n3027gat;
  wire n3028gat;
  wire n3029gat;
  wire n3030gat;
  wire n3031gat;
  wire n3032gat;
  wire n3034gat;
  wire n3035gat;
  wire n3036gat;
  wire n3037gat;
  wire n3039gat;
  wire n3040gat;
  wire n3041gat;
  wire n3042gat;
  wire n3043gat;
  wire n3044gat;
  wire n3046gat;
  wire n3047gat;
  wire n3048gat;
  wire n3049gat;
  wire n3050gat;
  wire n3051gat;
  wire n3052gat;
  wire n3053gat;
  wire n3054gat;
  wire n3055gat;
  wire n3056gat;
  wire n3057gat;
  wire n3058gat;
  wire n3059gat;
  wire n3060gat;
  wire n3061gat;
  wire n3062gat;
  wire n3063gat;
  wire n3064gat;
  input n3065gat;
  input n3066gat;
  input n3067gat;
  input n3068gat;
  input n3069gat;
  input n3070gat;
  input n3071gat;
  input n3072gat;
  input n3073gat;
  input n3074gat;
  input n3075gat;
  input n3076gat;
  input n3077gat;
  input n3078gat;
  input n3079gat;
  input n3080gat;
  input n3081gat;
  input n3082gat;
  input n3083gat;
  input n3084gat;
  input n3085gat;
  input n3086gat;
  input n3087gat;
  input n3088gat;
  input n3089gat;
  input n3090gat;
  input n3091gat;
  input n3092gat;
  input n3093gat;
  input n3094gat;
  input n3095gat;
  input n3097gat;
  input n3098gat;
  input n3099gat;
  input n3100gat;
  output n3104gat;
  output n3105gat;
  output n3106gat;
  output n3107gat;
  output n3108gat;
  output n3109gat;
  output n3110gat;
  output n3111gat;
  output n3112gat;
  output n3113gat;
  output n3114gat;
  output n3115gat;
  output n3116gat;
  output n3117gat;
  output n3118gat;
  output n3119gat;
  output n3120gat;
  output n3121gat;
  output n3122gat;
  output n3123gat;
  output n3124gat;
  output n3125gat;
  output n3126gat;
  output n3127gat;
  output n3128gat;
  output n3129gat;
  output n3130gat;
  output n3131gat;
  output n3132gat;
  output n3133gat;
  output n3134gat;
  output n3135gat;
  output n3136gat;
  output n3137gat;
  output n3138gat;
  output n3139gat;
  wire n313gat;
  output n3140gat;
  output n3141gat;
  output n3142gat;
  output n3143gat;
  output n3144gat;
  output n3145gat;
  output n3146gat;
  output n3147gat;
  output n3148gat;
  output n3149gat;
  wire n314gat;
  output n3150gat;
  output n3151gat;
  output n3152gat;
  wire n317gat;
  wire n318gat;
  wire n321gat;
  wire n322gat;
  wire n326gat;
  wire n327gat;
  wire n330gat;
  wire n331gat;
  wire n336gat;
  wire n337gat;
  wire n340gat;
  wire n341gat;
  wire n348gat;
  wire n349gat;
  wire n350gat;
  wire n365gat;
  wire n366gat;
  wire n383gat;
  wire n384gat;
  wire n387gat;
  wire n388gat;
  wire n393gat;
  wire n394gat;
  wire n397gat;
  wire n398gat;
  wire n401gat;
  wire n402gat;
  wire n43gat;
  wire n462gat;
  wire n463gat;
  wire n469gat;
  wire n470gat;
  wire n480gat;
  wire n481gat;
  wire n482gat;
  wire n490gat;
  wire n491gat;
  wire n498gat;
  wire n499gat;
  wire n500gat;
  wire n503gat;
  wire n504gat;
  wire n552gat;
  wire n553gat;
  wire n55gat;
  wire n560gat;
  wire n561gat;
  wire n566gat;
  wire n567gat;
  wire n579gat;
  wire n580gat;
  wire n583gat;
  wire n584gat;
  wire n591gat;
  wire n592gat;
  wire n593gat;
  wire n594gat;
  wire n595gat;
  wire n596gat;
  wire n612gat;
  wire n613gat;
  wire n614gat;
  wire n617gat;
  wire n618gat;
  wire n621gat;
  wire n622gat;
  wire n625gat;
  wire n626gat;
  wire n658gat;
  wire n659gat;
  wire n666gat;
  wire n667gat;
  wire n672gat;
  wire n673gat;
  wire n679gat;
  wire n680gat;
  wire n682gat;
  wire n683gat;
  wire n684gat;
  wire n691gat;
  wire n692gat;
  wire n693gat;
  wire n694gat;
  wire n695gat;
  wire n697gat;
  wire n698gat;
  wire n699gat;
  wire n702gat;
  wire n703gat;
  wire n705gat;
  wire n706gat;
  wire n707gat;
  wire n714gat;
  wire n715gat;
  wire n716gat;
  wire n717gat;
  wire n718gat;
  wire n719gat;
  wire n721gat;
  wire n722gat;
  wire n725gat;
  wire n726gat;
  wire n733gat;
  wire n734gat;
  wire n735gat;
  wire n736gat;
  wire n748gat;
  wire n776gat;
  wire n777gat;
  wire n784gat;
  wire n785gat;
  wire n786gat;
  wire n808gat;
  wire n809gat;
  wire n810gat;
  wire n815gat;
  wire n816gat;
  wire n818gat;
  wire n819gat;
  wire n820gat;
  wire n822gat;
  wire n823gat;
  wire n824gat;
  wire n827gat;
  wire n828gat;
  wire n829gat;
  wire n830gat;
  wire n832gat;
  wire n833gat;
  wire n834gat;
  wire n836gat;
  wire n837gat;
  wire n838gat;
  wire n841gat;
  wire n842gat;
  wire n845gat;
  wire n846gat;
  wire n850gat;
  wire n860gat;
  wire n861gat;
  wire n864gat;
  wire n865gat;
  wire n873gat;
  wire n875gat;
  wire n881gat;
  wire n882gat;
  wire n883gat;
  wire n911gat;
  wire n912gat;
  wire n913gat;
  wire n918gat;
  wire n919gat;
  wire n922gat;
  wire n923gat;
  wire n924gat;
  wire n927gat;
  wire n930gat;
  wire n931gat;
  wire n933gat;
  wire n949gat;
  wire n950gat;
  wire n951gat;
  wire n956gat;
  wire n957gat;
  wire n983gat;
  wire n985gat;
  al_inv _0553_ (
    .a(\DFF_16.Q ),
    .y(\DFF_17.D )
  );
  al_inv _0554_ (
    .a(\DFF_20.Q ),
    .y(\DFF_21.D )
  );
  al_inv _0555_ (
    .a(\DFF_43.Q ),
    .y(\DFF_157.D )
  );
  al_inv _0556_ (
    .a(\DFF_44.Q ),
    .y(\DFF_163.D )
  );
  al_inv _0557_ (
    .a(\DFF_42.Q ),
    .y(\DFF_165.D )
  );
  al_inv _0558_ (
    .a(\DFF_45.Q ),
    .y(\DFF_164.D )
  );
  al_inv _0559_ (
    .a(\DFF_46.Q ),
    .y(\DFF_156.D )
  );
  al_inv _0560_ (
    .a(\DFF_52.Q ),
    .y(\DFF_160.D )
  );
  al_inv _0561_ (
    .a(\DFF_53.Q ),
    .y(\DFF_159.D )
  );
  al_inv _0562_ (
    .a(\DFF_51.Q ),
    .y(\DFF_158.D )
  );
  al_inv _0563_ (
    .a(\DFF_55.Q ),
    .y(\DFF_161.D )
  );
  al_inv _0564_ (
    .a(\DFF_56.Q ),
    .y(\DFF_162.D )
  );
  al_inv _0565_ (
    .a(\DFF_93.Q ),
    .y(\DFF_155.D )
  );
  al_inv _0566_ (
    .a(\DFF_61.Q ),
    .y(\DFF_112.D )
  );
  al_inv _0567_ (
    .a(\DFF_59.Q ),
    .y(\DFF_111.D )
  );
  al_inv _0568_ (
    .a(\DFF_58.Q ),
    .y(\DFF_110.D )
  );
  al_inv _0569_ (
    .a(\DFF_95.Q ),
    .y(\DFF_148.D )
  );
  al_inv _0570_ (
    .a(\DFF_63.Q ),
    .y(\DFF_108.D )
  );
  al_inv _0571_ (
    .a(\DFF_64.Q ),
    .y(\DFF_107.D )
  );
  al_inv _0572_ (
    .a(\DFF_65.Q ),
    .y(\DFF_106.D )
  );
  al_inv _0573_ (
    .a(\DFF_100.Q ),
    .y(\DFF_154.D )
  );
  al_inv _0574_ (
    .a(\DFF_67.Q ),
    .y(\DFF_105.D )
  );
  al_inv _0575_ (
    .a(\DFF_66.Q ),
    .y(\DFF_109.D )
  );
  al_inv _0576_ (
    .a(\DFF_60.Q ),
    .y(\DFF_114.D )
  );
  al_inv _0577_ (
    .a(\DFF_62.Q ),
    .y(\DFF_113.D )
  );
  al_inv _0578_ (
    .a(\DFF_120.Q ),
    .y(\DFF_121.D )
  );
  al_or3 _0579_ (
    .a(\DFF_108.Q ),
    .b(\DFF_106.Q ),
    .c(\DFF_107.Q ),
    .y(_0096_)
  );
  al_and3fft _0580_ (
    .a(\DFF_105.Q ),
    .b(_0096_),
    .c(\DFF_109.Q ),
    .y(\DFF_172.D )
  );
  al_and3ftt _0581_ (
    .a(\DFF_106.Q ),
    .b(\DFF_109.Q ),
    .c(\DFF_107.Q ),
    .y(_0097_)
  );
  al_and3ftt _0582_ (
    .a(\DFF_108.Q ),
    .b(\DFF_105.Q ),
    .c(_0097_),
    .y(\DFF_171.D )
  );
  al_inv _0583_ (
    .a(\DFF_127.Q ),
    .y(\DFF_128.D )
  );
  al_inv _0584_ (
    .a(\DFF_129.Q ),
    .y(\DFF_130.D )
  );
  al_oa21 _0585_ (
    .a(\DFF_69.Q ),
    .b(\DFF_70.Q ),
    .c(\DFF_68.Q ),
    .y(_0098_)
  );
  al_inv _0586_ (
    .a(_0098_),
    .y(\DFF_71.D )
  );
  al_inv _0587_ (
    .a(\DFF_117.Q ),
    .y(\DFF_118.D )
  );
  al_and3 _0588_ (
    .a(\DFF_108.Q ),
    .b(\DFF_105.Q ),
    .c(_0097_),
    .y(\DFF_135.D )
  );
  al_inv _0589_ (
    .a(\DFF_139.Q ),
    .y(\DFF_140.D )
  );
  al_inv _0590_ (
    .a(\DFF_140.Q ),
    .y(\DFF_141.D )
  );
  al_inv _0591_ (
    .a(\DFF_131.Q ),
    .y(\DFF_133.D )
  );
  al_inv _0592_ (
    .a(\DFF_128.Q ),
    .y(\DFF_129.D )
  );
  al_inv _0593_ (
    .a(\DFF_144.Q ),
    .y(\DFF_145.D )
  );
  al_inv _0594_ (
    .a(\DFF_145.Q ),
    .y(\DFF_149.D )
  );
  al_inv _0595_ (
    .a(\DFF_146.Q ),
    .y(\DFF_147.D )
  );
  al_and2 _0596_ (
    .a(\DFF_9.Q ),
    .b(\DFF_92.Q ),
    .y(_0099_)
  );
  al_and3 _0597_ (
    .a(\DFF_94.Q ),
    .b(\DFF_99.Q ),
    .c(\DFF_101.Q ),
    .y(_0100_)
  );
  al_ao21 _0598_ (
    .a(_0100_),
    .b(_0099_),
    .c(n3100gat),
    .y(_0101_)
  );
  al_ao21ttf _0599_ (
    .a(\DFF_69.Q ),
    .b(\DFF_116.Q ),
    .c(\DFF_147.Q ),
    .y(_0102_)
  );
  al_and2 _0600_ (
    .a(\DFF_139.Q ),
    .b(\DFF_145.Q ),
    .y(_0103_)
  );
  al_and3 _0601_ (
    .a(_0102_),
    .b(_0103_),
    .c(_0101_),
    .y(\DFF_96.D )
  );
  al_and3fft _0602_ (
    .a(\DFF_114.Q ),
    .b(\DFF_113.Q ),
    .c(\DFF_110.Q ),
    .y(_0104_)
  );
  al_and2ft _0603_ (
    .a(\DFF_111.Q ),
    .b(\DFF_112.Q ),
    .y(_0105_)
  );
  al_and2ft _0604_ (
    .a(\DFF_112.Q ),
    .b(\DFF_111.Q ),
    .y(_0106_)
  );
  al_mux2l _0605_ (
    .a(_0106_),
    .b(_0105_),
    .s(_0098_),
    .y(_0107_)
  );
  al_and2 _0606_ (
    .a(_0104_),
    .b(_0107_),
    .y(_0108_)
  );
  al_and2 _0607_ (
    .a(\DFF_112.Q ),
    .b(\DFF_111.Q ),
    .y(_0109_)
  );
  al_and3fft _0608_ (
    .a(_0109_),
    .b(_0108_),
    .c(\DFF_96.D ),
    .y(\DFF_59.D )
  );
  al_inv _0609_ (
    .a(_0104_),
    .y(_0110_)
  );
  al_aoi21ftf _0610_ (
    .a(_0110_),
    .b(_0107_),
    .c(\DFF_96.D ),
    .y(\DFF_61.D )
  );
  al_or3 _0611_ (
    .a(\DFF_110.Q ),
    .b(\DFF_112.Q ),
    .c(\DFF_111.Q ),
    .y(_0111_)
  );
  al_oai21ttf _0612_ (
    .a(\DFF_114.Q ),
    .b(_0111_),
    .c(\DFF_113.Q ),
    .y(_0112_)
  );
  al_and3fft _0613_ (
    .a(\DFF_114.Q ),
    .b(_0111_),
    .c(\DFF_113.Q ),
    .y(_0113_)
  );
  al_aoi21ftf _0614_ (
    .a(_0113_),
    .b(_0112_),
    .c(\DFF_61.D ),
    .y(\DFF_62.D )
  );
  al_nor2 _0615_ (
    .a(\DFF_112.Q ),
    .b(\DFF_111.Q ),
    .y(_0114_)
  );
  al_nand3fft _0616_ (
    .a(\DFF_114.Q ),
    .b(\DFF_110.Q ),
    .c(_0114_),
    .y(_0115_)
  );
  al_and2 _0617_ (
    .a(\DFF_114.Q ),
    .b(_0111_),
    .y(_0116_)
  );
  al_and3ftt _0618_ (
    .a(_0116_),
    .b(_0115_),
    .c(\DFF_61.D ),
    .y(\DFF_60.D )
  );
  al_inv _0619_ (
    .a(\DFF_149.Q ),
    .y(\DFF_150.D )
  );
  al_inv _0620_ (
    .a(\DFF_150.Q ),
    .y(\DFF_151.D )
  );
  al_inv _0621_ (
    .a(\DFF_151.Q ),
    .y(\DFF_152.D )
  );
  al_inv _0622_ (
    .a(\DFF_152.Q ),
    .y(\DFF_153.D )
  );
  al_and3ftt _0623_ (
    .a(\DFF_151.Q ),
    .b(\DFF_153.Q ),
    .c(n3100gat),
    .y(\DFF_69.D )
  );
  al_inv _0624_ (
    .a(\DFF_133.Q ),
    .y(\DFF_166.D )
  );
  al_inv _0625_ (
    .a(\DFF_166.Q ),
    .y(\DFF_167.D )
  );
  al_nand2ft _0626_ (
    .a(\DFF_59.Q ),
    .b(\DFF_61.Q ),
    .y(_0117_)
  );
  al_and2ft _0627_ (
    .a(\DFF_61.Q ),
    .b(\DFF_59.Q ),
    .y(_0118_)
  );
  al_oai21ftf _0628_ (
    .a(_0117_),
    .b(_0118_),
    .c(\DFF_93.Q ),
    .y(_0119_)
  );
  al_nor3fft _0629_ (
    .a(\DFF_93.Q ),
    .b(_0117_),
    .c(_0118_),
    .y(_0120_)
  );
  al_nand2ft _0630_ (
    .a(\DFF_62.Q ),
    .b(\DFF_60.Q ),
    .y(_0121_)
  );
  al_nand2ft _0631_ (
    .a(\DFF_60.Q ),
    .b(\DFF_62.Q ),
    .y(_0122_)
  );
  al_and3ftt _0632_ (
    .a(\DFF_58.Q ),
    .b(_0121_),
    .c(_0122_),
    .y(_0123_)
  );
  al_ao21 _0633_ (
    .a(_0121_),
    .b(_0122_),
    .c(\DFF_110.D ),
    .y(_0124_)
  );
  al_nand2ft _0634_ (
    .a(_0123_),
    .b(_0124_),
    .y(_0125_)
  );
  al_and3ftt _0635_ (
    .a(_0120_),
    .b(_0119_),
    .c(_0125_),
    .y(_0126_)
  );
  al_ao21ftt _0636_ (
    .a(_0120_),
    .b(_0119_),
    .c(_0125_),
    .y(_0127_)
  );
  al_nand2ft _0637_ (
    .a(_0126_),
    .b(_0127_),
    .y(\DFF_94.D )
  );
  al_nor2 _0638_ (
    .a(\DFF_67.Q ),
    .b(\DFF_66.Q ),
    .y(_0128_)
  );
  al_nand2 _0639_ (
    .a(\DFF_67.Q ),
    .b(\DFF_66.Q ),
    .y(_0129_)
  );
  al_and2ft _0640_ (
    .a(_0128_),
    .b(_0129_),
    .y(_0130_)
  );
  al_and2ft _0641_ (
    .a(\DFF_64.Q ),
    .b(\DFF_63.Q ),
    .y(_0131_)
  );
  al_nand2ft _0642_ (
    .a(\DFF_63.Q ),
    .b(\DFF_64.Q ),
    .y(_0132_)
  );
  al_nor2 _0643_ (
    .a(\DFF_65.Q ),
    .b(\DFF_100.Q ),
    .y(_0133_)
  );
  al_nand2 _0644_ (
    .a(\DFF_65.Q ),
    .b(\DFF_100.Q ),
    .y(_0134_)
  );
  al_nand2ft _0645_ (
    .a(_0133_),
    .b(_0134_),
    .y(_0135_)
  );
  al_nand3ftt _0646_ (
    .a(_0131_),
    .b(_0132_),
    .c(_0135_),
    .y(_0136_)
  );
  al_ao21ftt _0647_ (
    .a(_0131_),
    .b(_0132_),
    .c(_0135_),
    .y(_0137_)
  );
  al_ao21 _0648_ (
    .a(_0136_),
    .b(_0137_),
    .c(_0130_),
    .y(_0138_)
  );
  al_and3 _0649_ (
    .a(_0130_),
    .b(_0136_),
    .c(_0137_),
    .y(_0139_)
  );
  al_nand2ft _0650_ (
    .a(_0139_),
    .b(_0138_),
    .y(\DFF_101.D )
  );
  al_and3 _0651_ (
    .a(\DFF_109.Q ),
    .b(\DFF_105.Q ),
    .c(\DFF_106.Q ),
    .y(_0140_)
  );
  al_and3ftt _0652_ (
    .a(\DFF_107.Q ),
    .b(\DFF_108.Q ),
    .c(_0140_),
    .y(\DFF_175.D )
  );
  al_and2ft _0653_ (
    .a(\DFF_97.Q ),
    .b(\DFF_96.Q ),
    .y(_0141_)
  );
  al_nand2ft _0654_ (
    .a(\DFF_96.Q ),
    .b(\DFF_97.Q ),
    .y(_0142_)
  );
  al_nand2 _0655_ (
    .a(\DFF_95.Q ),
    .b(\DFF_98.Q ),
    .y(_0143_)
  );
  al_nor2 _0656_ (
    .a(\DFF_95.Q ),
    .b(\DFF_98.Q ),
    .y(_0144_)
  );
  al_nand2ft _0657_ (
    .a(_0144_),
    .b(_0143_),
    .y(_0145_)
  );
  al_and3ftt _0658_ (
    .a(_0141_),
    .b(_0142_),
    .c(_0145_),
    .y(_0146_)
  );
  al_ao21ftt _0659_ (
    .a(_0141_),
    .b(_0142_),
    .c(_0145_),
    .y(_0147_)
  );
  al_nand2ft _0660_ (
    .a(_0146_),
    .b(_0147_),
    .y(\DFF_99.D )
  );
  al_nand2 _0661_ (
    .a(\DFF_78.Q ),
    .b(\DFF_79.Q ),
    .y(_0148_)
  );
  al_or2 _0662_ (
    .a(\DFF_78.Q ),
    .b(\DFF_79.Q ),
    .y(_0149_)
  );
  al_ao21ttf _0663_ (
    .a(_0149_),
    .b(_0148_),
    .c(\DFF_77.Q ),
    .y(_0150_)
  );
  al_and3ftt _0664_ (
    .a(\DFF_77.Q ),
    .b(_0149_),
    .c(_0148_),
    .y(_0151_)
  );
  al_and2ft _0665_ (
    .a(_0151_),
    .b(_0150_),
    .y(_0152_)
  );
  al_nand2ft _0666_ (
    .a(\DFF_75.Q ),
    .b(\DFF_76.Q ),
    .y(_0153_)
  );
  al_nand2ft _0667_ (
    .a(\DFF_76.Q ),
    .b(\DFF_75.Q ),
    .y(_0154_)
  );
  al_nand3 _0668_ (
    .a(\DFF_73.Q ),
    .b(_0153_),
    .c(_0154_),
    .y(_0155_)
  );
  al_ao21 _0669_ (
    .a(_0153_),
    .b(_0154_),
    .c(\DFF_73.Q ),
    .y(_0156_)
  );
  al_and2ft _0670_ (
    .a(\DFF_72.Q ),
    .b(\DFF_74.Q ),
    .y(_0157_)
  );
  al_nand2ft _0671_ (
    .a(\DFF_74.Q ),
    .b(\DFF_72.Q ),
    .y(_0158_)
  );
  al_nand2ft _0672_ (
    .a(_0157_),
    .b(_0158_),
    .y(_0159_)
  );
  al_ao21 _0673_ (
    .a(_0155_),
    .b(_0156_),
    .c(_0159_),
    .y(_0160_)
  );
  al_nand3 _0674_ (
    .a(_0155_),
    .b(_0156_),
    .c(_0159_),
    .y(_0161_)
  );
  al_aoi21 _0675_ (
    .a(_0160_),
    .b(_0161_),
    .c(_0152_),
    .y(_0162_)
  );
  al_nand3 _0676_ (
    .a(_0160_),
    .b(_0152_),
    .c(_0161_),
    .y(_0163_)
  );
  al_oai21ftt _0677_ (
    .a(_0163_),
    .b(_0162_),
    .c(\DFF_80.Q ),
    .y(_0164_)
  );
  al_and3fft _0678_ (
    .a(\DFF_80.Q ),
    .b(_0162_),
    .c(_0163_),
    .y(_0165_)
  );
  al_nand2ft _0679_ (
    .a(_0165_),
    .b(_0164_),
    .y(\DFF_81.D )
  );
  al_nand2ft _0680_ (
    .a(\DFF_89.Q ),
    .b(\DFF_88.Q ),
    .y(_0166_)
  );
  al_nand2ft _0681_ (
    .a(\DFF_88.Q ),
    .b(\DFF_89.Q ),
    .y(_0167_)
  );
  al_and3 _0682_ (
    .a(\DFF_90.Q ),
    .b(_0166_),
    .c(_0167_),
    .y(_0168_)
  );
  al_ao21 _0683_ (
    .a(_0166_),
    .b(_0167_),
    .c(\DFF_90.Q ),
    .y(_0169_)
  );
  al_nand2ft _0684_ (
    .a(_0168_),
    .b(_0169_),
    .y(_0170_)
  );
  al_nand2ft _0685_ (
    .a(\DFF_85.Q ),
    .b(\DFF_84.Q ),
    .y(_0171_)
  );
  al_and2ft _0686_ (
    .a(\DFF_84.Q ),
    .b(\DFF_85.Q ),
    .y(_0172_)
  );
  al_nor3fft _0687_ (
    .a(\DFF_83.Q ),
    .b(_0171_),
    .c(_0172_),
    .y(_0173_)
  );
  al_nand2 _0688_ (
    .a(\DFF_84.Q ),
    .b(\DFF_85.Q ),
    .y(_0174_)
  );
  al_or2 _0689_ (
    .a(\DFF_84.Q ),
    .b(\DFF_85.Q ),
    .y(_0175_)
  );
  al_nand3ftt _0690_ (
    .a(\DFF_83.Q ),
    .b(_0175_),
    .c(_0174_),
    .y(_0176_)
  );
  al_nand2ft _0691_ (
    .a(\DFF_87.Q ),
    .b(\DFF_86.Q ),
    .y(_0177_)
  );
  al_and2ft _0692_ (
    .a(\DFF_86.Q ),
    .b(\DFF_87.Q ),
    .y(_0178_)
  );
  al_and2ft _0693_ (
    .a(_0178_),
    .b(_0177_),
    .y(_0179_)
  );
  al_nand3ftt _0694_ (
    .a(_0173_),
    .b(_0176_),
    .c(_0179_),
    .y(_0180_)
  );
  al_oai21ftf _0695_ (
    .a(_0176_),
    .b(_0173_),
    .c(_0179_),
    .y(_0181_)
  );
  al_nand3ftt _0696_ (
    .a(_0170_),
    .b(_0180_),
    .c(_0181_),
    .y(_0182_)
  );
  al_ao21ttf _0697_ (
    .a(_0181_),
    .b(_0180_),
    .c(_0170_),
    .y(_0183_)
  );
  al_and3 _0698_ (
    .a(\DFF_82.Q ),
    .b(_0183_),
    .c(_0182_),
    .y(_0184_)
  );
  al_ao21 _0699_ (
    .a(_0181_),
    .b(_0180_),
    .c(_0170_),
    .y(_0185_)
  );
  al_nand3 _0700_ (
    .a(_0181_),
    .b(_0170_),
    .c(_0180_),
    .y(_0186_)
  );
  al_nand3ftt _0701_ (
    .a(\DFF_82.Q ),
    .b(_0185_),
    .c(_0186_),
    .y(_0187_)
  );
  al_nand2ft _0702_ (
    .a(_0184_),
    .b(_0187_),
    .y(\DFF_91.D )
  );
  al_nand2ft _0703_ (
    .a(\DFF_42.Q ),
    .b(\DFF_46.Q ),
    .y(_0188_)
  );
  al_and2ft _0704_ (
    .a(\DFF_46.Q ),
    .b(\DFF_42.Q ),
    .y(_0189_)
  );
  al_oai21ftf _0705_ (
    .a(_0188_),
    .b(_0189_),
    .c(\DFF_163.D ),
    .y(_0190_)
  );
  al_and3fft _0706_ (
    .a(\DFF_44.Q ),
    .b(_0189_),
    .c(_0188_),
    .y(_0191_)
  );
  al_nand2ft _0707_ (
    .a(_0191_),
    .b(_0190_),
    .y(_0192_)
  );
  al_nand2ft _0708_ (
    .a(\DFF_38.Q ),
    .b(\DFF_39.Q ),
    .y(_0193_)
  );
  al_nand2ft _0709_ (
    .a(\DFF_39.Q ),
    .b(\DFF_38.Q ),
    .y(_0194_)
  );
  al_nand2ft _0710_ (
    .a(\DFF_41.Q ),
    .b(\DFF_40.Q ),
    .y(_0195_)
  );
  al_and2ft _0711_ (
    .a(\DFF_40.Q ),
    .b(\DFF_41.Q ),
    .y(_0196_)
  );
  al_nand2ft _0712_ (
    .a(_0196_),
    .b(_0195_),
    .y(_0197_)
  );
  al_or3fft _0713_ (
    .a(_0193_),
    .b(_0194_),
    .c(_0197_),
    .y(_0198_)
  );
  al_ao21ttf _0714_ (
    .a(_0193_),
    .b(_0194_),
    .c(_0197_),
    .y(_0199_)
  );
  al_ao21 _0715_ (
    .a(_0199_),
    .b(_0198_),
    .c(_0192_),
    .y(_0200_)
  );
  al_nand3 _0716_ (
    .a(_0199_),
    .b(_0192_),
    .c(_0198_),
    .y(_0201_)
  );
  al_and2ft _0717_ (
    .a(\DFF_43.Q ),
    .b(\DFF_45.Q ),
    .y(_0202_)
  );
  al_nand2ft _0718_ (
    .a(\DFF_45.Q ),
    .b(\DFF_43.Q ),
    .y(_0203_)
  );
  al_nand2ft _0719_ (
    .a(_0202_),
    .b(_0203_),
    .y(_0204_)
  );
  al_and3 _0720_ (
    .a(_0204_),
    .b(_0200_),
    .c(_0201_),
    .y(_0205_)
  );
  al_ao21 _0721_ (
    .a(_0200_),
    .b(_0201_),
    .c(_0204_),
    .y(_0206_)
  );
  al_nand2ft _0722_ (
    .a(_0205_),
    .b(_0206_),
    .y(\DFF_47.D )
  );
  al_inv _0723_ (
    .a(\DFF_54.Q ),
    .y(_0207_)
  );
  al_nand2 _0724_ (
    .a(\DFF_53.Q ),
    .b(\DFF_56.Q ),
    .y(_0208_)
  );
  al_or2 _0725_ (
    .a(\DFF_53.Q ),
    .b(\DFF_56.Q ),
    .y(_0209_)
  );
  al_aoi21 _0726_ (
    .a(_0209_),
    .b(_0208_),
    .c(_0207_),
    .y(_0210_)
  );
  al_nand3ftt _0727_ (
    .a(\DFF_54.Q ),
    .b(_0209_),
    .c(_0208_),
    .y(_0211_)
  );
  al_nor2ft _0728_ (
    .a(_0211_),
    .b(_0210_),
    .y(_0212_)
  );
  al_nor2 _0729_ (
    .a(\DFF_49.Q ),
    .b(\DFF_50.Q ),
    .y(_0213_)
  );
  al_nand2 _0730_ (
    .a(\DFF_49.Q ),
    .b(\DFF_50.Q ),
    .y(_0214_)
  );
  al_and2ft _0731_ (
    .a(_0213_),
    .b(_0214_),
    .y(_0215_)
  );
  al_nor2 _0732_ (
    .a(\DFF_52.Q ),
    .b(\DFF_51.Q ),
    .y(_0216_)
  );
  al_and2 _0733_ (
    .a(\DFF_52.Q ),
    .b(\DFF_51.Q ),
    .y(_0217_)
  );
  al_nand2ft _0734_ (
    .a(\DFF_48.Q ),
    .b(\DFF_55.Q ),
    .y(_0218_)
  );
  al_and2ft _0735_ (
    .a(\DFF_55.Q ),
    .b(\DFF_48.Q ),
    .y(_0219_)
  );
  al_and2ft _0736_ (
    .a(_0219_),
    .b(_0218_),
    .y(_0220_)
  );
  al_nand3fft _0737_ (
    .a(_0216_),
    .b(_0217_),
    .c(_0220_),
    .y(_0221_)
  );
  al_oai21ttf _0738_ (
    .a(_0216_),
    .b(_0217_),
    .c(_0220_),
    .y(_0222_)
  );
  al_nand3 _0739_ (
    .a(_0215_),
    .b(_0221_),
    .c(_0222_),
    .y(_0223_)
  );
  al_ao21 _0740_ (
    .a(_0221_),
    .b(_0222_),
    .c(_0215_),
    .y(_0224_)
  );
  al_aoi21 _0741_ (
    .a(_0223_),
    .b(_0224_),
    .c(_0212_),
    .y(_0225_)
  );
  al_and3 _0742_ (
    .a(_0212_),
    .b(_0223_),
    .c(_0224_),
    .y(_0226_)
  );
  al_nor2 _0743_ (
    .a(_0226_),
    .b(_0225_),
    .y(\DFF_57.D )
  );
  al_nand2 _0744_ (
    .a(\DFF_30.Q ),
    .b(\DFF_28.Q ),
    .y(_0227_)
  );
  al_or2 _0745_ (
    .a(\DFF_30.Q ),
    .b(\DFF_28.Q ),
    .y(_0228_)
  );
  al_aoi21ttf _0746_ (
    .a(_0228_),
    .b(_0227_),
    .c(\DFF_36.Q ),
    .y(_0229_)
  );
  al_nand3ftt _0747_ (
    .a(\DFF_36.Q ),
    .b(_0228_),
    .c(_0227_),
    .y(_0230_)
  );
  al_nor2ft _0748_ (
    .a(_0230_),
    .b(_0229_),
    .y(_0231_)
  );
  al_nor2 _0749_ (
    .a(\DFF_29.Q ),
    .b(\DFF_32.Q ),
    .y(_0232_)
  );
  al_nand2 _0750_ (
    .a(\DFF_29.Q ),
    .b(\DFF_32.Q ),
    .y(_0233_)
  );
  al_and2ft _0751_ (
    .a(_0232_),
    .b(_0233_),
    .y(_0234_)
  );
  al_nor2 _0752_ (
    .a(\DFF_35.Q ),
    .b(\DFF_34.Q ),
    .y(_0235_)
  );
  al_and2 _0753_ (
    .a(\DFF_35.Q ),
    .b(\DFF_34.Q ),
    .y(_0236_)
  );
  al_nand2ft _0754_ (
    .a(\DFF_31.Q ),
    .b(\DFF_33.Q ),
    .y(_0237_)
  );
  al_and2ft _0755_ (
    .a(\DFF_33.Q ),
    .b(\DFF_31.Q ),
    .y(_0238_)
  );
  al_and2ft _0756_ (
    .a(_0238_),
    .b(_0237_),
    .y(_0239_)
  );
  al_nand3fft _0757_ (
    .a(_0235_),
    .b(_0236_),
    .c(_0239_),
    .y(_0240_)
  );
  al_oai21ttf _0758_ (
    .a(_0235_),
    .b(_0236_),
    .c(_0239_),
    .y(_0241_)
  );
  al_nand3 _0759_ (
    .a(_0234_),
    .b(_0240_),
    .c(_0241_),
    .y(_0242_)
  );
  al_ao21 _0760_ (
    .a(_0240_),
    .b(_0241_),
    .c(_0234_),
    .y(_0243_)
  );
  al_aoi21 _0761_ (
    .a(_0242_),
    .b(_0243_),
    .c(_0231_),
    .y(_0244_)
  );
  al_and3 _0762_ (
    .a(_0231_),
    .b(_0242_),
    .c(_0243_),
    .y(_0245_)
  );
  al_nor2 _0763_ (
    .a(_0245_),
    .b(_0244_),
    .y(\DFF_37.D )
  );
  al_and2ft _0764_ (
    .a(\DFF_22.Q ),
    .b(\DFF_24.Q ),
    .y(_0246_)
  );
  al_nand2ft _0765_ (
    .a(\DFF_24.Q ),
    .b(\DFF_22.Q ),
    .y(_0247_)
  );
  al_nand2ft _0766_ (
    .a(_0246_),
    .b(_0247_),
    .y(_0248_)
  );
  al_and2ft _0767_ (
    .a(\DFF_25.Q ),
    .b(\DFF_23.Q ),
    .y(_0249_)
  );
  al_nand2ft _0768_ (
    .a(\DFF_23.Q ),
    .b(\DFF_25.Q ),
    .y(_0250_)
  );
  al_or3ftt _0769_ (
    .a(_0250_),
    .b(_0249_),
    .c(_0197_),
    .y(_0251_)
  );
  al_aoi21ftf _0770_ (
    .a(_0249_),
    .b(_0250_),
    .c(_0197_),
    .y(_0252_)
  );
  al_oai21ftf _0771_ (
    .a(_0251_),
    .b(_0252_),
    .c(_0248_),
    .y(_0253_)
  );
  al_or3fft _0772_ (
    .a(_0248_),
    .b(_0251_),
    .c(_0252_),
    .y(_0254_)
  );
  al_nand3ftt _0773_ (
    .a(\DFF_26.Q ),
    .b(_0193_),
    .c(_0194_),
    .y(_0255_)
  );
  al_ao21ttf _0774_ (
    .a(_0193_),
    .b(_0194_),
    .c(\DFF_26.Q ),
    .y(_0256_)
  );
  al_nand2 _0775_ (
    .a(_0255_),
    .b(_0256_),
    .y(_0257_)
  );
  al_and3 _0776_ (
    .a(_0257_),
    .b(_0254_),
    .c(_0253_),
    .y(_0258_)
  );
  al_ao21 _0777_ (
    .a(_0254_),
    .b(_0253_),
    .c(_0257_),
    .y(_0259_)
  );
  al_nand2ft _0778_ (
    .a(_0258_),
    .b(_0259_),
    .y(\DFF_27.D )
  );
  al_or2 _0779_ (
    .a(n3084gat),
    .b(n3083gat),
    .y(_0260_)
  );
  al_nand2 _0780_ (
    .a(n3084gat),
    .b(n3083gat),
    .y(_0261_)
  );
  al_and3ftt _0781_ (
    .a(n3085gat),
    .b(_0260_),
    .c(_0261_),
    .y(_0262_)
  );
  al_ao21ttf _0782_ (
    .a(_0260_),
    .b(_0261_),
    .c(n3085gat),
    .y(_0263_)
  );
  al_nand2ft _0783_ (
    .a(_0262_),
    .b(_0263_),
    .y(_0264_)
  );
  al_and2ft _0784_ (
    .a(n3087gat),
    .b(n3086gat),
    .y(_0265_)
  );
  al_nand2ft _0785_ (
    .a(n3086gat),
    .b(n3087gat),
    .y(_0266_)
  );
  al_nand2ft _0786_ (
    .a(_0265_),
    .b(_0266_),
    .y(_0267_)
  );
  al_and2ft _0787_ (
    .a(n3089gat),
    .b(n3088gat),
    .y(_0268_)
  );
  al_nand2ft _0788_ (
    .a(n3088gat),
    .b(n3089gat),
    .y(_0269_)
  );
  al_nand3ftt _0789_ (
    .a(_0268_),
    .b(_0269_),
    .c(_0267_),
    .y(_0270_)
  );
  al_ao21ftt _0790_ (
    .a(_0268_),
    .b(_0269_),
    .c(_0267_),
    .y(_0271_)
  );
  al_aoi21ttf _0791_ (
    .a(_0270_),
    .b(_0271_),
    .c(_0264_),
    .y(_0272_)
  );
  al_or3fft _0792_ (
    .a(_0270_),
    .b(_0271_),
    .c(_0264_),
    .y(_0273_)
  );
  al_nand2ft _0793_ (
    .a(_0272_),
    .b(_0273_),
    .y(\DFF_9.D )
  );
  al_inv _0794_ (
    .a(\DFF_132.Q ),
    .y(n3106gat)
  );
  al_aoi21ttf _0795_ (
    .a(\DFF_131.Q ),
    .b(\DFF_168.Q ),
    .c(\DFF_132.Q ),
    .y(n3107gat)
  );
  al_nand2ft _0796_ (
    .a(_0162_),
    .b(_0163_),
    .y(n3116gat)
  );
  al_inv _0797_ (
    .a(\DFF_98.Q ),
    .y(\DFF_124.D )
  );
  al_inv _0798_ (
    .a(\DFF_97.Q ),
    .y(\DFF_123.D )
  );
  al_inv _0799_ (
    .a(\DFF_96.Q ),
    .y(\DFF_125.D )
  );
  al_and3fft _0800_ (
    .a(\DFF_38.Q ),
    .b(\DFF_142.Q ),
    .c(\DFF_39.Q ),
    .y(_0274_)
  );
  al_and3 _0801_ (
    .a(\DFF_40.Q ),
    .b(\DFF_41.Q ),
    .c(_0274_),
    .y(_0275_)
  );
  al_or3 _0802_ (
    .a(\DFF_142.Q ),
    .b(_0193_),
    .c(_0195_),
    .y(_0276_)
  );
  al_nor3ftt _0803_ (
    .a(\DFF_65.Q ),
    .b(_0132_),
    .c(_0129_),
    .y(_0277_)
  );
  al_nor2 _0804_ (
    .a(\DFF_60.Q ),
    .b(\DFF_62.Q ),
    .y(_0278_)
  );
  al_and3ftt _0805_ (
    .a(\DFF_61.Q ),
    .b(\DFF_59.Q ),
    .c(\DFF_58.Q ),
    .y(_0279_)
  );
  al_and3 _0806_ (
    .a(_0278_),
    .b(_0279_),
    .c(_0277_),
    .y(_0280_)
  );
  al_aoi21ftf _0807_ (
    .a(_0275_),
    .b(_0276_),
    .c(_0280_),
    .y(n3138gat)
  );
  al_and2 _0808_ (
    .a(\DFF_40.Q ),
    .b(\DFF_41.Q ),
    .y(_0281_)
  );
  al_aoi21ttf _0809_ (
    .a(_0281_),
    .b(_0274_),
    .c(_0276_),
    .y(_0282_)
  );
  al_and3fft _0810_ (
    .a(\DFF_40.Q ),
    .b(\DFF_142.Q ),
    .c(\DFF_39.Q ),
    .y(_0283_)
  );
  al_nand2 _0811_ (
    .a(\DFF_38.Q ),
    .b(_0283_),
    .y(_0284_)
  );
  al_inv _0812_ (
    .a(\DFF_142.Q ),
    .y(_0285_)
  );
  al_nor3fft _0813_ (
    .a(\DFF_38.Q ),
    .b(\DFF_39.Q ),
    .c(_0195_),
    .y(_0286_)
  );
  al_nand3fft _0814_ (
    .a(\DFF_142.Q ),
    .b(_0194_),
    .c(_0281_),
    .y(_0287_)
  );
  al_aoi21ttf _0815_ (
    .a(_0285_),
    .b(_0286_),
    .c(_0287_),
    .y(_0288_)
  );
  al_nand2 _0816_ (
    .a(_0284_),
    .b(_0288_),
    .y(\DFF_126.D )
  );
  al_and3 _0817_ (
    .a(\DFF_131.Q ),
    .b(\DFF_167.Q ),
    .c(\DFF_168.Q ),
    .y(_0289_)
  );
  al_and3fft _0818_ (
    .a(_0289_),
    .b(\DFF_126.D ),
    .c(_0282_),
    .y(n3145gat)
  );
  al_and3 _0819_ (
    .a(\DFF_140.Q ),
    .b(\DFF_150.Q ),
    .c(\DFF_141.Q ),
    .y(_0290_)
  );
  al_and3 _0820_ (
    .a(\DFF_149.Q ),
    .b(_0290_),
    .c(_0103_),
    .y(_0291_)
  );
  al_aoi21ftf _0821_ (
    .a(n3106gat),
    .b(_0289_),
    .c(_0291_),
    .y(n3146gat)
  );
  al_and2 _0822_ (
    .a(\DFF_38.Q ),
    .b(\DFF_39.Q ),
    .y(_0292_)
  );
  al_and3 _0823_ (
    .a(\DFF_40.Q ),
    .b(\DFF_41.Q ),
    .c(_0292_),
    .y(\DFF_16.D )
  );
  al_and2ft _0824_ (
    .a(n3099gat),
    .b(\DFF_17.Q ),
    .y(\DFF_19.D )
  );
  al_nor2 _0825_ (
    .a(\DFF_22.Q ),
    .b(\DFF_142.Q ),
    .y(\DFF_68.D )
  );
  al_nand2ft _0826_ (
    .a(\DFF_21.Q ),
    .b(\DFF_19.Q ),
    .y(_0293_)
  );
  al_and3 _0827_ (
    .a(\DFF_16.Q ),
    .b(n3100gat),
    .c(_0293_),
    .y(_0294_)
  );
  al_and2 _0828_ (
    .a(\DFF_68.D ),
    .b(_0294_),
    .y(\DFF_70.D )
  );
  al_nand3ftt _0829_ (
    .a(_0275_),
    .b(_0276_),
    .c(_0288_),
    .y(\DFF_119.D )
  );
  al_nor2 _0830_ (
    .a(\DFF_40.Q ),
    .b(\DFF_41.Q ),
    .y(_0295_)
  );
  al_and3fft _0831_ (
    .a(\DFF_142.Q ),
    .b(_0193_),
    .c(_0295_),
    .y(\DFF_102.D )
  );
  al_and3ftt _0832_ (
    .a(\DFF_40.Q ),
    .b(\DFF_41.Q ),
    .c(_0274_),
    .y(\DFF_103.D )
  );
  al_nand3 _0833_ (
    .a(\DFF_102.Q ),
    .b(\DFF_103.Q ),
    .c(\DFF_69.Q ),
    .y(\DFF_104.D )
  );
  al_nand2ft _0834_ (
    .a(\DFF_108.Q ),
    .b(\DFF_107.Q ),
    .y(_0296_)
  );
  al_and3ftt _0835_ (
    .a(\DFF_109.Q ),
    .b(\DFF_105.Q ),
    .c(\DFF_106.Q ),
    .y(_0297_)
  );
  al_nand3fft _0836_ (
    .a(_0296_),
    .b(_0098_),
    .c(_0297_),
    .y(_0298_)
  );
  al_nor2 _0837_ (
    .a(\DFF_108.Q ),
    .b(\DFF_107.Q ),
    .y(_0299_)
  );
  al_and2ft _0838_ (
    .a(\DFF_106.Q ),
    .b(\DFF_109.Q ),
    .y(_0300_)
  );
  al_and3 _0839_ (
    .a(\DFF_105.Q ),
    .b(_0300_),
    .c(_0299_),
    .y(_0301_)
  );
  al_nand2 _0840_ (
    .a(_0098_),
    .b(_0301_),
    .y(_0302_)
  );
  al_and2ft _0841_ (
    .a(\DFF_114.Q ),
    .b(\DFF_113.Q ),
    .y(_0303_)
  );
  al_and3ftt _0842_ (
    .a(\DFF_110.Q ),
    .b(_0105_),
    .c(_0303_),
    .y(_0304_)
  );
  al_aoi21ttf _0843_ (
    .a(_0298_),
    .b(_0302_),
    .c(_0304_),
    .y(\DFF_115.D )
  );
  al_nand3ftt _0844_ (
    .a(\DFF_113.Q ),
    .b(\DFF_114.Q ),
    .c(\DFF_110.Q ),
    .y(_0305_)
  );
  al_nor3fft _0845_ (
    .a(\DFF_112.Q ),
    .b(\DFF_111.Q ),
    .c(_0305_),
    .y(_0306_)
  );
  al_and3ftt _0846_ (
    .a(_0296_),
    .b(_0140_),
    .c(_0306_),
    .y(\DFF_117.D )
  );
  al_and3 _0847_ (
    .a(_0299_),
    .b(_0140_),
    .c(_0304_),
    .y(\DFF_120.D )
  );
  al_inv _0848_ (
    .a(_0282_),
    .y(\DFF_122.D )
  );
  al_and3 _0849_ (
    .a(_0196_),
    .b(_0274_),
    .c(_0294_),
    .y(\DFF_131.D )
  );
  al_and2 _0850_ (
    .a(\DFF_69.Q ),
    .b(\DFF_116.Q ),
    .y(_0307_)
  );
  al_and3fft _0851_ (
    .a(\DFF_113.Q ),
    .b(\DFF_110.Q ),
    .c(\DFF_114.Q ),
    .y(_0308_)
  );
  al_and3fft _0852_ (
    .a(_0193_),
    .b(_0195_),
    .c(_0106_),
    .y(_0309_)
  );
  al_nand3ftt _0853_ (
    .a(\DFF_38.Q ),
    .b(\DFF_39.Q ),
    .c(_0295_),
    .y(_0310_)
  );
  al_nand3ftt _0854_ (
    .a(_0193_),
    .b(_0105_),
    .c(_0196_),
    .y(_0311_)
  );
  al_oa21ftt _0855_ (
    .a(_0114_),
    .b(_0310_),
    .c(_0311_),
    .y(_0312_)
  );
  al_aoi21ftf _0856_ (
    .a(_0309_),
    .b(_0312_),
    .c(_0308_),
    .y(_0313_)
  );
  al_nand3ftt _0857_ (
    .a(_0193_),
    .b(_0281_),
    .c(_0308_),
    .y(_0314_)
  );
  al_aoi21ftf _0858_ (
    .a(_0305_),
    .b(\DFF_16.D ),
    .c(_0314_),
    .y(_0315_)
  );
  al_aoi21ttf _0859_ (
    .a(_0110_),
    .b(_0315_),
    .c(_0109_),
    .y(_0316_)
  );
  al_nand3 _0860_ (
    .a(_0114_),
    .b(_0292_),
    .c(_0295_),
    .y(_0317_)
  );
  al_nand3 _0861_ (
    .a(_0105_),
    .b(_0196_),
    .c(_0292_),
    .y(_0318_)
  );
  al_aoi21ttf _0862_ (
    .a(_0106_),
    .b(_0286_),
    .c(_0318_),
    .y(_0319_)
  );
  al_ao21 _0863_ (
    .a(_0317_),
    .b(_0319_),
    .c(_0305_),
    .y(_0320_)
  );
  al_nand3fft _0864_ (
    .a(_0313_),
    .b(_0316_),
    .c(_0320_),
    .y(_0321_)
  );
  al_and3 _0865_ (
    .a(\DFF_102.Q ),
    .b(\DFF_103.Q ),
    .c(\DFF_69.Q ),
    .y(_0322_)
  );
  al_aoi21 _0866_ (
    .a(_0298_),
    .b(_0302_),
    .c(_0322_),
    .y(_0323_)
  );
  al_aoi21 _0867_ (
    .a(_0323_),
    .b(_0321_),
    .c(_0307_),
    .y(\DFF_146.D )
  );
  al_aoi21ftf _0868_ (
    .a(\DFF_130.Q ),
    .b(\DFF_131.Q ),
    .c(_0101_),
    .y(_0324_)
  );
  al_and2 _0869_ (
    .a(_0324_),
    .b(\DFF_146.D ),
    .y(\DFF_132.D )
  );
  al_and3ftt _0870_ (
    .a(\DFF_105.Q ),
    .b(\DFF_109.Q ),
    .c(\DFF_106.Q ),
    .y(_0325_)
  );
  al_and3fft _0871_ (
    .a(_0296_),
    .b(_0098_),
    .c(_0325_),
    .y(\DFF_134.D )
  );
  al_nand3ftt _0872_ (
    .a(\DFF_141.Q ),
    .b(\DFF_130.Q ),
    .c(_0101_),
    .y(_0326_)
  );
  al_aoi21 _0873_ (
    .a(_0323_),
    .b(_0321_),
    .c(_0326_),
    .y(\DFF_142.D )
  );
  al_and3fft _0874_ (
    .a(\DFF_128.Q ),
    .b(\DFF_143.Q ),
    .c(\DFF_133.D ),
    .y(\DFF_144.D )
  );
  al_aoi21ttf _0875_ (
    .a(\DFF_125.Q ),
    .b(\DFF_123.Q ),
    .c(\DFF_96.D ),
    .y(\DFF_97.D )
  );
  al_or3 _0876_ (
    .a(\DFF_125.Q ),
    .b(\DFF_124.Q ),
    .c(\DFF_123.Q ),
    .y(_0327_)
  );
  al_oa21 _0877_ (
    .a(\DFF_125.Q ),
    .b(\DFF_123.Q ),
    .c(\DFF_124.Q ),
    .y(_0328_)
  );
  al_and3ftt _0878_ (
    .a(_0328_),
    .b(_0327_),
    .c(\DFF_96.D ),
    .y(\DFF_98.D )
  );
  al_oai21ttf _0879_ (
    .a(\DFF_105.Q ),
    .b(_0096_),
    .c(\DFF_109.Q ),
    .y(_0329_)
  );
  al_nand2ft _0880_ (
    .a(\DFF_172.D ),
    .b(_0329_),
    .y(_0330_)
  );
  al_nand3fft _0881_ (
    .a(\DFF_118.Q ),
    .b(\DFF_119.Q ),
    .c(_0098_),
    .y(_0331_)
  );
  al_nand3 _0882_ (
    .a(_0098_),
    .b(_0331_),
    .c(_0301_),
    .y(_0332_)
  );
  al_or2 _0883_ (
    .a(\DFF_121.Q ),
    .b(_0298_),
    .y(_0333_)
  );
  al_nand3ftt _0884_ (
    .a(_0098_),
    .b(\DFF_121.Q ),
    .c(\DFF_172.D ),
    .y(_0334_)
  );
  al_aoi21ftf _0885_ (
    .a(_0331_),
    .b(\DFF_171.D ),
    .c(_0334_),
    .y(_0335_)
  );
  al_and3 _0886_ (
    .a(_0332_),
    .b(_0333_),
    .c(_0335_),
    .y(_0336_)
  );
  al_and3 _0887_ (
    .a(\DFF_96.D ),
    .b(_0330_),
    .c(_0336_),
    .y(\DFF_66.D )
  );
  al_and2 _0888_ (
    .a(\DFF_96.D ),
    .b(_0336_),
    .y(\DFF_63.D )
  );
  al_nand3fft _0889_ (
    .a(\DFF_105.Q ),
    .b(\DFF_106.Q ),
    .c(_0299_),
    .y(_0337_)
  );
  al_and2 _0890_ (
    .a(\DFF_105.Q ),
    .b(_0096_),
    .y(_0338_)
  );
  al_nand2ft _0891_ (
    .a(_0338_),
    .b(_0337_),
    .y(_0339_)
  );
  al_and3ftt _0892_ (
    .a(_0339_),
    .b(\DFF_96.D ),
    .c(_0336_),
    .y(\DFF_67.D )
  );
  al_oa21 _0893_ (
    .a(\DFF_108.Q ),
    .b(\DFF_107.Q ),
    .c(\DFF_106.Q ),
    .y(_0340_)
  );
  al_nor2ft _0894_ (
    .a(_0096_),
    .b(_0340_),
    .y(_0341_)
  );
  al_and3 _0895_ (
    .a(\DFF_96.D ),
    .b(_0341_),
    .c(_0336_),
    .y(\DFF_65.D )
  );
  al_and2 _0896_ (
    .a(\DFF_108.Q ),
    .b(\DFF_107.Q ),
    .y(_0342_)
  );
  al_and3ftt _0897_ (
    .a(_0342_),
    .b(\DFF_96.D ),
    .c(_0336_),
    .y(\DFF_64.D )
  );
  al_oai21 _0898_ (
    .a(\DFF_112.Q ),
    .b(\DFF_111.Q ),
    .c(\DFF_110.Q ),
    .y(_0343_)
  );
  al_and3 _0899_ (
    .a(_0111_),
    .b(_0343_),
    .c(\DFF_61.D ),
    .y(\DFF_58.D )
  );
  al_nor3fft _0900_ (
    .a(_0285_),
    .b(_0294_),
    .c(_0310_),
    .y(\DFF_168.D )
  );
  al_and3 _0901_ (
    .a(\DFF_61.Q ),
    .b(\DFF_59.Q ),
    .c(\DFF_58.Q ),
    .y(_0344_)
  );
  al_and3ftt _0902_ (
    .a(_0121_),
    .b(_0344_),
    .c(_0277_),
    .y(\DFF_169.D )
  );
  al_aoi21ttf _0903_ (
    .a(_0323_),
    .b(_0321_),
    .c(_0301_),
    .y(\DFF_170.D )
  );
  al_and2 _0904_ (
    .a(\DFF_135.D ),
    .b(_0304_),
    .y(\DFF_173.D )
  );
  al_ao21 _0905_ (
    .a(_0104_),
    .b(_0105_),
    .c(_0298_),
    .y(_0345_)
  );
  al_aoi21 _0906_ (
    .a(\DFF_104.D ),
    .b(_0321_),
    .c(_0345_),
    .y(\DFF_174.D )
  );
  al_and3ftt _0907_ (
    .a(\DFF_110.Q ),
    .b(_0106_),
    .c(_0303_),
    .y(_0346_)
  );
  al_and3ftt _0908_ (
    .a(_0337_),
    .b(\DFF_109.Q ),
    .c(_0346_),
    .y(\DFF_176.D )
  );
  al_and2 _0909_ (
    .a(_0301_),
    .b(_0346_),
    .y(\DFF_177.D )
  );
  al_nor3fft _0910_ (
    .a(\DFF_130.Q ),
    .b(_0140_),
    .c(_0296_),
    .y(\DFF_178.D )
  );
  al_nand2 _0911_ (
    .a(n3072gat),
    .b(n3093gat),
    .y(_0347_)
  );
  al_ao21ttf _0912_ (
    .a(n3081gat),
    .b(n3095gat),
    .c(_0347_),
    .y(\DFF_33.D )
  );
  al_nand2 _0913_ (
    .a(n3065gat),
    .b(n3093gat),
    .y(_0348_)
  );
  al_ao21ttf _0914_ (
    .a(n3074gat),
    .b(n3095gat),
    .c(_0348_),
    .y(\DFF_28.D )
  );
  al_nand2 _0915_ (
    .a(n3076gat),
    .b(n3095gat),
    .y(_0349_)
  );
  al_ao21ttf _0916_ (
    .a(n3067gat),
    .b(n3093gat),
    .c(_0349_),
    .y(\DFF_29.D )
  );
  al_nand2 _0917_ (
    .a(n3075gat),
    .b(n3095gat),
    .y(_0350_)
  );
  al_ao21ttf _0918_ (
    .a(n3066gat),
    .b(n3093gat),
    .c(_0350_),
    .y(\DFF_30.D )
  );
  al_nand2 _0919_ (
    .a(n3071gat),
    .b(n3093gat),
    .y(_0351_)
  );
  al_ao21ttf _0920_ (
    .a(n3080gat),
    .b(n3095gat),
    .c(_0351_),
    .y(\DFF_31.D )
  );
  al_nand2 _0921_ (
    .a(n3073gat),
    .b(n3093gat),
    .y(_0352_)
  );
  al_ao21ttf _0922_ (
    .a(n3082gat),
    .b(n3095gat),
    .c(_0352_),
    .y(\DFF_32.D )
  );
  al_nand2 _0923_ (
    .a(n3068gat),
    .b(n3093gat),
    .y(_0353_)
  );
  al_ao21ttf _0924_ (
    .a(n3077gat),
    .b(n3095gat),
    .c(_0353_),
    .y(\DFF_34.D )
  );
  al_nand2 _0925_ (
    .a(n3070gat),
    .b(n3093gat),
    .y(_0354_)
  );
  al_ao21ttf _0926_ (
    .a(n3079gat),
    .b(n3095gat),
    .c(_0354_),
    .y(\DFF_35.D )
  );
  al_nand2 _0927_ (
    .a(n3069gat),
    .b(n3093gat),
    .y(_0355_)
  );
  al_ao21ttf _0928_ (
    .a(n3078gat),
    .b(n3095gat),
    .c(_0355_),
    .y(\DFF_36.D )
  );
  al_and3fft _0929_ (
    .a(n3084gat),
    .b(n3083gat),
    .c(n3093gat),
    .y(_0356_)
  );
  al_nand2ft _0930_ (
    .a(n3088gat),
    .b(n3087gat),
    .y(_0357_)
  );
  al_nor3fft _0931_ (
    .a(\DFF_132.Q ),
    .b(_0356_),
    .c(_0357_),
    .y(_0358_)
  );
  al_or2 _0932_ (
    .a(n3091gat),
    .b(n3092gat),
    .y(_0359_)
  );
  al_and3ftt _0933_ (
    .a(n3086gat),
    .b(n3085gat),
    .c(_0359_),
    .y(_0360_)
  );
  al_and3 _0934_ (
    .a(n3065gat),
    .b(_0360_),
    .c(_0358_),
    .y(_0361_)
  );
  al_or3 _0935_ (
    .a(n3085gat),
    .b(n3084gat),
    .c(n3083gat),
    .y(_0362_)
  );
  al_nand2 _0936_ (
    .a(n3086gat),
    .b(n3095gat),
    .y(_0363_)
  );
  al_and2 _0937_ (
    .a(n3094gat),
    .b(\DFF_132.Q ),
    .y(_0364_)
  );
  al_nand3fft _0938_ (
    .a(_0362_),
    .b(_0363_),
    .c(_0364_),
    .y(_0365_)
  );
  al_and3fft _0939_ (
    .a(n3087gat),
    .b(_0365_),
    .c(n3088gat),
    .y(_0366_)
  );
  al_ao21 _0940_ (
    .a(n3074gat),
    .b(_0366_),
    .c(_0361_),
    .y(\DFF_48.D )
  );
  al_and3 _0941_ (
    .a(n3067gat),
    .b(_0360_),
    .c(_0358_),
    .y(_0367_)
  );
  al_ao21 _0942_ (
    .a(n3076gat),
    .b(_0366_),
    .c(_0367_),
    .y(\DFF_49.D )
  );
  al_and3 _0943_ (
    .a(n3066gat),
    .b(_0360_),
    .c(_0358_),
    .y(_0368_)
  );
  al_ao21 _0944_ (
    .a(n3075gat),
    .b(_0366_),
    .c(_0368_),
    .y(\DFF_50.D )
  );
  al_and3 _0945_ (
    .a(n3068gat),
    .b(_0360_),
    .c(_0358_),
    .y(_0369_)
  );
  al_ao21 _0946_ (
    .a(n3077gat),
    .b(_0366_),
    .c(_0369_),
    .y(\DFF_54.D )
  );
  al_nand3 _0947_ (
    .a(n3085gat),
    .b(n3086gat),
    .c(_0359_),
    .y(_0370_)
  );
  al_and2ft _0948_ (
    .a(n3087gat),
    .b(n3088gat),
    .y(_0371_)
  );
  al_and3 _0949_ (
    .a(\DFF_132.Q ),
    .b(_0356_),
    .c(_0371_),
    .y(_0372_)
  );
  al_inv _0950_ (
    .a(n3088gat),
    .y(_0373_)
  );
  al_and2 _0951_ (
    .a(n3095gat),
    .b(\DFF_132.Q ),
    .y(_0374_)
  );
  al_and2 _0952_ (
    .a(n3086gat),
    .b(n3094gat),
    .y(_0375_)
  );
  al_and3ftt _0953_ (
    .a(_0362_),
    .b(_0374_),
    .c(_0375_),
    .y(_0376_)
  );
  al_nand2 _0954_ (
    .a(n3087gat),
    .b(n3095gat),
    .y(_0377_)
  );
  al_nor3ftt _0955_ (
    .a(\DFF_132.Q ),
    .b(_0362_),
    .c(_0377_),
    .y(_0378_)
  );
  al_nand3 _0956_ (
    .a(_0373_),
    .b(_0378_),
    .c(_0376_),
    .y(_0379_)
  );
  al_aoi21ftf _0957_ (
    .a(_0370_),
    .b(_0372_),
    .c(_0379_),
    .y(_0380_)
  );
  al_or3ftt _0958_ (
    .a(\DFF_66.Q ),
    .b(\DFF_65.Q ),
    .c(\DFF_62.Q ),
    .y(_0381_)
  );
  al_aoi21 _0959_ (
    .a(_0279_),
    .b(_0278_),
    .c(_0381_),
    .y(_0382_)
  );
  al_and3ftt _0960_ (
    .a(\DFF_59.Q ),
    .b(\DFF_61.Q ),
    .c(\DFF_58.Q ),
    .y(_0383_)
  );
  al_nand3fft _0961_ (
    .a(\DFF_60.Q ),
    .b(\DFF_62.Q ),
    .c(_0383_),
    .y(_0384_)
  );
  al_and2 _0962_ (
    .a(\DFF_71.Q ),
    .b(\DFF_67.Q ),
    .y(_0385_)
  );
  al_nand3fft _0963_ (
    .a(\DFF_71.Q ),
    .b(\DFF_67.Q ),
    .c(_0131_),
    .y(_0386_)
  );
  al_ao21ftf _0964_ (
    .a(_0132_),
    .b(_0385_),
    .c(_0386_),
    .y(_0387_)
  );
  al_and3 _0965_ (
    .a(_0384_),
    .b(_0382_),
    .c(_0387_),
    .y(_0388_)
  );
  al_ao21ttf _0966_ (
    .a(_0282_),
    .b(_0288_),
    .c(_0388_),
    .y(_0389_)
  );
  al_oai21ftt _0967_ (
    .a(n3065gat),
    .b(_0380_),
    .c(_0389_),
    .y(\DFF_72.D )
  );
  al_oai21ftt _0968_ (
    .a(n3067gat),
    .b(_0380_),
    .c(_0389_),
    .y(\DFF_73.D )
  );
  al_oai21ftt _0969_ (
    .a(n3066gat),
    .b(_0380_),
    .c(_0389_),
    .y(\DFF_74.D )
  );
  al_oai21ftt _0970_ (
    .a(n3071gat),
    .b(_0380_),
    .c(_0389_),
    .y(\DFF_75.D )
  );
  al_oai21ftt _0971_ (
    .a(n3072gat),
    .b(_0380_),
    .c(_0389_),
    .y(\DFF_76.D )
  );
  al_oai21ftt _0972_ (
    .a(n3068gat),
    .b(_0380_),
    .c(_0389_),
    .y(\DFF_77.D )
  );
  al_oai21ftt _0973_ (
    .a(n3070gat),
    .b(_0380_),
    .c(_0389_),
    .y(\DFF_78.D )
  );
  al_oai21ftt _0974_ (
    .a(n3069gat),
    .b(_0380_),
    .c(_0389_),
    .y(\DFF_79.D )
  );
  al_oai21ftt _0975_ (
    .a(n3073gat),
    .b(_0380_),
    .c(_0389_),
    .y(\DFF_80.D )
  );
  al_ao21 _0976_ (
    .a(_0388_),
    .b(\DFF_119.D ),
    .c(\DFF_32.D ),
    .y(\DFF_82.D )
  );
  al_ao21 _0977_ (
    .a(_0388_),
    .b(\DFF_119.D ),
    .c(\DFF_28.D ),
    .y(\DFF_83.D )
  );
  al_ao21 _0978_ (
    .a(_0388_),
    .b(\DFF_119.D ),
    .c(\DFF_29.D ),
    .y(\DFF_84.D )
  );
  al_ao21 _0979_ (
    .a(_0388_),
    .b(\DFF_119.D ),
    .c(\DFF_30.D ),
    .y(\DFF_85.D )
  );
  al_ao21 _0980_ (
    .a(_0388_),
    .b(\DFF_119.D ),
    .c(\DFF_31.D ),
    .y(\DFF_86.D )
  );
  al_ao21 _0981_ (
    .a(_0388_),
    .b(\DFF_119.D ),
    .c(\DFF_33.D ),
    .y(\DFF_87.D )
  );
  al_ao21 _0982_ (
    .a(_0388_),
    .b(\DFF_119.D ),
    .c(\DFF_34.D ),
    .y(\DFF_88.D )
  );
  al_ao21 _0983_ (
    .a(_0388_),
    .b(\DFF_119.D ),
    .c(\DFF_35.D ),
    .y(\DFF_89.D )
  );
  al_ao21 _0984_ (
    .a(_0388_),
    .b(\DFF_119.D ),
    .c(\DFF_36.D ),
    .y(\DFF_90.D )
  );
  al_nand3ftt _0985_ (
    .a(n3090gat),
    .b(\DFF_81.Q ),
    .c(\DFF_91.Q ),
    .y(_0390_)
  );
  al_nand2 _0986_ (
    .a(\DFF_27.Q ),
    .b(\DFF_37.Q ),
    .y(_0391_)
  );
  al_and2 _0987_ (
    .a(\DFF_47.Q ),
    .b(\DFF_57.Q ),
    .y(_0392_)
  );
  al_nand3fft _0988_ (
    .a(_0390_),
    .b(_0391_),
    .c(_0392_),
    .y(\DFF_92.D )
  );
  al_nand3 _0989_ (
    .a(_0284_),
    .b(_0282_),
    .c(_0288_),
    .y(\DFF_143.D )
  );
  al_oa21 _0990_ (
    .a(\DFF_122.Q ),
    .b(_0327_),
    .c(\DFF_126.Q ),
    .y(_0393_)
  );
  al_and3fft _0991_ (
    .a(_0393_),
    .b(_0336_),
    .c(_0108_),
    .y(\DFF_127.D )
  );
  al_inv _0992_ (
    .a(\DFF_157.Q ),
    .y(_0394_)
  );
  al_oai21ttf _0993_ (
    .a(\DFF_156.Q ),
    .b(_0276_),
    .c(_0394_),
    .y(_0395_)
  );
  al_and3fft _0994_ (
    .a(\DFF_156.Q ),
    .b(_0276_),
    .c(_0394_),
    .y(_0396_)
  );
  al_and2ft _0995_ (
    .a(_0396_),
    .b(_0395_),
    .y(_0397_)
  );
  al_and3 _0996_ (
    .a(n3088gat),
    .b(\DFF_132.Q ),
    .c(_0356_),
    .y(_0398_)
  );
  al_nand3 _0997_ (
    .a(n3087gat),
    .b(_0360_),
    .c(_0398_),
    .y(_0399_)
  );
  al_aoi21ttf _0998_ (
    .a(_0371_),
    .b(_0376_),
    .c(_0399_),
    .y(_0400_)
  );
  al_mux2h _0999_ (
    .a(n3067gat),
    .b(_0397_),
    .s(_0400_),
    .y(\DFF_43.D )
  );
  al_or2 _1000_ (
    .a(\DFF_156.Q ),
    .b(_0276_),
    .y(_0401_)
  );
  al_and2 _1001_ (
    .a(\DFF_156.Q ),
    .b(_0276_),
    .y(_0402_)
  );
  al_and2ft _1002_ (
    .a(_0402_),
    .b(_0401_),
    .y(_0403_)
  );
  al_mux2h _1003_ (
    .a(n3068gat),
    .b(_0403_),
    .s(_0400_),
    .y(\DFF_46.D )
  );
  al_nand2 _1004_ (
    .a(_0360_),
    .b(_0358_),
    .y(_0404_)
  );
  al_aoi21ftf _1005_ (
    .a(_0365_),
    .b(_0371_),
    .c(_0404_),
    .y(_0405_)
  );
  al_inv _1006_ (
    .a(\DFF_159.Q ),
    .y(_0406_)
  );
  al_inv _1007_ (
    .a(\DFF_158.Q ),
    .y(_0407_)
  );
  al_and3 _1008_ (
    .a(_0406_),
    .b(_0407_),
    .c(_0275_),
    .y(_0408_)
  );
  al_ao21 _1009_ (
    .a(_0406_),
    .b(_0275_),
    .c(_0407_),
    .y(_0409_)
  );
  al_and2ft _1010_ (
    .a(_0408_),
    .b(_0409_),
    .y(_0410_)
  );
  al_and3 _1011_ (
    .a(n3071gat),
    .b(_0360_),
    .c(_0358_),
    .y(_0411_)
  );
  al_ao21 _1012_ (
    .a(n3080gat),
    .b(_0366_),
    .c(_0411_),
    .y(_0412_)
  );
  al_ao21 _1013_ (
    .a(_0405_),
    .b(_0410_),
    .c(_0412_),
    .y(\DFF_51.D )
  );
  al_and3ftt _1014_ (
    .a(\DFF_159.Q ),
    .b(_0274_),
    .c(_0281_),
    .y(_0413_)
  );
  al_ao21 _1015_ (
    .a(_0274_),
    .b(_0281_),
    .c(_0406_),
    .y(_0414_)
  );
  al_and2ft _1016_ (
    .a(_0413_),
    .b(_0414_),
    .y(_0415_)
  );
  al_and3 _1017_ (
    .a(n3072gat),
    .b(_0360_),
    .c(_0358_),
    .y(_0416_)
  );
  al_aoi21 _1018_ (
    .a(n3081gat),
    .b(_0366_),
    .c(_0416_),
    .y(_0417_)
  );
  al_ao21ttf _1019_ (
    .a(_0415_),
    .b(_0405_),
    .c(_0417_),
    .y(\DFF_53.D )
  );
  al_oai21ftf _1020_ (
    .a(\DFF_161.Q ),
    .b(\DFF_158.Q ),
    .c(\DFF_159.Q ),
    .y(_0418_)
  );
  al_and3 _1021_ (
    .a(\DFF_160.Q ),
    .b(_0418_),
    .c(_0275_),
    .y(_0419_)
  );
  al_ao21 _1022_ (
    .a(_0418_),
    .b(_0275_),
    .c(\DFF_160.Q ),
    .y(_0420_)
  );
  al_nand2ft _1023_ (
    .a(_0419_),
    .b(_0420_),
    .y(_0421_)
  );
  al_or3fft _1024_ (
    .a(n3082gat),
    .b(_0371_),
    .c(_0365_),
    .y(_0422_)
  );
  al_oai21ftt _1025_ (
    .a(n3073gat),
    .b(_0404_),
    .c(_0422_),
    .y(_0423_)
  );
  al_ao21 _1026_ (
    .a(_0421_),
    .b(_0405_),
    .c(_0423_),
    .y(\DFF_52.D )
  );
  al_inv _1027_ (
    .a(\DFF_161.Q ),
    .y(_0424_)
  );
  al_and3 _1028_ (
    .a(_0407_),
    .b(_0424_),
    .c(_0413_),
    .y(_0425_)
  );
  al_ao21 _1029_ (
    .a(_0407_),
    .b(_0413_),
    .c(_0424_),
    .y(_0426_)
  );
  al_and2ft _1030_ (
    .a(_0425_),
    .b(_0426_),
    .y(_0427_)
  );
  al_and3 _1031_ (
    .a(n3070gat),
    .b(_0360_),
    .c(_0358_),
    .y(_0428_)
  );
  al_aoi21 _1032_ (
    .a(n3079gat),
    .b(_0366_),
    .c(_0428_),
    .y(_0429_)
  );
  al_ao21ttf _1033_ (
    .a(_0405_),
    .b(_0427_),
    .c(_0429_),
    .y(\DFF_55.D )
  );
  al_ao21ftf _1034_ (
    .a(\DFF_162.Q ),
    .b(_0425_),
    .c(_0405_),
    .y(_0430_)
  );
  al_ao21ftt _1035_ (
    .a(_0425_),
    .b(\DFF_162.Q ),
    .c(_0430_),
    .y(_0431_)
  );
  al_and3 _1036_ (
    .a(n3078gat),
    .b(_0371_),
    .c(_0376_),
    .y(_0432_)
  );
  al_oa21ftf _1037_ (
    .a(n3069gat),
    .b(_0404_),
    .c(_0432_),
    .y(_0433_)
  );
  al_nand2 _1038_ (
    .a(_0433_),
    .b(_0431_),
    .y(\DFF_56.D )
  );
  al_oa21ftf _1039_ (
    .a(\DFF_163.Q ),
    .b(\DFF_157.Q ),
    .c(\DFF_156.Q ),
    .y(_0434_)
  );
  al_and3fft _1040_ (
    .a(_0434_),
    .b(_0276_),
    .c(\DFF_164.Q ),
    .y(_0435_)
  );
  al_oai21ttf _1041_ (
    .a(_0434_),
    .b(_0276_),
    .c(\DFF_164.Q ),
    .y(_0436_)
  );
  al_nand2ft _1042_ (
    .a(_0435_),
    .b(_0436_),
    .y(_0437_)
  );
  al_mux2h _1043_ (
    .a(n3073gat),
    .b(_0437_),
    .s(_0400_),
    .y(\DFF_45.D )
  );
  al_inv _1044_ (
    .a(\DFF_163.Q ),
    .y(_0438_)
  );
  al_nand2 _1045_ (
    .a(_0438_),
    .b(_0396_),
    .y(_0439_)
  );
  al_or2 _1046_ (
    .a(_0438_),
    .b(_0396_),
    .y(_0440_)
  );
  al_nand3 _1047_ (
    .a(_0400_),
    .b(_0439_),
    .c(_0440_),
    .y(_0441_)
  );
  al_ao21ftf _1048_ (
    .a(_0400_),
    .b(n3066gat),
    .c(_0441_),
    .y(\DFF_44.D )
  );
  al_nand3fft _1049_ (
    .a(\DFF_163.Q ),
    .b(\DFF_165.Q ),
    .c(_0396_),
    .y(_0442_)
  );
  al_ao21ttf _1050_ (
    .a(_0438_),
    .b(_0396_),
    .c(\DFF_165.Q ),
    .y(_0443_)
  );
  al_nand3 _1051_ (
    .a(_0400_),
    .b(_0442_),
    .c(_0443_),
    .y(_0444_)
  );
  al_ao21ftf _1052_ (
    .a(_0400_),
    .b(n3065gat),
    .c(_0444_),
    .y(\DFF_42.D )
  );
  al_nand3ftt _1053_ (
    .a(n3085gat),
    .b(_0265_),
    .c(_0398_),
    .y(_0445_)
  );
  al_nand3fft _1054_ (
    .a(n3088gat),
    .b(n3086gat),
    .c(_0378_),
    .y(_0446_)
  );
  al_nand3 _1055_ (
    .a(_0342_),
    .b(_0445_),
    .c(_0446_),
    .y(n3151gat)
  );
  al_inv _1056_ (
    .a(\DFF_24.Q ),
    .y(_0447_)
  );
  al_ao21ftt _1057_ (
    .a(\DFF_142.Q ),
    .b(_0447_),
    .c(_0341_),
    .y(n3150gat)
  );
  al_nand2ft _1058_ (
    .a(\DFF_84.Q ),
    .b(_0383_),
    .y(_0448_)
  );
  al_nand2ft _1059_ (
    .a(\DFF_85.Q ),
    .b(_0279_),
    .y(_0449_)
  );
  al_and3ftt _1060_ (
    .a(\DFF_58.Q ),
    .b(\DFF_61.Q ),
    .c(\DFF_59.Q ),
    .y(_0450_)
  );
  al_nand2ft _1061_ (
    .a(\DFF_90.Q ),
    .b(_0450_),
    .y(_0451_)
  );
  al_aoi21ftf _1062_ (
    .a(\DFF_83.Q ),
    .b(_0344_),
    .c(_0451_),
    .y(_0452_)
  );
  al_and3 _1063_ (
    .a(_0448_),
    .b(_0449_),
    .c(_0452_),
    .y(_0453_)
  );
  al_and3fft _1064_ (
    .a(\DFF_61.Q ),
    .b(\DFF_59.Q ),
    .c(\DFF_58.Q ),
    .y(_0454_)
  );
  al_and3fft _1065_ (
    .a(\DFF_59.Q ),
    .b(\DFF_58.Q ),
    .c(\DFF_61.Q ),
    .y(_0455_)
  );
  al_nand2ft _1066_ (
    .a(\DFF_86.Q ),
    .b(_0455_),
    .y(_0456_)
  );
  al_aoi21ftf _1067_ (
    .a(\DFF_88.Q ),
    .b(_0454_),
    .c(_0456_),
    .y(_0457_)
  );
  al_or3 _1068_ (
    .a(\DFF_61.Q ),
    .b(\DFF_59.Q ),
    .c(\DFF_58.Q ),
    .y(_0458_)
  );
  al_or2 _1069_ (
    .a(\DFF_87.Q ),
    .b(_0458_),
    .y(_0459_)
  );
  al_and3fft _1070_ (
    .a(\DFF_61.Q ),
    .b(\DFF_58.Q ),
    .c(\DFF_59.Q ),
    .y(_0460_)
  );
  al_nand2ft _1071_ (
    .a(\DFF_89.Q ),
    .b(_0460_),
    .y(_0461_)
  );
  al_and3 _1072_ (
    .a(_0459_),
    .b(_0461_),
    .c(_0457_),
    .y(_0462_)
  );
  al_ao21 _1073_ (
    .a(_0453_),
    .b(_0462_),
    .c(_0121_),
    .y(_0463_)
  );
  al_nand3ftt _1074_ (
    .a(\DFF_142.Q ),
    .b(_0295_),
    .c(_0292_),
    .y(_0464_)
  );
  al_nand3ftt _1075_ (
    .a(_0464_),
    .b(_0185_),
    .c(_0186_),
    .y(_0465_)
  );
  al_nand3 _1076_ (
    .a(_0464_),
    .b(_0183_),
    .c(_0182_),
    .y(_0466_)
  );
  al_nand3fft _1077_ (
    .a(\DFF_60.Q ),
    .b(\DFF_62.Q ),
    .c(_0344_),
    .y(_0467_)
  );
  al_ao21 _1078_ (
    .a(_0466_),
    .b(_0465_),
    .c(_0467_),
    .y(_0468_)
  );
  al_ao21 _1079_ (
    .a(_0463_),
    .b(_0468_),
    .c(_0284_),
    .y(_0469_)
  );
  al_and2 _1080_ (
    .a(\DFF_60.Q ),
    .b(\DFF_62.Q ),
    .y(_0470_)
  );
  al_and3ftt _1081_ (
    .a(\DFF_36.Q ),
    .b(\DFF_60.Q ),
    .c(\DFF_62.Q ),
    .y(_0471_)
  );
  al_ao21 _1082_ (
    .a(_0471_),
    .b(_0455_),
    .c(_0322_),
    .y(_0472_)
  );
  al_nand2ft _1083_ (
    .a(\DFF_43.Q ),
    .b(_0450_),
    .y(_0473_)
  );
  al_aoi21ftf _1084_ (
    .a(\DFF_46.Q ),
    .b(_0460_),
    .c(_0473_),
    .y(_0474_)
  );
  al_nand2ft _1085_ (
    .a(\DFF_42.Q ),
    .b(_0383_),
    .y(_0475_)
  );
  al_aoi21ftf _1086_ (
    .a(\DFF_44.Q ),
    .b(_0454_),
    .c(_0475_),
    .y(_0476_)
  );
  al_ao21ttf _1087_ (
    .a(_0474_),
    .b(_0476_),
    .c(_0472_),
    .y(_0477_)
  );
  al_nand2ft _1088_ (
    .a(\DFF_31.Q ),
    .b(_0344_),
    .y(_0478_)
  );
  al_and2ft _1089_ (
    .a(\DFF_23.Q ),
    .b(_0450_),
    .y(_0479_)
  );
  al_nand2ft _1090_ (
    .a(\DFF_26.Q ),
    .b(_0460_),
    .y(_0480_)
  );
  al_and3ftt _1091_ (
    .a(_0479_),
    .b(_0478_),
    .c(_0480_),
    .y(_0481_)
  );
  al_nand2ft _1092_ (
    .a(\DFF_33.Q ),
    .b(_0279_),
    .y(_0482_)
  );
  al_and2ft _1093_ (
    .a(\DFF_22.Q ),
    .b(_0383_),
    .y(_0483_)
  );
  al_aoi21ftf _1094_ (
    .a(\DFF_24.Q ),
    .b(_0454_),
    .c(\DFF_104.D ),
    .y(_0484_)
  );
  al_and3ftt _1095_ (
    .a(_0483_),
    .b(_0482_),
    .c(_0484_),
    .y(_0485_)
  );
  al_aoi21ftf _1096_ (
    .a(\DFF_53.Q ),
    .b(_0279_),
    .c(_0322_),
    .y(_0486_)
  );
  al_aoi21ftf _1097_ (
    .a(\DFF_51.Q ),
    .b(_0344_),
    .c(_0486_),
    .y(_0487_)
  );
  al_ao21 _1098_ (
    .a(_0481_),
    .b(_0485_),
    .c(_0487_),
    .y(_0488_)
  );
  al_ao21 _1099_ (
    .a(_0477_),
    .b(_0488_),
    .c(_0122_),
    .y(_0489_)
  );
  al_nand2ft _1100_ (
    .a(\DFF_29.Q ),
    .b(_0450_),
    .y(_0490_)
  );
  al_aoi21ftf _1101_ (
    .a(\DFF_34.Q ),
    .b(_0460_),
    .c(_0490_),
    .y(_0491_)
  );
  al_nand2ft _1102_ (
    .a(\DFF_28.Q ),
    .b(_0383_),
    .y(_0492_)
  );
  al_aoi21ftf _1103_ (
    .a(\DFF_30.Q ),
    .b(_0454_),
    .c(_0492_),
    .y(_0493_)
  );
  al_aoi21 _1104_ (
    .a(_0491_),
    .b(_0493_),
    .c(_0322_),
    .y(_0494_)
  );
  al_nand2 _1105_ (
    .a(\DFF_35.Q ),
    .b(\DFF_104.D ),
    .y(_0495_)
  );
  al_nand2 _1106_ (
    .a(\DFF_55.Q ),
    .b(_0322_),
    .y(_0496_)
  );
  al_and3ftt _1107_ (
    .a(_0458_),
    .b(_0495_),
    .c(_0496_),
    .y(_0497_)
  );
  al_ao21ttf _1108_ (
    .a(\DFF_104.Q ),
    .b(_0287_),
    .c(_0344_),
    .y(_0498_)
  );
  al_ao21ttf _1109_ (
    .a(_0284_),
    .b(_0287_),
    .c(_0279_),
    .y(_0499_)
  );
  al_nand3ftt _1110_ (
    .a(_0497_),
    .b(_0498_),
    .c(_0499_),
    .y(_0500_)
  );
  al_aoi21ttf _1111_ (
    .a(\DFF_56.Q ),
    .b(_0322_),
    .c(_0455_),
    .y(_0501_)
  );
  al_nand2ft _1112_ (
    .a(\DFF_49.Q ),
    .b(_0450_),
    .y(_0502_)
  );
  al_ao21ftf _1113_ (
    .a(\DFF_54.Q ),
    .b(_0460_),
    .c(_0502_),
    .y(_0503_)
  );
  al_nand2ft _1114_ (
    .a(\DFF_48.Q ),
    .b(_0383_),
    .y(_0504_)
  );
  al_aoi21ftf _1115_ (
    .a(\DFF_50.Q ),
    .b(_0454_),
    .c(_0504_),
    .y(_0505_)
  );
  al_nand3fft _1116_ (
    .a(_0501_),
    .b(_0503_),
    .c(_0505_),
    .y(_0506_)
  );
  al_nand2 _1117_ (
    .a(_0472_),
    .b(_0506_),
    .y(_0507_)
  );
  al_nand3fft _1118_ (
    .a(_0494_),
    .b(_0500_),
    .c(_0507_),
    .y(_0508_)
  );
  al_ao21ttf _1119_ (
    .a(_0470_),
    .b(_0508_),
    .c(_0489_),
    .y(_0509_)
  );
  al_nand3fft _1120_ (
    .a(\DFF_133.Q ),
    .b(\DFF_33.Q ),
    .c(\DFF_132.Q ),
    .y(_0510_)
  );
  al_or3 _1121_ (
    .a(\DFF_134.Q ),
    .b(_0322_),
    .c(_0098_),
    .y(_0511_)
  );
  al_nand3ftt _1122_ (
    .a(\DFF_135.Q ),
    .b(\DFF_104.D ),
    .c(_0098_),
    .y(_0512_)
  );
  al_ao21 _1123_ (
    .a(_0512_),
    .b(_0511_),
    .c(\DFF_117.Q ),
    .y(_0513_)
  );
  al_nand2 _1124_ (
    .a(_0510_),
    .b(_0513_),
    .y(_0514_)
  );
  al_aoi21 _1125_ (
    .a(\DFF_115.Q ),
    .b(_0509_),
    .c(_0514_),
    .y(_0515_)
  );
  al_nand3 _1126_ (
    .a(\DFF_94.D ),
    .b(_0515_),
    .c(_0469_),
    .y(n3144gat)
  );
  al_nand3 _1127_ (
    .a(\DFF_101.D ),
    .b(_0515_),
    .c(_0469_),
    .y(n3143gat)
  );
  al_nor2 _1128_ (
    .a(_0322_),
    .b(_0098_),
    .y(_0516_)
  );
  al_and3ftt _1129_ (
    .a(\DFF_173.Q ),
    .b(\DFF_71.D ),
    .c(\DFF_143.D ),
    .y(_0517_)
  );
  al_oai21ttf _1130_ (
    .a(_0516_),
    .b(_0517_),
    .c(\DFF_174.Q ),
    .y(_0518_)
  );
  al_ao21ttf _1131_ (
    .a(_0322_),
    .b(_0284_),
    .c(_0098_),
    .y(_0519_)
  );
  al_nor2 _1132_ (
    .a(\DFF_170.Q ),
    .b(_0519_),
    .y(_0520_)
  );
  al_and3fft _1133_ (
    .a(\DFF_172.Q ),
    .b(_0098_),
    .c(\DFF_173.Q ),
    .y(_0521_)
  );
  al_or2 _1134_ (
    .a(\DFF_117.Q ),
    .b(\DFF_171.Q ),
    .y(_0522_)
  );
  al_ao21ftf _1135_ (
    .a(\DFF_170.Q ),
    .b(\DFF_169.Q ),
    .c(_0522_),
    .y(_0523_)
  );
  al_nand3 _1136_ (
    .a(_0098_),
    .b(_0523_),
    .c(\DFF_119.D ),
    .y(_0524_)
  );
  al_nand3fft _1137_ (
    .a(_0520_),
    .b(_0521_),
    .c(_0524_),
    .y(_0525_)
  );
  al_nand2ft _1138_ (
    .a(_0525_),
    .b(_0518_),
    .y(n3141gat)
  );
  al_oa21 _1139_ (
    .a(n3085gat),
    .b(n3086gat),
    .c(_0356_),
    .y(_0526_)
  );
  al_and2 _1140_ (
    .a(n3088gat),
    .b(n3087gat),
    .y(_0527_)
  );
  al_nand3fft _1141_ (
    .a(_0362_),
    .b(_0363_),
    .c(_0527_),
    .y(_0528_)
  );
  al_aoi21ftf _1142_ (
    .a(n3088gat),
    .b(_0526_),
    .c(_0528_),
    .y(_0529_)
  );
  al_nand2 _1143_ (
    .a(n3087gat),
    .b(n3093gat),
    .y(_0530_)
  );
  al_aoi21ttf _1144_ (
    .a(n3088gat),
    .b(n3095gat),
    .c(_0530_),
    .y(_0531_)
  );
  al_ao21ttf _1145_ (
    .a(n3086gat),
    .b(n3093gat),
    .c(_0377_),
    .y(_0532_)
  );
  al_ao21ttf _1146_ (
    .a(n3085gat),
    .b(n3093gat),
    .c(_0363_),
    .y(_0533_)
  );
  al_and3fft _1147_ (
    .a(_0532_),
    .b(_0531_),
    .c(_0533_),
    .y(_0534_)
  );
  al_and3ftt _1148_ (
    .a(_0531_),
    .b(_0532_),
    .c(_0533_),
    .y(_0535_)
  );
  al_or3ftt _1149_ (
    .a(_0532_),
    .b(\DFF_33.Q ),
    .c(_0533_),
    .y(_0536_)
  );
  al_and3 _1150_ (
    .a(_0532_),
    .b(_0531_),
    .c(_0533_),
    .y(_0537_)
  );
  al_aoi21ftf _1151_ (
    .a(\DFF_87.Q ),
    .b(_0537_),
    .c(_0536_),
    .y(_0538_)
  );
  al_aoi21ftf _1152_ (
    .a(\DFF_41.Q ),
    .b(_0535_),
    .c(_0538_),
    .y(_0539_)
  );
  al_ao21ftf _1153_ (
    .a(\DFF_53.Q ),
    .b(_0534_),
    .c(_0539_),
    .y(_0540_)
  );
  al_nand2ft _1154_ (
    .a(\DFF_76.Q ),
    .b(_0537_),
    .y(_0541_)
  );
  al_or3ftt _1155_ (
    .a(_0532_),
    .b(_0531_),
    .c(_0533_),
    .y(_0542_)
  );
  al_oai21ftf _1156_ (
    .a(_0542_),
    .b(_0534_),
    .c(\DFF_41.Q ),
    .y(_0543_)
  );
  al_ao21 _1157_ (
    .a(_0363_),
    .b(_0377_),
    .c(_0362_),
    .y(_0544_)
  );
  al_nand3 _1158_ (
    .a(n3085gat),
    .b(n3087gat),
    .c(n3086gat),
    .y(_0545_)
  );
  al_and3 _1159_ (
    .a(n3088gat),
    .b(n3093gat),
    .c(_0545_),
    .y(_0546_)
  );
  al_aoi21ttf _1160_ (
    .a(_0546_),
    .b(_0526_),
    .c(_0544_),
    .y(_0547_)
  );
  al_ao21 _1161_ (
    .a(_0541_),
    .b(_0543_),
    .c(_0547_),
    .y(_0548_)
  );
  al_ao21ftf _1162_ (
    .a(_0529_),
    .b(_0540_),
    .c(_0548_),
    .y(n3137gat)
  );
  al_nand2 _1163_ (
    .a(\DFF_158.D ),
    .b(_0534_),
    .y(_0549_)
  );
  al_aoi21ftf _1164_ (
    .a(\DFF_40.Q ),
    .b(_0535_),
    .c(_0549_),
    .y(_0550_)
  );
  al_nand2ft _1165_ (
    .a(\DFF_86.Q ),
    .b(_0537_),
    .y(_0551_)
  );
  al_and2ft _1166_ (
    .a(_0533_),
    .b(_0532_),
    .y(_0552_)
  );
  al_nand3fft _1167_ (
    .a(\DFF_31.Q ),
    .b(_0531_),
    .c(_0552_),
    .y(_0000_)
  );
  al_nand3 _1168_ (
    .a(_0551_),
    .b(_0000_),
    .c(_0550_),
    .y(_0001_)
  );
  al_nand2ft _1169_ (
    .a(\DFF_75.Q ),
    .b(_0537_),
    .y(_0002_)
  );
  al_oai21ftf _1170_ (
    .a(_0542_),
    .b(_0534_),
    .c(\DFF_40.Q ),
    .y(_0003_)
  );
  al_ao21 _1171_ (
    .a(_0002_),
    .b(_0003_),
    .c(_0547_),
    .y(_0004_)
  );
  al_ao21ftf _1172_ (
    .a(_0529_),
    .b(_0001_),
    .c(_0004_),
    .y(n3136gat)
  );
  al_nand2ft _1173_ (
    .a(\DFF_78.Q ),
    .b(_0537_),
    .y(_0005_)
  );
  al_oai21ftf _1174_ (
    .a(_0542_),
    .b(_0534_),
    .c(\DFF_38.Q ),
    .y(_0006_)
  );
  al_ao21 _1175_ (
    .a(_0005_),
    .b(_0006_),
    .c(_0547_),
    .y(_0007_)
  );
  al_nand2 _1176_ (
    .a(\DFF_161.D ),
    .b(_0534_),
    .y(_0008_)
  );
  al_aoi21ftf _1177_ (
    .a(\DFF_38.Q ),
    .b(_0535_),
    .c(_0008_),
    .y(_0009_)
  );
  al_nand3fft _1178_ (
    .a(\DFF_35.Q ),
    .b(_0531_),
    .c(_0552_),
    .y(_0010_)
  );
  al_nand2ft _1179_ (
    .a(\DFF_89.Q ),
    .b(_0537_),
    .y(_0011_)
  );
  al_nand3 _1180_ (
    .a(_0011_),
    .b(_0010_),
    .c(_0009_),
    .y(_0012_)
  );
  al_ao21ftf _1181_ (
    .a(_0529_),
    .b(_0012_),
    .c(_0007_),
    .y(n3135gat)
  );
  al_nand2ft _1182_ (
    .a(\DFF_79.Q ),
    .b(_0537_),
    .y(_0013_)
  );
  al_oai21ftf _1183_ (
    .a(_0542_),
    .b(_0534_),
    .c(\DFF_39.Q ),
    .y(_0014_)
  );
  al_ao21 _1184_ (
    .a(_0013_),
    .b(_0014_),
    .c(_0547_),
    .y(_0015_)
  );
  al_and2ft _1185_ (
    .a(\DFF_90.Q ),
    .b(_0537_),
    .y(_0016_)
  );
  al_nor2 _1186_ (
    .a(\DFF_36.Q ),
    .b(_0542_),
    .y(_0017_)
  );
  al_nand2 _1187_ (
    .a(\DFF_162.D ),
    .b(_0534_),
    .y(_0018_)
  );
  al_aoi21ftf _1188_ (
    .a(\DFF_39.Q ),
    .b(_0535_),
    .c(_0018_),
    .y(_0019_)
  );
  al_nand3fft _1189_ (
    .a(_0016_),
    .b(_0017_),
    .c(_0019_),
    .y(_0020_)
  );
  al_ao21ftf _1190_ (
    .a(_0529_),
    .b(_0020_),
    .c(_0015_),
    .y(n3134gat)
  );
  al_and2ft _1191_ (
    .a(\DFF_88.Q ),
    .b(_0537_),
    .y(_0021_)
  );
  al_nor2 _1192_ (
    .a(\DFF_34.Q ),
    .b(_0542_),
    .y(_0022_)
  );
  al_nand2 _1193_ (
    .a(_0207_),
    .b(_0534_),
    .y(_0023_)
  );
  al_aoi21ftf _1194_ (
    .a(\DFF_26.Q ),
    .b(_0535_),
    .c(_0023_),
    .y(_0024_)
  );
  al_nand3fft _1195_ (
    .a(_0021_),
    .b(_0022_),
    .c(_0024_),
    .y(_0025_)
  );
  al_nand3fft _1196_ (
    .a(\DFF_26.Q ),
    .b(_0531_),
    .c(_0552_),
    .y(_0026_)
  );
  al_nand2 _1197_ (
    .a(\DFF_156.D ),
    .b(_0534_),
    .y(_0027_)
  );
  al_aoi21ftf _1198_ (
    .a(\DFF_77.Q ),
    .b(_0537_),
    .c(_0027_),
    .y(_0028_)
  );
  al_ao21 _1199_ (
    .a(_0026_),
    .b(_0028_),
    .c(_0547_),
    .y(_0029_)
  );
  al_ao21ftf _1200_ (
    .a(_0529_),
    .b(_0025_),
    .c(_0029_),
    .y(n3133gat)
  );
  al_nand2ft _1201_ (
    .a(\DFF_49.Q ),
    .b(_0534_),
    .y(_0030_)
  );
  al_aoi21ftf _1202_ (
    .a(\DFF_84.Q ),
    .b(_0537_),
    .c(_0030_),
    .y(_0031_)
  );
  al_nand3fft _1203_ (
    .a(\DFF_29.Q ),
    .b(_0531_),
    .c(_0552_),
    .y(_0032_)
  );
  al_nand2ft _1204_ (
    .a(\DFF_23.Q ),
    .b(_0535_),
    .y(_0033_)
  );
  al_nand3 _1205_ (
    .a(_0032_),
    .b(_0033_),
    .c(_0031_),
    .y(_0034_)
  );
  al_nand2 _1206_ (
    .a(\DFF_157.D ),
    .b(_0534_),
    .y(_0035_)
  );
  al_nand3fft _1207_ (
    .a(\DFF_23.Q ),
    .b(_0531_),
    .c(_0552_),
    .y(_0036_)
  );
  al_aoi21ftf _1208_ (
    .a(\DFF_73.Q ),
    .b(_0537_),
    .c(_0036_),
    .y(_0037_)
  );
  al_ao21 _1209_ (
    .a(_0035_),
    .b(_0037_),
    .c(_0547_),
    .y(_0038_)
  );
  al_ao21ftf _1210_ (
    .a(_0529_),
    .b(_0034_),
    .c(_0038_),
    .y(n3132gat)
  );
  al_and2ft _1211_ (
    .a(\DFF_50.Q ),
    .b(_0534_),
    .y(_0039_)
  );
  al_and2ft _1212_ (
    .a(\DFF_85.Q ),
    .b(_0537_),
    .y(_0040_)
  );
  al_nand3fft _1213_ (
    .a(\DFF_30.Q ),
    .b(_0531_),
    .c(_0552_),
    .y(_0041_)
  );
  al_aoi21ftf _1214_ (
    .a(\DFF_24.Q ),
    .b(_0535_),
    .c(_0041_),
    .y(_0042_)
  );
  al_nand3fft _1215_ (
    .a(_0039_),
    .b(_0040_),
    .c(_0042_),
    .y(_0043_)
  );
  al_inv _1216_ (
    .a(\DFF_74.Q ),
    .y(_0044_)
  );
  al_nand2 _1217_ (
    .a(_0044_),
    .b(_0537_),
    .y(_0045_)
  );
  al_nand2 _1218_ (
    .a(\DFF_163.D ),
    .b(_0534_),
    .y(_0046_)
  );
  al_aoi21ftf _1219_ (
    .a(_0542_),
    .b(_0447_),
    .c(_0046_),
    .y(_0047_)
  );
  al_ao21 _1220_ (
    .a(_0045_),
    .b(_0047_),
    .c(_0547_),
    .y(_0048_)
  );
  al_ao21ftf _1221_ (
    .a(_0529_),
    .b(_0043_),
    .c(_0048_),
    .y(n3131gat)
  );
  al_nor2 _1222_ (
    .a(\DFF_28.Q ),
    .b(_0542_),
    .y(_0049_)
  );
  al_and2ft _1223_ (
    .a(\DFF_83.Q ),
    .b(_0537_),
    .y(_0050_)
  );
  al_nand2ft _1224_ (
    .a(\DFF_48.Q ),
    .b(_0534_),
    .y(_0051_)
  );
  al_aoi21ftf _1225_ (
    .a(\DFF_22.Q ),
    .b(_0535_),
    .c(_0051_),
    .y(_0052_)
  );
  al_nand3fft _1226_ (
    .a(_0049_),
    .b(_0050_),
    .c(_0052_),
    .y(_0053_)
  );
  al_nand3fft _1227_ (
    .a(\DFF_22.Q ),
    .b(_0531_),
    .c(_0552_),
    .y(_0054_)
  );
  al_nand2 _1228_ (
    .a(\DFF_165.D ),
    .b(_0534_),
    .y(_0055_)
  );
  al_aoi21ftf _1229_ (
    .a(\DFF_72.Q ),
    .b(_0537_),
    .c(_0055_),
    .y(_0056_)
  );
  al_ao21 _1230_ (
    .a(_0054_),
    .b(_0056_),
    .c(_0547_),
    .y(_0057_)
  );
  al_ao21ftf _1231_ (
    .a(_0529_),
    .b(_0053_),
    .c(_0057_),
    .y(n3130gat)
  );
  al_nand3 _1232_ (
    .a(_0537_),
    .b(_0183_),
    .c(_0182_),
    .y(_0058_)
  );
  al_nand2ft _1233_ (
    .a(_0532_),
    .b(_0533_),
    .y(_0059_)
  );
  al_or3fft _1234_ (
    .a(\DFF_33.Q ),
    .b(_0532_),
    .c(_0533_),
    .y(_0060_)
  );
  al_ao21ttf _1235_ (
    .a(_0060_),
    .b(_0059_),
    .c(_0531_),
    .y(_0061_)
  );
  al_nand2ft _1236_ (
    .a(\DFF_25.Q ),
    .b(_0535_),
    .y(_0062_)
  );
  al_nand3fft _1237_ (
    .a(\DFF_32.Q ),
    .b(_0531_),
    .c(_0552_),
    .y(_0063_)
  );
  al_aoi21ftf _1238_ (
    .a(\DFF_52.Q ),
    .b(_0534_),
    .c(_0063_),
    .y(_0064_)
  );
  al_and3 _1239_ (
    .a(_0062_),
    .b(_0061_),
    .c(_0064_),
    .y(_0065_)
  );
  al_ao21 _1240_ (
    .a(_0058_),
    .b(_0065_),
    .c(_0529_),
    .y(_0066_)
  );
  al_nand3fft _1241_ (
    .a(\DFF_25.Q ),
    .b(_0531_),
    .c(_0552_),
    .y(_0067_)
  );
  al_aoi21ftf _1242_ (
    .a(\DFF_45.Q ),
    .b(_0534_),
    .c(_0067_),
    .y(_0068_)
  );
  al_ao21ttf _1243_ (
    .a(_0537_),
    .b(n3116gat),
    .c(_0068_),
    .y(_0069_)
  );
  al_ao21ftf _1244_ (
    .a(_0547_),
    .b(_0069_),
    .c(_0066_),
    .y(n3129gat)
  );
  al_ao21 _1245_ (
    .a(_0058_),
    .b(_0065_),
    .c(_0544_),
    .y(_0070_)
  );
  al_nand2 _1246_ (
    .a(\DFF_99.D ),
    .b(_0070_),
    .y(n3125gat)
  );
  al_ao21ftf _1247_ (
    .a(_0544_),
    .b(_0540_),
    .c(\DFF_81.D ),
    .y(n3124gat)
  );
  al_ao21ftf _1248_ (
    .a(_0544_),
    .b(_0001_),
    .c(\DFF_91.D ),
    .y(n3123gat)
  );
  al_ao21ftf _1249_ (
    .a(_0544_),
    .b(_0012_),
    .c(\DFF_47.D ),
    .y(n3122gat)
  );
  al_ao21ftf _1250_ (
    .a(_0544_),
    .b(_0020_),
    .c(\DFF_57.D ),
    .y(n3121gat)
  );
  al_ao21ftf _1251_ (
    .a(_0544_),
    .b(_0025_),
    .c(\DFF_27.D ),
    .y(n3120gat)
  );
  al_ao21ftf _1252_ (
    .a(_0544_),
    .b(_0034_),
    .c(\DFF_37.D ),
    .y(n3119gat)
  );
  al_ao21ftf _1253_ (
    .a(_0544_),
    .b(_0043_),
    .c(\DFF_27.D ),
    .y(n3118gat)
  );
  al_ao21ftf _1254_ (
    .a(_0544_),
    .b(_0053_),
    .c(\DFF_9.D ),
    .y(n3117gat)
  );
  al_nand3 _1255_ (
    .a(\DFF_125.Q ),
    .b(\DFF_123.Q ),
    .c(\DFF_75.Q ),
    .y(n3114gat)
  );
  al_oai21ftt _1256_ (
    .a(_0327_),
    .b(_0328_),
    .c(\DFF_78.Q ),
    .y(n3113gat)
  );
  al_nand3 _1257_ (
    .a(\DFF_112.Q ),
    .b(\DFF_111.Q ),
    .c(\DFF_77.Q ),
    .y(n3111gat)
  );
  al_ao21ttf _1258_ (
    .a(_0111_),
    .b(_0343_),
    .c(\DFF_73.Q ),
    .y(n3110gat)
  );
  al_oai21ftf _1259_ (
    .a(_0115_),
    .b(_0116_),
    .c(_0044_),
    .y(n3109gat)
  );
  al_or3fft _1260_ (
    .a(\DFF_72.Q ),
    .b(_0112_),
    .c(_0113_),
    .y(n3108gat)
  );
  al_and3ftt _1261_ (
    .a(n3087gat),
    .b(_0360_),
    .c(_0398_),
    .y(_0071_)
  );
  al_or3fft _1262_ (
    .a(_0373_),
    .b(_0376_),
    .c(_0378_),
    .y(_0072_)
  );
  al_nand3ftt _1263_ (
    .a(_0071_),
    .b(_0339_),
    .c(_0072_),
    .y(n3105gat)
  );
  al_oa21ftf _1264_ (
    .a(n3094gat),
    .b(_0446_),
    .c(_0330_),
    .y(_0073_)
  );
  al_ao21ftf _1265_ (
    .a(_0445_),
    .b(_0359_),
    .c(_0073_),
    .y(n3104gat)
  );
  al_inv _1266_ (
    .a(\DFF_19.Q ),
    .y(\DFF_20.D )
  );
  al_nand3ftt _1267_ (
    .a(_0283_),
    .b(_0282_),
    .c(_0288_),
    .y(\DFF_116.D )
  );
  al_nand2ft _1268_ (
    .a(_0370_),
    .b(_0358_),
    .y(_0074_)
  );
  al_ao21ftf _1269_ (
    .a(_0365_),
    .b(_0527_),
    .c(_0074_),
    .y(\DFF_139.D )
  );
  al_oai21ftt _1270_ (
    .a(\DFF_123.Q ),
    .b(\DFF_125.Q ),
    .c(\DFF_148.Q ),
    .y(_0075_)
  );
  al_or3ftt _1271_ (
    .a(\DFF_123.Q ),
    .b(\DFF_125.Q ),
    .c(\DFF_148.Q ),
    .y(_0076_)
  );
  al_nand3 _1272_ (
    .a(_0075_),
    .b(_0076_),
    .c(\DFF_96.D ),
    .y(\DFF_95.D )
  );
  al_or3ftt _1273_ (
    .a(\DFF_105.Q ),
    .b(\DFF_108.Q ),
    .c(\DFF_106.Q ),
    .y(_0077_)
  );
  al_nand3 _1274_ (
    .a(\DFF_154.Q ),
    .b(_0296_),
    .c(_0077_),
    .y(_0078_)
  );
  al_ao21 _1275_ (
    .a(_0296_),
    .b(_0077_),
    .c(\DFF_154.Q ),
    .y(_0079_)
  );
  al_nand3 _1276_ (
    .a(_0078_),
    .b(_0079_),
    .c(\DFF_63.D ),
    .y(\DFF_100.D )
  );
  al_oai21ftf _1277_ (
    .a(\DFF_114.Q ),
    .b(\DFF_110.Q ),
    .c(\DFF_111.Q ),
    .y(_0080_)
  );
  al_nand3fft _1278_ (
    .a(\DFF_112.Q ),
    .b(\DFF_155.Q ),
    .c(_0080_),
    .y(_0081_)
  );
  al_ao21ftf _1279_ (
    .a(\DFF_112.Q ),
    .b(_0080_),
    .c(\DFF_155.Q ),
    .y(_0082_)
  );
  al_nand3 _1280_ (
    .a(_0081_),
    .b(_0082_),
    .c(\DFF_61.D ),
    .y(\DFF_93.D )
  );
  al_nand3fft _1281_ (
    .a(\DFF_118.D ),
    .b(\DFF_176.Q ),
    .c(_0516_),
    .y(_0083_)
  );
  al_ao21ttf _1282_ (
    .a(_0384_),
    .b(_0517_),
    .c(_0083_),
    .y(_0084_)
  );
  al_or2 _1283_ (
    .a(\DFF_177.Q ),
    .b(\DFF_135.Q ),
    .y(_0085_)
  );
  al_ao21 _1284_ (
    .a(\DFF_118.D ),
    .b(_0284_),
    .c(_0085_),
    .y(_0086_)
  );
  al_ao21ftf _1285_ (
    .a(\DFF_178.Q ),
    .b(\DFF_177.Q ),
    .c(_0086_),
    .y(_0087_)
  );
  al_nor2 _1286_ (
    .a(\DFF_117.Q ),
    .b(\DFF_175.Q ),
    .y(_0088_)
  );
  al_ao21 _1287_ (
    .a(_0088_),
    .b(\DFF_119.D ),
    .c(_0087_),
    .y(_0089_)
  );
  al_and2 _1288_ (
    .a(n3097gat),
    .b(\DFF_21.Q ),
    .y(_0090_)
  );
  al_ao21 _1289_ (
    .a(_0307_),
    .b(_0090_),
    .c(\DFF_20.D ),
    .y(_0091_)
  );
  al_and3fft _1290_ (
    .a(\DFF_131.Q ),
    .b(n3098gat),
    .c(\DFF_132.Q ),
    .y(_0092_)
  );
  al_and3fft _1291_ (
    .a(\DFF_135.Q ),
    .b(_0098_),
    .c(\DFF_176.Q ),
    .y(_0093_)
  );
  al_ao21 _1292_ (
    .a(_0092_),
    .b(_0091_),
    .c(_0093_),
    .y(_0094_)
  );
  al_aoi21 _1293_ (
    .a(_0098_),
    .b(_0089_),
    .c(_0094_),
    .y(_0095_)
  );
  al_ao21ftf _1294_ (
    .a(\DFF_134.Q ),
    .b(_0084_),
    .c(_0095_),
    .y(n3140gat)
  );
  al_ao21ftf _1295_ (
    .a(\DFF_134.Q ),
    .b(_0084_),
    .c(_0095_),
    .y(n3139gat)
  );
  al_dffl _1296_ (
    .clk(CK),
    .d(\DFF_9.D ),
    .q(\DFF_9.Q )
  );
  al_dffl _1297_ (
    .clk(CK),
    .d(\DFF_16.D ),
    .q(\DFF_16.Q )
  );
  al_dffl _1298_ (
    .clk(CK),
    .d(\DFF_17.D ),
    .q(\DFF_17.Q )
  );
  al_dffl _1299_ (
    .clk(CK),
    .d(\DFF_19.D ),
    .q(\DFF_19.Q )
  );
  al_dffl _1300_ (
    .clk(CK),
    .d(\DFF_20.D ),
    .q(\DFF_20.Q )
  );
  al_dffl _1301_ (
    .clk(CK),
    .d(\DFF_21.D ),
    .q(\DFF_21.Q )
  );
  al_dffl _1302_ (
    .clk(CK),
    .d(n3065gat),
    .q(\DFF_22.Q )
  );
  al_dffl _1303_ (
    .clk(CK),
    .d(n3067gat),
    .q(\DFF_23.Q )
  );
  al_dffl _1304_ (
    .clk(CK),
    .d(n3066gat),
    .q(\DFF_24.Q )
  );
  al_dffl _1305_ (
    .clk(CK),
    .d(n3073gat),
    .q(\DFF_25.Q )
  );
  al_dffl _1306_ (
    .clk(CK),
    .d(n3068gat),
    .q(\DFF_26.Q )
  );
  al_dffl _1307_ (
    .clk(CK),
    .d(\DFF_27.D ),
    .q(\DFF_27.Q )
  );
  al_dffl _1308_ (
    .clk(CK),
    .d(\DFF_28.D ),
    .q(\DFF_28.Q )
  );
  al_dffl _1309_ (
    .clk(CK),
    .d(\DFF_29.D ),
    .q(\DFF_29.Q )
  );
  al_dffl _1310_ (
    .clk(CK),
    .d(\DFF_30.D ),
    .q(\DFF_30.Q )
  );
  al_dffl _1311_ (
    .clk(CK),
    .d(\DFF_31.D ),
    .q(\DFF_31.Q )
  );
  al_dffl _1312_ (
    .clk(CK),
    .d(\DFF_32.D ),
    .q(\DFF_32.Q )
  );
  al_dffl _1313_ (
    .clk(CK),
    .d(\DFF_33.D ),
    .q(\DFF_33.Q )
  );
  al_dffl _1314_ (
    .clk(CK),
    .d(\DFF_34.D ),
    .q(\DFF_34.Q )
  );
  al_dffl _1315_ (
    .clk(CK),
    .d(\DFF_35.D ),
    .q(\DFF_35.Q )
  );
  al_dffl _1316_ (
    .clk(CK),
    .d(\DFF_36.D ),
    .q(\DFF_36.Q )
  );
  al_dffl _1317_ (
    .clk(CK),
    .d(\DFF_37.D ),
    .q(\DFF_37.Q )
  );
  al_dffl _1318_ (
    .clk(CK),
    .d(n3070gat),
    .q(\DFF_38.Q )
  );
  al_dffl _1319_ (
    .clk(CK),
    .d(n3069gat),
    .q(\DFF_39.Q )
  );
  al_dffl _1320_ (
    .clk(CK),
    .d(n3071gat),
    .q(\DFF_40.Q )
  );
  al_dffl _1321_ (
    .clk(CK),
    .d(n3072gat),
    .q(\DFF_41.Q )
  );
  al_dffl _1322_ (
    .clk(CK),
    .d(\DFF_42.D ),
    .q(\DFF_42.Q )
  );
  al_dffl _1323_ (
    .clk(CK),
    .d(\DFF_43.D ),
    .q(\DFF_43.Q )
  );
  al_dffl _1324_ (
    .clk(CK),
    .d(\DFF_44.D ),
    .q(\DFF_44.Q )
  );
  al_dffl _1325_ (
    .clk(CK),
    .d(\DFF_45.D ),
    .q(\DFF_45.Q )
  );
  al_dffl _1326_ (
    .clk(CK),
    .d(\DFF_46.D ),
    .q(\DFF_46.Q )
  );
  al_dffl _1327_ (
    .clk(CK),
    .d(\DFF_47.D ),
    .q(\DFF_47.Q )
  );
  al_dffl _1328_ (
    .clk(CK),
    .d(\DFF_48.D ),
    .q(\DFF_48.Q )
  );
  al_dffl _1329_ (
    .clk(CK),
    .d(\DFF_49.D ),
    .q(\DFF_49.Q )
  );
  al_dffl _1330_ (
    .clk(CK),
    .d(\DFF_50.D ),
    .q(\DFF_50.Q )
  );
  al_dffl _1331_ (
    .clk(CK),
    .d(\DFF_51.D ),
    .q(\DFF_51.Q )
  );
  al_dffl _1332_ (
    .clk(CK),
    .d(\DFF_52.D ),
    .q(\DFF_52.Q )
  );
  al_dffl _1333_ (
    .clk(CK),
    .d(\DFF_53.D ),
    .q(\DFF_53.Q )
  );
  al_dffl _1334_ (
    .clk(CK),
    .d(\DFF_54.D ),
    .q(\DFF_54.Q )
  );
  al_dffl _1335_ (
    .clk(CK),
    .d(\DFF_55.D ),
    .q(\DFF_55.Q )
  );
  al_dffl _1336_ (
    .clk(CK),
    .d(\DFF_56.D ),
    .q(\DFF_56.Q )
  );
  al_dffl _1337_ (
    .clk(CK),
    .d(\DFF_57.D ),
    .q(\DFF_57.Q )
  );
  al_dffl _1338_ (
    .clk(CK),
    .d(\DFF_58.D ),
    .q(\DFF_58.Q )
  );
  al_dffl _1339_ (
    .clk(CK),
    .d(\DFF_59.D ),
    .q(\DFF_59.Q )
  );
  al_dffl _1340_ (
    .clk(CK),
    .d(\DFF_60.D ),
    .q(\DFF_60.Q )
  );
  al_dffl _1341_ (
    .clk(CK),
    .d(\DFF_61.D ),
    .q(\DFF_61.Q )
  );
  al_dffl _1342_ (
    .clk(CK),
    .d(\DFF_62.D ),
    .q(\DFF_62.Q )
  );
  al_dffl _1343_ (
    .clk(CK),
    .d(\DFF_63.D ),
    .q(\DFF_63.Q )
  );
  al_dffl _1344_ (
    .clk(CK),
    .d(\DFF_64.D ),
    .q(\DFF_64.Q )
  );
  al_dffl _1345_ (
    .clk(CK),
    .d(\DFF_65.D ),
    .q(\DFF_65.Q )
  );
  al_dffl _1346_ (
    .clk(CK),
    .d(\DFF_66.D ),
    .q(\DFF_66.Q )
  );
  al_dffl _1347_ (
    .clk(CK),
    .d(\DFF_67.D ),
    .q(\DFF_67.Q )
  );
  al_dffl _1348_ (
    .clk(CK),
    .d(\DFF_68.D ),
    .q(\DFF_68.Q )
  );
  al_dffl _1349_ (
    .clk(CK),
    .d(\DFF_69.D ),
    .q(\DFF_69.Q )
  );
  al_dffl _1350_ (
    .clk(CK),
    .d(\DFF_70.D ),
    .q(\DFF_70.Q )
  );
  al_dffl _1351_ (
    .clk(CK),
    .d(\DFF_71.D ),
    .q(\DFF_71.Q )
  );
  al_dffl _1352_ (
    .clk(CK),
    .d(\DFF_72.D ),
    .q(\DFF_72.Q )
  );
  al_dffl _1353_ (
    .clk(CK),
    .d(\DFF_73.D ),
    .q(\DFF_73.Q )
  );
  al_dffl _1354_ (
    .clk(CK),
    .d(\DFF_74.D ),
    .q(\DFF_74.Q )
  );
  al_dffl _1355_ (
    .clk(CK),
    .d(\DFF_75.D ),
    .q(\DFF_75.Q )
  );
  al_dffl _1356_ (
    .clk(CK),
    .d(\DFF_76.D ),
    .q(\DFF_76.Q )
  );
  al_dffl _1357_ (
    .clk(CK),
    .d(\DFF_77.D ),
    .q(\DFF_77.Q )
  );
  al_dffl _1358_ (
    .clk(CK),
    .d(\DFF_78.D ),
    .q(\DFF_78.Q )
  );
  al_dffl _1359_ (
    .clk(CK),
    .d(\DFF_79.D ),
    .q(\DFF_79.Q )
  );
  al_dffl _1360_ (
    .clk(CK),
    .d(\DFF_80.D ),
    .q(\DFF_80.Q )
  );
  al_dffl _1361_ (
    .clk(CK),
    .d(\DFF_81.D ),
    .q(\DFF_81.Q )
  );
  al_dffl _1362_ (
    .clk(CK),
    .d(\DFF_82.D ),
    .q(\DFF_82.Q )
  );
  al_dffl _1363_ (
    .clk(CK),
    .d(\DFF_83.D ),
    .q(\DFF_83.Q )
  );
  al_dffl _1364_ (
    .clk(CK),
    .d(\DFF_84.D ),
    .q(\DFF_84.Q )
  );
  al_dffl _1365_ (
    .clk(CK),
    .d(\DFF_85.D ),
    .q(\DFF_85.Q )
  );
  al_dffl _1366_ (
    .clk(CK),
    .d(\DFF_86.D ),
    .q(\DFF_86.Q )
  );
  al_dffl _1367_ (
    .clk(CK),
    .d(\DFF_87.D ),
    .q(\DFF_87.Q )
  );
  al_dffl _1368_ (
    .clk(CK),
    .d(\DFF_88.D ),
    .q(\DFF_88.Q )
  );
  al_dffl _1369_ (
    .clk(CK),
    .d(\DFF_89.D ),
    .q(\DFF_89.Q )
  );
  al_dffl _1370_ (
    .clk(CK),
    .d(\DFF_90.D ),
    .q(\DFF_90.Q )
  );
  al_dffl _1371_ (
    .clk(CK),
    .d(\DFF_91.D ),
    .q(\DFF_91.Q )
  );
  al_dffl _1372_ (
    .clk(CK),
    .d(\DFF_92.D ),
    .q(\DFF_92.Q )
  );
  al_dffl _1373_ (
    .clk(CK),
    .d(\DFF_93.D ),
    .q(\DFF_93.Q )
  );
  al_dffl _1374_ (
    .clk(CK),
    .d(\DFF_94.D ),
    .q(\DFF_94.Q )
  );
  al_dffl _1375_ (
    .clk(CK),
    .d(\DFF_95.D ),
    .q(\DFF_95.Q )
  );
  al_dffl _1376_ (
    .clk(CK),
    .d(\DFF_96.D ),
    .q(\DFF_96.Q )
  );
  al_dffl _1377_ (
    .clk(CK),
    .d(\DFF_97.D ),
    .q(\DFF_97.Q )
  );
  al_dffl _1378_ (
    .clk(CK),
    .d(\DFF_98.D ),
    .q(\DFF_98.Q )
  );
  al_dffl _1379_ (
    .clk(CK),
    .d(\DFF_99.D ),
    .q(\DFF_99.Q )
  );
  al_dffl _1380_ (
    .clk(CK),
    .d(\DFF_100.D ),
    .q(\DFF_100.Q )
  );
  al_dffl _1381_ (
    .clk(CK),
    .d(\DFF_101.D ),
    .q(\DFF_101.Q )
  );
  al_dffl _1382_ (
    .clk(CK),
    .d(\DFF_102.D ),
    .q(\DFF_102.Q )
  );
  al_dffl _1383_ (
    .clk(CK),
    .d(\DFF_103.D ),
    .q(\DFF_103.Q )
  );
  al_dffl _1384_ (
    .clk(CK),
    .d(\DFF_104.D ),
    .q(\DFF_104.Q )
  );
  al_dffl _1385_ (
    .clk(CK),
    .d(\DFF_105.D ),
    .q(\DFF_105.Q )
  );
  al_dffl _1386_ (
    .clk(CK),
    .d(\DFF_106.D ),
    .q(\DFF_106.Q )
  );
  al_dffl _1387_ (
    .clk(CK),
    .d(\DFF_107.D ),
    .q(\DFF_107.Q )
  );
  al_dffl _1388_ (
    .clk(CK),
    .d(\DFF_108.D ),
    .q(\DFF_108.Q )
  );
  al_dffl _1389_ (
    .clk(CK),
    .d(\DFF_109.D ),
    .q(\DFF_109.Q )
  );
  al_dffl _1390_ (
    .clk(CK),
    .d(\DFF_110.D ),
    .q(\DFF_110.Q )
  );
  al_dffl _1391_ (
    .clk(CK),
    .d(\DFF_111.D ),
    .q(\DFF_111.Q )
  );
  al_dffl _1392_ (
    .clk(CK),
    .d(\DFF_112.D ),
    .q(\DFF_112.Q )
  );
  al_dffl _1393_ (
    .clk(CK),
    .d(\DFF_113.D ),
    .q(\DFF_113.Q )
  );
  al_dffl _1394_ (
    .clk(CK),
    .d(\DFF_114.D ),
    .q(\DFF_114.Q )
  );
  al_dffl _1395_ (
    .clk(CK),
    .d(\DFF_115.D ),
    .q(\DFF_115.Q )
  );
  al_dffl _1396_ (
    .clk(CK),
    .d(\DFF_116.D ),
    .q(\DFF_116.Q )
  );
  al_dffl _1397_ (
    .clk(CK),
    .d(\DFF_117.D ),
    .q(\DFF_117.Q )
  );
  al_dffl _1398_ (
    .clk(CK),
    .d(\DFF_118.D ),
    .q(\DFF_118.Q )
  );
  al_dffl _1399_ (
    .clk(CK),
    .d(\DFF_119.D ),
    .q(\DFF_119.Q )
  );
  al_dffl _1400_ (
    .clk(CK),
    .d(\DFF_120.D ),
    .q(\DFF_120.Q )
  );
  al_dffl _1401_ (
    .clk(CK),
    .d(\DFF_121.D ),
    .q(\DFF_121.Q )
  );
  al_dffl _1402_ (
    .clk(CK),
    .d(\DFF_122.D ),
    .q(\DFF_122.Q )
  );
  al_dffl _1403_ (
    .clk(CK),
    .d(\DFF_123.D ),
    .q(\DFF_123.Q )
  );
  al_dffl _1404_ (
    .clk(CK),
    .d(\DFF_124.D ),
    .q(\DFF_124.Q )
  );
  al_dffl _1405_ (
    .clk(CK),
    .d(\DFF_125.D ),
    .q(\DFF_125.Q )
  );
  al_dffl _1406_ (
    .clk(CK),
    .d(\DFF_126.D ),
    .q(\DFF_126.Q )
  );
  al_dffl _1407_ (
    .clk(CK),
    .d(\DFF_127.D ),
    .q(\DFF_127.Q )
  );
  al_dffl _1408_ (
    .clk(CK),
    .d(\DFF_128.D ),
    .q(\DFF_128.Q )
  );
  al_dffl _1409_ (
    .clk(CK),
    .d(\DFF_129.D ),
    .q(\DFF_129.Q )
  );
  al_dffl _1410_ (
    .clk(CK),
    .d(\DFF_130.D ),
    .q(\DFF_130.Q )
  );
  al_dffl _1411_ (
    .clk(CK),
    .d(\DFF_131.D ),
    .q(\DFF_131.Q )
  );
  al_dffl _1412_ (
    .clk(CK),
    .d(\DFF_132.D ),
    .q(\DFF_132.Q )
  );
  al_dffl _1413_ (
    .clk(CK),
    .d(\DFF_133.D ),
    .q(\DFF_133.Q )
  );
  al_dffl _1414_ (
    .clk(CK),
    .d(\DFF_134.D ),
    .q(\DFF_134.Q )
  );
  al_dffl _1415_ (
    .clk(CK),
    .d(\DFF_135.D ),
    .q(\DFF_135.Q )
  );
  al_dffl _1416_ (
    .clk(CK),
    .d(\DFF_139.D ),
    .q(\DFF_139.Q )
  );
  al_dffl _1417_ (
    .clk(CK),
    .d(\DFF_140.D ),
    .q(\DFF_140.Q )
  );
  al_dffl _1418_ (
    .clk(CK),
    .d(\DFF_141.D ),
    .q(\DFF_141.Q )
  );
  al_dffl _1419_ (
    .clk(CK),
    .d(\DFF_142.D ),
    .q(\DFF_142.Q )
  );
  al_dffl _1420_ (
    .clk(CK),
    .d(\DFF_143.D ),
    .q(\DFF_143.Q )
  );
  al_dffl _1421_ (
    .clk(CK),
    .d(\DFF_144.D ),
    .q(\DFF_144.Q )
  );
  al_dffl _1422_ (
    .clk(CK),
    .d(\DFF_145.D ),
    .q(\DFF_145.Q )
  );
  al_dffl _1423_ (
    .clk(CK),
    .d(\DFF_146.D ),
    .q(\DFF_146.Q )
  );
  al_dffl _1424_ (
    .clk(CK),
    .d(\DFF_147.D ),
    .q(\DFF_147.Q )
  );
  al_dffl _1425_ (
    .clk(CK),
    .d(\DFF_148.D ),
    .q(\DFF_148.Q )
  );
  al_dffl _1426_ (
    .clk(CK),
    .d(\DFF_149.D ),
    .q(\DFF_149.Q )
  );
  al_dffl _1427_ (
    .clk(CK),
    .d(\DFF_150.D ),
    .q(\DFF_150.Q )
  );
  al_dffl _1428_ (
    .clk(CK),
    .d(\DFF_151.D ),
    .q(\DFF_151.Q )
  );
  al_dffl _1429_ (
    .clk(CK),
    .d(\DFF_152.D ),
    .q(\DFF_152.Q )
  );
  al_dffl _1430_ (
    .clk(CK),
    .d(\DFF_153.D ),
    .q(\DFF_153.Q )
  );
  al_dffl _1431_ (
    .clk(CK),
    .d(\DFF_154.D ),
    .q(\DFF_154.Q )
  );
  al_dffl _1432_ (
    .clk(CK),
    .d(\DFF_155.D ),
    .q(\DFF_155.Q )
  );
  al_dffl _1433_ (
    .clk(CK),
    .d(\DFF_156.D ),
    .q(\DFF_156.Q )
  );
  al_dffl _1434_ (
    .clk(CK),
    .d(\DFF_157.D ),
    .q(\DFF_157.Q )
  );
  al_dffl _1435_ (
    .clk(CK),
    .d(\DFF_158.D ),
    .q(\DFF_158.Q )
  );
  al_dffl _1436_ (
    .clk(CK),
    .d(\DFF_159.D ),
    .q(\DFF_159.Q )
  );
  al_dffl _1437_ (
    .clk(CK),
    .d(\DFF_160.D ),
    .q(\DFF_160.Q )
  );
  al_dffl _1438_ (
    .clk(CK),
    .d(\DFF_161.D ),
    .q(\DFF_161.Q )
  );
  al_dffl _1439_ (
    .clk(CK),
    .d(\DFF_162.D ),
    .q(\DFF_162.Q )
  );
  al_dffl _1440_ (
    .clk(CK),
    .d(\DFF_163.D ),
    .q(\DFF_163.Q )
  );
  al_dffl _1441_ (
    .clk(CK),
    .d(\DFF_164.D ),
    .q(\DFF_164.Q )
  );
  al_dffl _1442_ (
    .clk(CK),
    .d(\DFF_165.D ),
    .q(\DFF_165.Q )
  );
  al_dffl _1443_ (
    .clk(CK),
    .d(\DFF_166.D ),
    .q(\DFF_166.Q )
  );
  al_dffl _1444_ (
    .clk(CK),
    .d(\DFF_167.D ),
    .q(\DFF_167.Q )
  );
  al_dffl _1445_ (
    .clk(CK),
    .d(\DFF_168.D ),
    .q(\DFF_168.Q )
  );
  al_dffl _1446_ (
    .clk(CK),
    .d(\DFF_169.D ),
    .q(\DFF_169.Q )
  );
  al_dffl _1447_ (
    .clk(CK),
    .d(\DFF_170.D ),
    .q(\DFF_170.Q )
  );
  al_dffl _1448_ (
    .clk(CK),
    .d(\DFF_171.D ),
    .q(\DFF_171.Q )
  );
  al_dffl _1449_ (
    .clk(CK),
    .d(\DFF_172.D ),
    .q(\DFF_172.Q )
  );
  al_dffl _1450_ (
    .clk(CK),
    .d(\DFF_173.D ),
    .q(\DFF_173.Q )
  );
  al_dffl _1451_ (
    .clk(CK),
    .d(\DFF_174.D ),
    .q(\DFF_174.Q )
  );
  al_dffl _1452_ (
    .clk(CK),
    .d(\DFF_175.D ),
    .q(\DFF_175.Q )
  );
  al_dffl _1453_ (
    .clk(CK),
    .d(\DFF_176.D ),
    .q(\DFF_176.Q )
  );
  al_dffl _1454_ (
    .clk(CK),
    .d(\DFF_177.D ),
    .q(\DFF_177.Q )
  );
  al_dffl _1455_ (
    .clk(CK),
    .d(\DFF_178.D ),
    .q(\DFF_178.Q )
  );
  assign \DFF_0.CK  = CK;
  assign \DFF_0.D  = \DFF_33.D ;
  assign \DFF_0.Q  = \DFF_33.Q ;
  assign \DFF_1.CK  = CK;
  assign \DFF_1.D  = n3069gat;
  assign \DFF_1.Q  = \DFF_39.Q ;
  assign \DFF_10.CK  = CK;
  assign \DFF_10.D  = n3065gat;
  assign \DFF_10.Q  = \DFF_22.Q ;
  assign \DFF_100.CK  = CK;
  assign \DFF_101.CK  = CK;
  assign \DFF_102.CK  = CK;
  assign \DFF_103.CK  = CK;
  assign \DFF_104.CK  = CK;
  assign \DFF_105.CK  = CK;
  assign \DFF_106.CK  = CK;
  assign \DFF_107.CK  = CK;
  assign \DFF_108.CK  = CK;
  assign \DFF_109.CK  = CK;
  assign \DFF_11.CK  = CK;
  assign \DFF_11.D  = n3067gat;
  assign \DFF_11.Q  = \DFF_23.Q ;
  assign \DFF_110.CK  = CK;
  assign \DFF_111.CK  = CK;
  assign \DFF_112.CK  = CK;
  assign \DFF_113.CK  = CK;
  assign \DFF_114.CK  = CK;
  assign \DFF_115.CK  = CK;
  assign \DFF_116.CK  = CK;
  assign \DFF_117.CK  = CK;
  assign \DFF_118.CK  = CK;
  assign \DFF_119.CK  = CK;
  assign \DFF_12.CK  = CK;
  assign \DFF_12.D  = n3066gat;
  assign \DFF_12.Q  = \DFF_24.Q ;
  assign \DFF_120.CK  = CK;
  assign \DFF_121.CK  = CK;
  assign \DFF_122.CK  = CK;
  assign \DFF_123.CK  = CK;
  assign \DFF_124.CK  = CK;
  assign \DFF_125.CK  = CK;
  assign \DFF_126.CK  = CK;
  assign \DFF_127.CK  = CK;
  assign \DFF_128.CK  = CK;
  assign \DFF_129.CK  = CK;
  assign \DFF_13.CK  = CK;
  assign \DFF_13.D  = n3073gat;
  assign \DFF_13.Q  = \DFF_25.Q ;
  assign \DFF_130.CK  = CK;
  assign \DFF_131.CK  = CK;
  assign \DFF_132.CK  = CK;
  assign \DFF_133.CK  = CK;
  assign \DFF_134.CK  = CK;
  assign \DFF_135.CK  = CK;
  assign \DFF_136.CK  = CK;
  assign \DFF_137.CK  = CK;
  assign \DFF_138.CK  = CK;
  assign \DFF_139.CK  = CK;
  assign \DFF_14.CK  = CK;
  assign \DFF_14.D  = n3068gat;
  assign \DFF_14.Q  = \DFF_26.Q ;
  assign \DFF_140.CK  = CK;
  assign \DFF_141.CK  = CK;
  assign \DFF_142.CK  = CK;
  assign \DFF_143.CK  = CK;
  assign \DFF_144.CK  = CK;
  assign \DFF_145.CK  = CK;
  assign \DFF_146.CK  = CK;
  assign \DFF_147.CK  = CK;
  assign \DFF_148.CK  = CK;
  assign \DFF_149.CK  = CK;
  assign \DFF_15.CK  = CK;
  assign \DFF_15.D  = \DFF_27.D ;
  assign \DFF_15.Q  = \DFF_27.Q ;
  assign \DFF_150.CK  = CK;
  assign \DFF_151.CK  = CK;
  assign \DFF_152.CK  = CK;
  assign \DFF_153.CK  = CK;
  assign \DFF_154.CK  = CK;
  assign \DFF_155.CK  = CK;
  assign \DFF_156.CK  = CK;
  assign \DFF_157.CK  = CK;
  assign \DFF_158.CK  = CK;
  assign \DFF_159.CK  = CK;
  assign \DFF_16.CK  = CK;
  assign \DFF_160.CK  = CK;
  assign \DFF_161.CK  = CK;
  assign \DFF_162.CK  = CK;
  assign \DFF_163.CK  = CK;
  assign \DFF_164.CK  = CK;
  assign \DFF_165.CK  = CK;
  assign \DFF_166.CK  = CK;
  assign \DFF_167.CK  = CK;
  assign \DFF_168.CK  = CK;
  assign \DFF_169.CK  = CK;
  assign \DFF_17.CK  = CK;
  assign \DFF_170.CK  = CK;
  assign \DFF_171.CK  = CK;
  assign \DFF_172.CK  = CK;
  assign \DFF_173.CK  = CK;
  assign \DFF_174.CK  = CK;
  assign \DFF_175.CK  = CK;
  assign \DFF_176.CK  = CK;
  assign \DFF_177.CK  = CK;
  assign \DFF_178.CK  = CK;
  assign \DFF_18.CK  = CK;
  assign \DFF_18.D  = \DFF_19.D ;
  assign \DFF_18.Q  = \DFF_19.Q ;
  assign \DFF_19.CK  = CK;
  assign \DFF_2.CK  = CK;
  assign \DFF_2.D  = n3070gat;
  assign \DFF_2.Q  = \DFF_38.Q ;
  assign \DFF_20.CK  = CK;
  assign \DFF_21.CK  = CK;
  assign \DFF_22.CK  = CK;
  assign \DFF_22.D  = n3065gat;
  assign \DFF_23.CK  = CK;
  assign \DFF_23.D  = n3067gat;
  assign \DFF_24.CK  = CK;
  assign \DFF_24.D  = n3066gat;
  assign \DFF_25.CK  = CK;
  assign \DFF_25.D  = n3073gat;
  assign \DFF_26.CK  = CK;
  assign \DFF_26.D  = n3068gat;
  assign \DFF_27.CK  = CK;
  assign \DFF_28.CK  = CK;
  assign \DFF_29.CK  = CK;
  assign \DFF_3.CK  = CK;
  assign \DFF_3.D  = n3072gat;
  assign \DFF_3.Q  = \DFF_41.Q ;
  assign \DFF_30.CK  = CK;
  assign \DFF_31.CK  = CK;
  assign \DFF_32.CK  = CK;
  assign \DFF_33.CK  = CK;
  assign \DFF_34.CK  = CK;
  assign \DFF_35.CK  = CK;
  assign \DFF_36.CK  = CK;
  assign \DFF_37.CK  = CK;
  assign \DFF_38.CK  = CK;
  assign \DFF_38.D  = n3070gat;
  assign \DFF_39.CK  = CK;
  assign \DFF_39.D  = n3069gat;
  assign \DFF_4.CK  = CK;
  assign \DFF_4.D  = n3071gat;
  assign \DFF_4.Q  = \DFF_40.Q ;
  assign \DFF_40.CK  = CK;
  assign \DFF_40.D  = n3071gat;
  assign \DFF_41.CK  = CK;
  assign \DFF_41.D  = n3072gat;
  assign \DFF_42.CK  = CK;
  assign \DFF_43.CK  = CK;
  assign \DFF_44.CK  = CK;
  assign \DFF_45.CK  = CK;
  assign \DFF_46.CK  = CK;
  assign \DFF_47.CK  = CK;
  assign \DFF_48.CK  = CK;
  assign \DFF_49.CK  = CK;
  assign \DFF_5.CK  = CK;
  assign \DFF_5.D  = n3069gat;
  assign \DFF_5.Q  = \DFF_39.Q ;
  assign \DFF_50.CK  = CK;
  assign \DFF_51.CK  = CK;
  assign \DFF_52.CK  = CK;
  assign \DFF_53.CK  = CK;
  assign \DFF_54.CK  = CK;
  assign \DFF_55.CK  = CK;
  assign \DFF_56.CK  = CK;
  assign \DFF_57.CK  = CK;
  assign \DFF_58.CK  = CK;
  assign \DFF_59.CK  = CK;
  assign \DFF_6.CK  = CK;
  assign \DFF_6.D  = n3070gat;
  assign \DFF_6.Q  = \DFF_38.Q ;
  assign \DFF_60.CK  = CK;
  assign \DFF_61.CK  = CK;
  assign \DFF_62.CK  = CK;
  assign \DFF_63.CK  = CK;
  assign \DFF_64.CK  = CK;
  assign \DFF_65.CK  = CK;
  assign \DFF_66.CK  = CK;
  assign \DFF_67.CK  = CK;
  assign \DFF_68.CK  = CK;
  assign \DFF_69.CK  = CK;
  assign \DFF_7.CK  = CK;
  assign \DFF_7.D  = n3072gat;
  assign \DFF_7.Q  = \DFF_41.Q ;
  assign \DFF_70.CK  = CK;
  assign \DFF_71.CK  = CK;
  assign \DFF_72.CK  = CK;
  assign \DFF_73.CK  = CK;
  assign \DFF_74.CK  = CK;
  assign \DFF_75.CK  = CK;
  assign \DFF_76.CK  = CK;
  assign \DFF_77.CK  = CK;
  assign \DFF_78.CK  = CK;
  assign \DFF_79.CK  = CK;
  assign \DFF_8.CK  = CK;
  assign \DFF_8.D  = n3071gat;
  assign \DFF_8.Q  = \DFF_40.Q ;
  assign \DFF_80.CK  = CK;
  assign \DFF_81.CK  = CK;
  assign \DFF_82.CK  = CK;
  assign \DFF_83.CK  = CK;
  assign \DFF_84.CK  = CK;
  assign \DFF_85.CK  = CK;
  assign \DFF_86.CK  = CK;
  assign \DFF_87.CK  = CK;
  assign \DFF_88.CK  = CK;
  assign \DFF_89.CK  = CK;
  assign \DFF_9.CK  = CK;
  assign \DFF_90.CK  = CK;
  assign \DFF_91.CK  = CK;
  assign \DFF_92.CK  = CK;
  assign \DFF_93.CK  = CK;
  assign \DFF_94.CK  = CK;
  assign \DFF_95.CK  = CK;
  assign \DFF_96.CK  = CK;
  assign \DFF_97.CK  = CK;
  assign \DFF_98.CK  = CK;
  assign \DFF_99.CK  = CK;
  assign II1007 = \DFF_35.Q ;
  assign II1011 = \DFF_36.Q ;
  assign II1016 = \DFF_34.Q ;
  assign II1067 = \DFF_38.Q ;
  assign II1079 = \DFF_39.Q ;
  assign II1103 = \DFF_40.Q ;
  assign II1115 = \DFF_41.Q ;
  assign II1138 = \DFF_165.D ;
  assign II1141 = \DFF_165.D ;
  assign II1152 = \DFF_157.D ;
  assign II1155 = \DFF_157.D ;
  assign II1166 = \DFF_163.D ;
  assign II1169 = \DFF_163.D ;
  assign II1174 = \DFF_43.Q ;
  assign II1178 = \DFF_44.Q ;
  assign II1183 = \DFF_42.Q ;
  assign II1201 = \DFF_164.D ;
  assign II1204 = \DFF_164.D ;
  assign II1209 = \DFF_45.Q ;
  assign II1227 = \DFF_156.D ;
  assign II1230 = \DFF_156.D ;
  assign II1236 = \DFF_46.Q ;
  assign II1344 = \DFF_49.Q ;
  assign II1348 = \DFF_50.Q ;
  assign II1353 = \DFF_48.Q ;
  assign II1371 = \DFF_158.D ;
  assign II1374 = \DFF_158.D ;
  assign II1385 = \DFF_160.D ;
  assign II1388 = \DFF_160.D ;
  assign II1399 = \DFF_159.D ;
  assign II1402 = \DFF_159.D ;
  assign II1407 = \DFF_52.Q ;
  assign II1411 = \DFF_53.Q ;
  assign II1416 = \DFF_51.Q ;
  assign II1450 = \DFF_161.D ;
  assign II1453 = \DFF_161.D ;
  assign II1464 = \DFF_162.D ;
  assign II1467 = \DFF_162.D ;
  assign II1472 = \DFF_55.Q ;
  assign II1476 = \DFF_56.Q ;
  assign II1481 = \DFF_54.Q ;
  assign II1538 = \DFF_110.D ;
  assign II1550 = \DFF_111.D ;
  assign II1606 = \DFF_107.D ;
  assign II1617 = \DFF_106.D ;
  assign II1630 = \DFF_109.D ;
  assign II1703 = \DFF_108.D ;
  assign II1708 = \DFF_105.D ;
  assign II1719 = \DFF_112.D ;
  assign II1791 = \DFF_73.Q ;
  assign II1795 = \DFF_74.Q ;
  assign II1800 = \DFF_72.Q ;
  assign II1899 = \DFF_78.Q ;
  assign II1903 = \DFF_79.Q ;
  assign II1908 = \DFF_77.Q ;
  assign II196 = n3083gat;
  assign II1961 = \DFF_81.Q ;
  assign II203 = n3085gat;
  assign II2040 = \DFF_84.Q ;
  assign II2044 = \DFF_85.Q ;
  assign II2049 = \DFF_83.Q ;
  assign II210 = n3084gat;
  assign II2153 = \DFF_89.Q ;
  assign II2157 = \DFF_90.Q ;
  assign II2162 = \DFF_88.Q ;
  assign II2213 = \DFF_111.D ;
  assign II2225 = \DFF_93.Q ;
  assign II2228 = \DFF_112.D ;
  assign II2232 = \DFF_155.D ;
  assign II2235 = \DFF_155.D ;
  assign II2238 = \DFF_61.Q ;
  assign II2242 = \DFF_59.Q ;
  assign II2251 = \DFF_113.D ;
  assign II2254 = \DFF_113.D ;
  assign II2257 = \DFF_110.D ;
  assign II2260 = \DFF_114.D ;
  assign II2263 = \DFF_114.D ;
  assign II2268 = \DFF_58.Q ;
  assign II2271 = \DFF_60.Q ;
  assign II2275 = \DFF_62.Q ;
  assign II2316 = \DFF_125.D ;
  assign II2319 = \DFF_148.D ;
  assign II2344 = \DFF_124.D ;
  assign II2349 = \DFF_123.D ;
  assign II2372 = \DFF_106.D ;
  assign II2376 = \DFF_63.Q ;
  assign II2380 = \DFF_107.D ;
  assign II2385 = \DFF_108.D ;
  assign II2389 = \DFF_64.Q ;
  assign II2394 = \DFF_65.Q ;
  assign II2403 = \DFF_109.D ;
  assign II2414 = \DFF_154.D ;
  assign II2417 = \DFF_154.D ;
  assign II2420 = \DFF_105.D ;
  assign II2425 = \DFF_100.Q ;
  assign II2428 = \DFF_67.Q ;
  assign II2433 = \DFF_66.Q ;
  assign II2813 = \DFF_143.D ;
  assign II3143 = \DFF_166.D ;
  assign II3168 = \DFF_118.D ;
  assign II3315 = \DFF_132.Q ;
  assign II3318 = \DFF_132.Q ;
  assign II3339 = \DFF_133.D ;
  assign II3342 = \DFF_129.D ;
  assign II3394 = \DFF_125.Q ;
  assign II3461 = \DFF_108.Q ;
  assign II3509 = \DFF_112.Q ;
  assign II3587 = \DFF_152.D ;
  assign II359 = \DFF_23.Q ;
  assign II363 = \DFF_24.Q ;
  assign II368 = \DFF_22.Q ;
  assign II406 = \DFF_25.Q ;
  assign II409 = \DFF_41.Q ;
  assign II4117 = n3141gat;
  assign II4122 = n3141gat;
  assign II414 = \DFF_40.Q ;
  assign II4222 = n3140gat;
  assign II4227 = n3139gat;
  assign II4482 = \DFF_96.Q ;
  assign II4485 = \DFF_96.Q ;
  assign II4489 = \DFF_97.Q ;
  assign II4492 = \DFF_97.Q ;
  assign II4496 = \DFF_98.Q ;
  assign II4499 = \DFF_98.Q ;
  assign II453 = \DFF_38.Q ;
  assign II4558 = n3116gat;
  assign II456 = \DFF_39.Q ;
  assign II461 = \DFF_26.Q ;
  assign II4626 = n3106gat;
  assign II4630 = \DFF_132.Q ;
  assign II4633 = \DFF_132.Q ;
  assign II4660 = \DFF_132.Q ;
  assign II4720 = \DFF_98.Q ;
  assign II4723 = \DFF_97.Q ;
  assign II4726 = \DFF_96.Q ;
  assign II642 = \DFF_23.Q ;
  assign II646 = \DFF_24.Q ;
  assign II651 = \DFF_22.Q ;
  assign II683 = \DFF_25.Q ;
  assign II687 = \DFF_41.Q ;
  assign II692 = \DFF_40.Q ;
  assign II726 = \DFF_38.Q ;
  assign II729 = \DFF_39.Q ;
  assign II734 = \DFF_26.Q ;
  assign II842 = \DFF_29.Q ;
  assign II846 = \DFF_30.Q ;
  assign II851 = \DFF_28.Q ;
  assign II921 = \DFF_32.Q ;
  assign II925 = \DFF_33.Q ;
  assign II930 = \DFF_31.Q ;
  assign n1018gat = \DFF_40.Q ;
  assign n1019gat = \DFF_25.Q ;
  assign n1020gat = \DFF_41.Q ;
  assign n1025gat = \DFF_25.Q ;
  assign n1026gat = \DFF_25.Q ;
  assign n1034gat = \DFF_72.Q ;
  assign n1035gat = \DFF_72.Q ;
  assign n1044gat = \DFF_79.Q ;
  assign n1045gat = \DFF_79.Q ;
  assign n1055gat = \DFF_34.Q ;
  assign n1056gat = \DFF_35.Q ;
  assign n1057gat = \DFF_36.Q ;
  assign n1067gat = \DFF_28.Q ;
  assign n1068gat = \DFF_28.Q ;
  assign n1071gat = \DFF_74.Q ;
  assign n1072gat = \DFF_74.Q ;
  assign n1079gat = \DFF_35.Q ;
  assign n1080gat = \DFF_35.Q ;
  assign n1084gat = \DFF_83.Q ;
  assign n1085gat = \DFF_84.Q ;
  assign n1086gat = n3106gat;
  assign n1118gat = \DFF_72.Q ;
  assign n1120gat = \DFF_73.Q ;
  assign n1121gat = \DFF_73.Q ;
  assign n1134gat = \DFF_78.Q ;
  assign n1135gat = \DFF_78.Q ;
  assign n1147gat = \DFF_36.Q ;
  assign n1148gat = \DFF_36.Q ;
  assign n1150gat = \DFF_90.Q ;
  assign n1189gat = \DFF_72.Q ;
  assign n1190gat = \DFF_73.Q ;
  assign n1191gat = \DFF_74.Q ;
  assign n1196gat = \DFF_80.Q ;
  assign n1197gat = \DFF_80.Q ;
  assign n1206gat = \DFF_77.Q ;
  assign n1207gat = \DFF_78.Q ;
  assign n1208gat = \DFF_79.Q ;
  assign n1221gat = n3085gat;
  assign n1222gat = n3084gat;
  assign n1223gat = n3083gat;
  assign n1225gat = \DFF_76.Q ;
  assign n1226gat = \DFF_76.Q ;
  assign n1233gat = \DFF_31.Q ;
  assign n1234gat = \DFF_32.Q ;
  assign n1235gat = \DFF_33.Q ;
  assign n1240gat = \DFF_32.Q ;
  assign n1241gat = \DFF_32.Q ;
  assign n1269gat = n3116gat;
  assign n1281gat = \DFF_75.Q ;
  assign n1282gat = \DFF_75.Q ;
  assign n1293gat = \DFF_31.Q ;
  assign n1294gat = \DFF_31.Q ;
  assign n1297gat = \DFF_33.Q ;
  assign n1298gat = \DFF_33.Q ;
  assign n1311gat = \DFF_130.Q ;
  assign n1312gat = \DFF_130.Q ;
  assign n1314gat = \DFF_129.D ;
  assign n1315gat = \DFF_128.Q ;
  assign n1316gat = \DFF_128.Q ;
  assign n1328gat = \DFF_76.Q ;
  assign n1330gat = \DFF_121.D ;
  assign n1332gat = \DFF_120.Q ;
  assign n1336gat = \DFF_169.Q ;
  assign n1339gat = \DFF_173.Q ;
  assign n1340gat = \DFF_173.Q ;
  assign n1350gat = \DFF_104.D ;
  assign n1361gat = \DFF_130.D ;
  assign n1363gat = \DFF_129.Q ;
  assign n1382gat = \DFF_75.Q ;
  assign n1389gat = \DFF_115.Q ;
  assign n1391gat = \DFF_169.D ;
  assign n1392gat = \DFF_118.D ;
  assign n1393gat = \DFF_117.Q ;
  assign n1394gat = \DFF_117.Q ;
  assign n1431gat = \DFF_128.D ;
  assign n1433gat = \DFF_127.Q ;
  assign n1442gat = \DFF_104.D ;
  assign n1455gat = \DFF_174.Q ;
  assign n1456gat = \DFF_174.Q ;
  assign n1461gat = \DFF_176.Q ;
  assign n1462gat = \DFF_176.Q ;
  assign n147gat = \DFF_165.Q ;
  assign n148gat = \DFF_165.Q ;
  assign n1495gat = \DFF_118.Q ;
  assign n1496gat = \DFF_118.Q ;
  assign n1507gat = \DFF_134.Q ;
  assign n1508gat = \DFF_134.Q ;
  assign n1516gat = \DFF_117.D ;
  assign n1518gat = \DFF_143.D ;
  assign n151gat = \DFF_157.Q ;
  assign n1524gat = \DFF_175.Q ;
  assign n1525gat = \DFF_175.Q ;
  assign n152gat = \DFF_157.Q ;
  assign n155gat = \DFF_156.Q ;
  assign n1564gat = \DFF_174.D ;
  assign n1565gat = \DFF_120.D ;
  assign n1567gat = \DFF_173.D ;
  assign n156gat = \DFF_156.Q ;
  assign n1587gat = \DFF_178.Q ;
  assign n1588gat = \DFF_178.Q ;
  assign n1593gat = \DFF_178.D ;
  assign n1595gat = \DFF_177.Q ;
  assign n1596gat = \DFF_177.Q ;
  assign n159gat = \DFF_23.Q ;
  assign n1603gat = \DFF_104.D ;
  assign n1606gat = \DFF_68.D ;
  assign n160gat = \DFF_23.Q ;
  assign n1610gat = \DFF_70.D ;
  assign n1613gat = \DFF_168.D ;
  assign n1620gat = \DFF_16.D ;
  assign n1625gat = \DFF_102.D ;
  assign n1626gat = \DFF_103.D ;
  assign n1631gat = \DFF_109.Q ;
  assign n1632gat = \DFF_175.D ;
  assign n1633gat = \DFF_107.Q ;
  assign n1636gat = \DFF_134.D ;
  assign n164gat = \DFF_23.Q ;
  assign n1658gat = \DFF_113.Q ;
  assign n165gat = \DFF_23.Q ;
  assign n1674gat = \DFF_171.Q ;
  assign n1675gat = \DFF_171.Q ;
  assign n1677gat = \DFF_135.Q ;
  assign n1678gat = \DFF_135.Q ;
  assign n1685gat = \DFF_119.D ;
  assign n1691gat = \DFF_142.Q ;
  assign n1696gat = \DFF_131.D ;
  assign n1699gat = \DFF_142.Q ;
  assign n1708gat = \DFF_124.D ;
  assign n1712gat = \DFF_135.D ;
  assign n1713gat = \DFF_171.D ;
  assign n1717gat = \DFF_172.D ;
  assign n1721gat = n3138gat;
  assign n172gat = \DFF_22.Q ;
  assign n1739gat = \DFF_121.Q ;
  assign n173gat = \DFF_23.Q ;
  assign n1740gat = \DFF_121.Q ;
  assign n1742gat = \DFF_113.Q ;
  assign n1745gat = n3107gat;
  assign n1747gat = \DFF_170.Q ;
  assign n1748gat = \DFF_170.Q ;
  assign n174gat = \DFF_24.Q ;
  assign n1762gat = \DFF_70.Q ;
  assign n1763gat = \DFF_70.Q ;
  assign n1767gat = \DFF_103.Q ;
  assign n1771gat = \DFF_168.Q ;
  assign n1773gat = \DFF_133.D ;
  assign n1774gat = \DFF_131.Q ;
  assign n1775gat = \DFF_131.Q ;
  assign n1777gat = \DFF_143.D ;
  assign n1781gat = \DFF_116.D ;
  assign n1783gat = \DFF_109.Q ;
  assign n1785gat = \DFF_106.Q ;
  assign n1787gat = \DFF_105.Q ;
  assign n1793gat = \DFF_115.D ;
  assign n1800gat = \DFF_177.D ;
  assign n1806gat = \DFF_172.Q ;
  assign n1807gat = \DFF_172.Q ;
  assign n1816gat = \DFF_20.D ;
  assign n1821gat = \DFF_19.Q ;
  assign n1825gat = \DFF_19.Q ;
  assign n1827gat = \DFF_19.D ;
  assign n1828gat = \DFF_21.Q ;
  assign n1829gat = \DFF_21.Q ;
  assign n1834gat = \DFF_102.Q ;
  assign n1836gat = \DFF_126.D ;
  assign n1845gat = \DFF_105.Q ;
  assign n1849gat = \DFF_109.Q ;
  assign n1850gat = \DFF_109.Q ;
  assign n1858gat = \DFF_71.D ;
  assign n1869gat = n3106gat;
  assign n1870gat = \DFF_132.Q ;
  assign n1871gat = \DFF_132.Q ;
  assign n1879gat = \DFF_69.Q ;
  assign n1880gat = \DFF_69.Q ;
  assign n1882gat = \DFF_69.D ;
  assign n1884gat = \DFF_108.Q ;
  assign n1886gat = \DFF_108.Q ;
  assign n1891gat = \DFF_106.Q ;
  assign n1898gat = \DFF_108.Q ;
  assign n1899gat = \DFF_108.Q ;
  assign n1915gat = \DFF_176.D ;
  assign n1918gat = \DFF_111.Q ;
  assign n1927gat = \DFF_170.D ;
  assign n1945gat = \DFF_122.D ;
  assign n1954gat = \DFF_108.Q ;
  assign n1955gat = \DFF_108.Q ;
  assign n1963gat = \DFF_107.Q ;
  assign n1974gat = \DFF_154.Q ;
  assign n1975gat = \DFF_154.Q ;
  assign n1988gat = \DFF_114.Q ;
  assign n1989gat = \DFF_110.Q ;
  assign n2009gat = \DFF_132.D ;
  assign n2015gat = \DFF_144.D ;
  assign n2017gat = \DFF_146.D ;
  assign n2021gat = \DFF_116.Q ;
  assign n2023gat = \DFF_147.D ;
  assign n2025gat = \DFF_146.Q ;
  assign n2027gat = \DFF_21.D ;
  assign n2029gat = \DFF_20.Q ;
  assign n2031gat = \DFF_150.D ;
  assign n2033gat = \DFF_149.Q ;
  assign n2035gat = \DFF_149.D ;
  assign n2037gat = \DFF_145.Q ;
  assign n2039gat = \DFF_143.Q ;
  assign n2040gat = \DFF_143.Q ;
  assign n2042gat = \DFF_145.D ;
  assign n2044gat = \DFF_144.Q ;
  assign n2046gat = \DFF_123.D ;
  assign n2057gat = \DFF_98.D ;
  assign n2060gat = \DFF_106.Q ;
  assign n2061gat = \DFF_106.Q ;
  assign n2084gat = \DFF_104.Q ;
  assign n2090gat = \DFF_119.Q ;
  assign n2091gat = \DFF_119.Q ;
  assign n2093gat = \DFF_140.D ;
  assign n2095gat = \DFF_139.Q ;
  assign n2099gat = \DFF_147.Q ;
  assign n2101gat = \DFF_68.Q ;
  assign n2102gat = \DFF_68.Q ;
  assign n2108gat = \DFF_151.D ;
  assign n2110gat = \DFF_150.Q ;
  assign n2117gat = \DFF_153.Q ;
  assign n2119gat = \DFF_153.D ;
  assign n2121gat = \DFF_152.Q ;
  assign n2123gat = \DFF_152.D ;
  assign n2124gat = \DFF_151.Q ;
  assign n2125gat = \DFF_151.Q ;
  assign n2127gat = \DFF_125.D ;
  assign n2134gat = \DFF_124.Q ;
  assign n2135gat = \DFF_124.Q ;
  assign n2138gat = \DFF_107.Q ;
  assign n2139gat = \DFF_107.Q ;
  assign n2142gat = \DFF_105.Q ;
  assign n2143gat = \DFF_105.Q ;
  assign n2154gat = \DFF_71.Q ;
  assign n2155gat = \DFF_71.Q ;
  assign n2163gat = \DFF_142.D ;
  assign n2168gat = \DFF_141.Q ;
  assign n2169gat = \DFF_141.Q ;
  assign n2174gat = \DFF_141.D ;
  assign n2176gat = \DFF_140.Q ;
  assign n2178gat = \DFF_122.Q ;
  assign n2179gat = \DFF_122.Q ;
  assign n2181gat = \DFF_126.Q ;
  assign n2182gat = \DFF_126.Q ;
  assign n2189gat = \DFF_123.Q ;
  assign n2190gat = \DFF_123.Q ;
  assign n2192gat = \DFF_96.D ;
  assign n2194gat = \DFF_97.D ;
  assign n2196gat = \DFF_60.D ;
  assign n2197gat = \DFF_62.D ;
  assign n2198gat = \DFF_59.D ;
  assign n2201gat = \DFF_114.D ;
  assign n2202gat = \DFF_60.Q ;
  assign n2203gat = \DFF_60.Q ;
  assign n2205gat = \DFF_113.D ;
  assign n2206gat = \DFF_62.Q ;
  assign n2207gat = \DFF_62.Q ;
  assign n2214gat = \DFF_62.Q ;
  assign n2217gat = \DFF_113.D ;
  assign n2251gat = \DFF_125.Q ;
  assign n2252gat = \DFF_125.Q ;
  assign n2261gat = \DFF_125.Q ;
  assign n2262gat = \DFF_125.Q ;
  assign n2265gat = \DFF_148.Q ;
  assign n2266gat = \DFF_148.Q ;
  assign n2268gat = \DFF_123.D ;
  assign n2269gat = \DFF_97.Q ;
  assign n226gat = \DFF_88.Q ;
  assign n2270gat = \DFF_97.Q ;
  assign n227gat = \DFF_89.Q ;
  assign n2283gat = \DFF_112.Q ;
  assign n2284gat = \DFF_111.D ;
  assign n2285gat = \DFF_58.Q ;
  assign n228gat = \DFF_90.Q ;
  assign n2290gat = \DFF_114.D ;
  assign n2319gat = \DFF_17.Q ;
  assign n2330gat = \DFF_64.D ;
  assign n2332gat = \DFF_112.Q ;
  assign n2333gat = \DFF_112.Q ;
  assign n2337gat = \DFF_124.D ;
  assign n2338gat = \DFF_98.Q ;
  assign n2339gat = \DFF_98.Q ;
  assign n2341gat = \DFF_111.D ;
  assign n2342gat = \DFF_59.Q ;
  assign n2343gat = \DFF_59.Q ;
  assign n2346gat = \DFF_114.Q ;
  assign n2347gat = \DFF_114.Q ;
  assign n2351gat = \DFF_113.Q ;
  assign n2353gat = \DFF_110.D ;
  assign n2354gat = \DFF_60.Q ;
  assign n2355gat = \DFF_59.Q ;
  assign n2356gat = \DFF_61.Q ;
  assign n2387gat = \DFF_65.D ;
  assign n2388gat = \DFF_125.D ;
  assign n2389gat = \DFF_96.Q ;
  assign n2390gat = \DFF_96.Q ;
  assign n2393gat = \DFF_111.Q ;
  assign n2394gat = \DFF_111.Q ;
  assign n2396gat = \DFF_58.D ;
  assign n2397gat = \DFF_110.D ;
  assign n2398gat = \DFF_58.Q ;
  assign n2399gat = \DFF_58.Q ;
  assign n2402gat = \DFF_110.Q ;
  assign n2403gat = \DFF_110.Q ;
  assign n2406gat = \DFF_113.Q ;
  assign n2407gat = \DFF_113.Q ;
  assign n2414gat = \DFF_62.Q ;
  assign n2415gat = \DFF_58.Q ;
  assign n2416gat = \DFF_60.Q ;
  assign n2417gat = \DFF_110.D ;
  assign n2418gat = \DFF_114.D ;
  assign n2419gat = \DFF_113.D ;
  assign n2429gat = \DFF_67.Q ;
  assign n2436gat = \DFF_67.D ;
  assign n2439gat = \DFF_112.Q ;
  assign n2440gat = \DFF_112.Q ;
  assign n2443gat = \DFF_112.D ;
  assign n2454gat = \DFF_142.Q ;
  assign n2456gat = \DFF_167.D ;
  assign n2458gat = \DFF_166.Q ;
  assign n2464gat = \DFF_57.Q ;
  assign n2468gat = \DFF_37.Q ;
  assign n2470gat = \DFF_17.D ;
  assign n2472gat = \DFF_16.Q ;
  assign n2476gat = \DFF_27.Q ;
  assign n2482gat = \DFF_105.D ;
  assign n2486gat = \DFF_109.D ;
  assign n2487gat = \DFF_107.D ;
  assign n2488gat = \DFF_107.D ;
  assign n2489gat = \DFF_64.Q ;
  assign n2490gat = \DFF_64.Q ;
  assign n2492gat = \DFF_95.D ;
  assign n2493gat = \DFF_148.D ;
  assign n2494gat = \DFF_95.Q ;
  assign n2495gat = \DFF_95.Q ;
  assign n2498gat = \DFF_61.D ;
  assign n2502gat = \DFF_99.Q ;
  assign n2506gat = \DFF_101.Q ;
  assign n2510gat = \DFF_9.Q ;
  assign n2514gat = \DFF_167.Q ;
  assign n2518gat = \DFF_81.Q ;
  assign n2522gat = \DFF_27.Q ;
  assign n2526gat = \DFF_47.Q ;
  assign n2532gat = \DFF_108.D ;
  assign n2536gat = \DFF_63.Q ;
  assign n2539gat = \DFF_63.D ;
  assign n2540gat = \DFF_64.Q ;
  assign n2541gat = \DFF_105.D ;
  assign n2542gat = \DFF_67.Q ;
  assign n2543gat = \DFF_67.Q ;
  assign n2550gat = \DFF_66.Q ;
  assign n2551gat = \DFF_100.Q ;
  assign n2552gat = \DFF_67.Q ;
  assign n2553gat = \DFF_154.D ;
  assign n2554gat = \DFF_105.D ;
  assign n2555gat = \DFF_109.D ;
  assign n2556gat = \DFF_66.D ;
  assign n2557gat = \DFF_106.D ;
  assign n2558gat = \DFF_100.D ;
  assign n255gat = \DFF_163.Q ;
  assign n2560gat = \DFF_112.D ;
  assign n2561gat = \DFF_61.Q ;
  assign n2562gat = \DFF_61.Q ;
  assign n256gat = \DFF_163.Q ;
  assign n2573gat = \DFF_59.Q ;
  assign n2574gat = \DFF_155.D ;
  assign n2575gat = \DFF_61.Q ;
  assign n2576gat = \DFF_93.Q ;
  assign n2577gat = \DFF_112.D ;
  assign n2578gat = \DFF_111.D ;
  assign n2579gat = \DFF_94.D ;
  assign n2588gat = \DFF_92.Q ;
  assign n2590gat = \DFF_166.D ;
  assign n2591gat = \DFF_133.Q ;
  assign n2592gat = \DFF_133.Q ;
  assign n2599gat = \DFF_91.Q ;
  assign n2606gat = \DFF_65.Q ;
  assign n2607gat = \DFF_108.D ;
  assign n2608gat = \DFF_64.Q ;
  assign n2609gat = \DFF_63.Q ;
  assign n2610gat = \DFF_107.D ;
  assign n2611gat = \DFF_106.D ;
  assign n2612gat = \DFF_65.Q ;
  assign n2613gat = \DFF_101.D ;
  assign n2620gat = \DFF_106.D ;
  assign n2621gat = \DFF_65.Q ;
  assign n2622gat = \DFF_65.Q ;
  assign n2624gat = \DFF_108.D ;
  assign n2625gat = \DFF_63.Q ;
  assign n2626gat = \DFF_63.Q ;
  assign n2628gat = \DFF_109.D ;
  assign n2629gat = \DFF_66.Q ;
  assign n2630gat = \DFF_66.Q ;
  assign n2632gat = \DFF_154.D ;
  assign n2633gat = \DFF_100.Q ;
  assign n2634gat = \DFF_100.Q ;
  assign n2636gat = \DFF_93.D ;
  assign n2638gat = \DFF_155.D ;
  assign n2639gat = \DFF_93.Q ;
  assign n263gat = \DFF_22.Q ;
  assign n2640gat = \DFF_93.Q ;
  assign n2643gat = \DFF_155.Q ;
  assign n2644gat = \DFF_155.Q ;
  assign n2646gat = \DFF_99.D ;
  assign n264gat = \DFF_23.Q ;
  assign n2658gat = \DFF_94.Q ;
  assign n265gat = \DFF_24.Q ;
  assign n2667gat = n3095gat;
  assign n2668gat = n3095gat;
  assign n2670gat = n3072gat;
  assign n2671gat = n3072gat;
  assign n2673gat = n3073gat;
  assign n2674gat = n3073gat;
  assign n2677gat = \DFF_123.D ;
  assign n2678gat = \DFF_125.D ;
  assign n2680gat = n3150gat;
  assign n2681gat = \DFF_123.D ;
  assign n2682gat = \DFF_125.D ;
  assign n2684gat = n3150gat;
  assign n2685gat = n3116gat;
  assign n2686gat = \DFF_124.D ;
  assign n2688gat = \DFF_124.D ;
  assign n2689gat = n3114gat;
  assign n2691gat = n3146gat;
  assign n2692gat = \DFF_104.D ;
  assign n2693gat = n3114gat;
  assign n2696gat = \DFF_104.D ;
  assign n2698gat = n3113gat;
  assign n2699gat = n3145gat;
  assign n2700gat = n3151gat;
  assign n2702gat = n3113gat;
  assign n2704gat = n3151gat;
  assign n2705gat = n3110gat;
  assign n2706gat = n3111gat;
  assign n2708gat = n3110gat;
  assign n2709gat = n3111gat;
  assign n270gat = \DFF_22.Q ;
  assign n2712gat = n3075gat;
  assign n2716gat = n3088gat;
  assign n2717gat = n3088gat;
  assign n2719gat = n3074gat;
  assign n271gat = \DFF_22.Q ;
  assign n2721gat = n3094gat;
  assign n2722gat = n3094gat;
  assign n2724gat = n3087gat;
  assign n2725gat = n3087gat;
  assign n2727gat = n3086gat;
  assign n2728gat = n3086gat;
  assign n2729gat = n3099gat;
  assign n2730gat = n3099gat;
  assign n2732gat = n3065gat;
  assign n2733gat = n3065gat;
  assign n2735gat = n3066gat;
  assign n2736gat = n3066gat;
  assign n2737gat = n3117gat;
  assign n2738gat = n3118gat;
  assign n2739gat = n3139gat;
  assign n2740gat = n3144gat;
  assign n2741gat = n3117gat;
  assign n2742gat = n3118gat;
  assign n2744gat = n3144gat;
  assign n2745gat = n3119gat;
  assign n2746gat = n3120gat;
  assign n2747gat = n3140gat;
  assign n2748gat = n3141gat;
  assign n2749gat = n3119gat;
  assign n274gat = \DFF_26.Q ;
  assign n2750gat = n3120gat;
  assign n2753gat = n3121gat;
  assign n2754gat = n3122gat;
  assign n2755gat = n3141gat;
  assign n2756gat = n3121gat;
  assign n2757gat = n3122gat;
  assign n2759gat = n3123gat;
  assign n275gat = \DFF_26.Q ;
  assign n2760gat = n3124gat;
  assign n2761gat = n3123gat;
  assign n2762gat = n3124gat;
  assign n2763gat = n3125gat;
  assign n2764gat = n3125gat;
  assign n2765gat = n3098gat;
  assign n2766gat = n3098gat;
  assign n2767gat = n3093gat;
  assign n2768gat = n3093gat;
  assign n2776gat = n3067gat;
  assign n2777gat = n3067gat;
  assign n2779gat = n3068gat;
  assign n2780gat = n3068gat;
  assign n2782gat = n3069gat;
  assign n2783gat = n3069gat;
  assign n278gat = \DFF_24.Q ;
  assign n2790gat = n3070gat;
  assign n2791gat = n3070gat;
  assign n2793gat = n3071gat;
  assign n2794gat = n3071gat;
  assign n2795gat = n3108gat;
  assign n2796gat = n3109gat;
  assign n2797gat = n3143gat;
  assign n2798gat = n3108gat;
  assign n2799gat = n3109gat;
  assign n279gat = \DFF_24.Q ;
  assign n2800gat = n3143gat;
  assign n2801gat = n3106gat;
  assign n2802gat = n3107gat;
  assign n2803gat = n3129gat;
  assign n2804gat = n3138gat;
  assign n2805gat = n3106gat;
  assign n2806gat = n3107gat;
  assign n2807gat = n3129gat;
  assign n2808gat = n3138gat;
  assign n2809gat = n3105gat;
  assign n2810gat = n3136gat;
  assign n2811gat = n3137gat;
  assign n2812gat = n3105gat;
  assign n2813gat = n3136gat;
  assign n2814gat = n3137gat;
  assign n2815gat = n3134gat;
  assign n2816gat = n3135gat;
  assign n2817gat = n3134gat;
  assign n2818gat = n3135gat;
  assign n2819gat = n3104gat;
  assign n2820gat = n3132gat;
  assign n2821gat = n3133gat;
  assign n2822gat = n3104gat;
  assign n2823gat = n3132gat;
  assign n2824gat = n3133gat;
  assign n2825gat = n3130gat;
  assign n2826gat = n3131gat;
  assign n2828gat = n3130gat;
  assign n2829gat = n3131gat;
  assign n282gat = \DFF_22.Q ;
  assign n2831gat = n3090gat;
  assign n2832gat = n3090gat;
  assign n2837gat = n3077gat;
  assign n2839gat = n3076gat;
  assign n283gat = \DFF_22.Q ;
  assign n2841gat = n3079gat;
  assign n2843gat = n3078gat;
  assign n2845gat = n3081gat;
  assign n2847gat = n3080gat;
  assign n2850gat = n3100gat;
  assign n2851gat = n3100gat;
  assign n2853gat = n3082gat;
  assign n2855gat = n3083gat;
  assign n2856gat = n3083gat;
  assign n2858gat = n3097gat;
  assign n2860gat = n3085gat;
  assign n2861gat = n3085gat;
  assign n2863gat = n3084gat;
  assign n2864gat = n3084gat;
  assign n2868gat = n3089gat;
  assign n2869gat = n3089gat;
  assign n2886gat = \DFF_90.D ;
  assign n2887gat = \DFF_89.D ;
  assign n2888gat = \DFF_88.D ;
  assign n2890gat = \DFF_87.D ;
  assign n2891gat = \DFF_83.D ;
  assign n2892gat = \DFF_46.D ;
  assign n2894gat = \DFF_34.D ;
  assign n2895gat = \DFF_36.D ;
  assign n2896gat = \DFF_31.D ;
  assign n2897gat = \DFF_33.D ;
  assign n2898gat = \DFF_54.D ;
  assign n2899gat = \DFF_56.D ;
  assign n2900gat = \DFF_51.D ;
  assign n2901gat = \DFF_86.D ;
  assign n2903gat = \DFF_84.D ;
  assign n2904gat = \DFF_82.D ;
  assign n2905gat = \DFF_50.D ;
  assign n2907gat = \DFF_76.D ;
  assign n2908gat = \DFF_80.D ;
  assign n2909gat = \DFF_79.D ;
  assign n2910gat = \DFF_75.D ;
  assign n2911gat = \DFF_77.D ;
  assign n2912gat = \DFF_78.D ;
  assign n2913gat = \DFF_48.D ;
  assign n2914gat = \DFF_28.D ;
  assign n2915gat = \DFF_85.D ;
  assign n2916gat = \DFF_55.D ;
  assign n2917gat = \DFF_43.D ;
  assign n2918gat = \DFF_72.D ;
  assign n2919gat = \DFF_74.D ;
  assign n2920gat = \DFF_49.D ;
  assign n2921gat = \DFF_35.D ;
  assign n2922gat = \DFF_32.D ;
  assign n2923gat = \DFF_42.D ;
  assign n2924gat = \DFF_44.D ;
  assign n2925gat = \DFF_52.D ;
  assign n2926gat = \DFF_45.D ;
  assign n2927gat = \DFF_30.D ;
  assign n2928gat = \DFF_29.D ;
  assign n2929gat = \DFF_53.D ;
  assign n2935gat = n3135gat;
  assign n2936gat = n3131gat;
  assign n2937gat = n3134gat;
  assign n2938gat = n3132gat;
  assign n2941gat = n3137gat;
  assign n2950gat = n3136gat;
  assign n2951gat = n3129gat;
  assign n2952gat = \DFF_73.D ;
  assign n2955gat = n3130gat;
  assign n2956gat = n3133gat;
  assign n2971gat = \DFF_81.D ;
  assign n2980gat = n3141gat;
  assign n2983gat = \DFF_127.D ;
  assign n2989gat = \DFF_71.D ;
  assign n3010gat = \DFF_91.D ;
  assign n3016gat = \DFF_92.D ;
  assign n3020gat = \DFF_142.Q ;
  assign n3021gat = \DFF_142.Q ;
  assign n3022gat = \DFF_142.Q ;
  assign n3023gat = \DFF_142.Q ;
  assign n3024gat = \DFF_142.Q ;
  assign n3025gat = \DFF_142.Q ;
  assign n3026gat = \DFF_142.Q ;
  assign n3027gat = \DFF_142.Q ;
  assign n3028gat = \DFF_142.Q ;
  assign n3029gat = n3106gat;
  assign n3030gat = n3106gat;
  assign n3031gat = \DFF_97.D ;
  assign n3032gat = \DFF_125.Q ;
  assign n3034gat = \DFF_96.D ;
  assign n3035gat = \DFF_98.D ;
  assign n3036gat = \DFF_95.D ;
  assign n3037gat = \DFF_66.D ;
  assign n3039gat = \DFF_108.Q ;
  assign n3040gat = \DFF_63.D ;
  assign n3041gat = \DFF_67.D ;
  assign n3042gat = \DFF_65.D ;
  assign n3043gat = \DFF_107.Q ;
  assign n3044gat = \DFF_64.D ;
  assign n3046gat = \DFF_112.Q ;
  assign n3047gat = \DFF_61.D ;
  assign n3048gat = \DFF_58.D ;
  assign n3049gat = \DFF_59.D ;
  assign n3050gat = \DFF_62.D ;
  assign n3051gat = \DFF_60.D ;
  assign n3052gat = \DFF_69.D ;
  assign n3053gat = \DFF_100.D ;
  assign n3054gat = \DFF_93.D ;
  assign n3055gat = \DFF_43.D ;
  assign n3056gat = \DFF_46.D ;
  assign n3057gat = \DFF_51.D ;
  assign n3058gat = \DFF_53.D ;
  assign n3059gat = \DFF_52.D ;
  assign n3060gat = \DFF_55.D ;
  assign n3061gat = \DFF_56.D ;
  assign n3062gat = \DFF_45.D ;
  assign n3063gat = \DFF_44.D ;
  assign n3064gat = \DFF_42.D ;
  assign n3112gat = 1'b1;
  assign n3115gat = 1'b1;
  assign n3126gat = \DFF_124.D ;
  assign n3127gat = \DFF_123.D ;
  assign n3128gat = \DFF_125.D ;
  assign n313gat = \DFF_90.Q ;
  assign n3142gat = n3141gat;
  assign n3147gat = 1'b1;
  assign n3148gat = 1'b1;
  assign n3149gat = \DFF_104.D ;
  assign n314gat = \DFF_90.Q ;
  assign n3152gat = 1'b1;
  assign n317gat = \DFF_89.Q ;
  assign n318gat = \DFF_89.Q ;
  assign n321gat = \DFF_88.Q ;
  assign n322gat = \DFF_88.Q ;
  assign n326gat = \DFF_161.Q ;
  assign n327gat = \DFF_161.Q ;
  assign n330gat = \DFF_158.Q ;
  assign n331gat = \DFF_158.Q ;
  assign n336gat = \DFF_24.Q ;
  assign n337gat = \DFF_24.Q ;
  assign n340gat = \DFF_26.Q ;
  assign n341gat = \DFF_26.Q ;
  assign n348gat = \DFF_26.Q ;
  assign n349gat = \DFF_38.Q ;
  assign n350gat = \DFF_39.Q ;
  assign n365gat = \DFF_87.Q ;
  assign n366gat = \DFF_87.Q ;
  assign n383gat = \DFF_162.Q ;
  assign n384gat = \DFF_162.Q ;
  assign n387gat = \DFF_159.Q ;
  assign n388gat = \DFF_159.Q ;
  assign n393gat = \DFF_39.Q ;
  assign n394gat = \DFF_39.Q ;
  assign n397gat = \DFF_39.Q ;
  assign n398gat = \DFF_39.Q ;
  assign n401gat = \DFF_38.Q ;
  assign n402gat = \DFF_38.Q ;
  assign n43gat = \DFF_27.D ;
  assign n462gat = \DFF_160.Q ;
  assign n463gat = \DFF_160.Q ;
  assign n469gat = \DFF_164.Q ;
  assign n470gat = \DFF_164.Q ;
  assign n480gat = \DFF_26.Q ;
  assign n481gat = \DFF_38.Q ;
  assign n482gat = \DFF_39.Q ;
  assign n490gat = \DFF_39.Q ;
  assign n491gat = \DFF_39.Q ;
  assign n498gat = \DFF_46.Q ;
  assign n499gat = \DFF_38.Q ;
  assign n500gat = \DFF_39.Q ;
  assign n503gat = \DFF_156.D ;
  assign n504gat = \DFF_47.D ;
  assign n552gat = \DFF_84.Q ;
  assign n553gat = \DFF_84.Q ;
  assign n55gat = \DFF_27.D ;
  assign n560gat = \DFF_86.Q ;
  assign n561gat = \DFF_86.Q ;
  assign n566gat = \DFF_87.Q ;
  assign n567gat = \DFF_57.D ;
  assign n579gat = \DFF_50.Q ;
  assign n580gat = \DFF_50.Q ;
  assign n583gat = \DFF_54.Q ;
  assign n584gat = \DFF_54.Q ;
  assign n591gat = \DFF_51.Q ;
  assign n592gat = \DFF_52.Q ;
  assign n593gat = \DFF_53.Q ;
  assign n594gat = \DFF_160.D ;
  assign n595gat = \DFF_159.D ;
  assign n596gat = \DFF_158.D ;
  assign n612gat = \DFF_156.D ;
  assign n613gat = \DFF_46.Q ;
  assign n614gat = \DFF_46.Q ;
  assign n617gat = \DFF_38.Q ;
  assign n618gat = \DFF_38.Q ;
  assign n621gat = \DFF_40.Q ;
  assign n622gat = \DFF_40.Q ;
  assign n625gat = \DFF_41.Q ;
  assign n626gat = \DFF_41.Q ;
  assign n658gat = \DFF_83.Q ;
  assign n659gat = \DFF_83.Q ;
  assign n666gat = \DFF_82.Q ;
  assign n667gat = \DFF_82.Q ;
  assign n672gat = \DFF_33.Q ;
  assign n673gat = \DFF_33.Q ;
  assign n679gat = \DFF_48.Q ;
  assign n680gat = \DFF_48.Q ;
  assign n682gat = \DFF_161.D ;
  assign n683gat = \DFF_55.Q ;
  assign n684gat = \DFF_55.Q ;
  assign n691gat = \DFF_54.Q ;
  assign n692gat = \DFF_55.Q ;
  assign n693gat = \DFF_56.Q ;
  assign n694gat = \DFF_161.D ;
  assign n695gat = \DFF_162.D ;
  assign n697gat = \DFF_162.D ;
  assign n698gat = \DFF_56.Q ;
  assign n699gat = \DFF_56.Q ;
  assign n702gat = \DFF_38.Q ;
  assign n703gat = \DFF_38.Q ;
  assign n705gat = \DFF_157.D ;
  assign n706gat = \DFF_43.Q ;
  assign n707gat = \DFF_43.Q ;
  assign n714gat = \DFF_42.Q ;
  assign n715gat = \DFF_43.Q ;
  assign n716gat = \DFF_44.Q ;
  assign n717gat = \DFF_157.D ;
  assign n718gat = \DFF_163.D ;
  assign n719gat = \DFF_165.D ;
  assign n721gat = \DFF_41.Q ;
  assign n722gat = \DFF_41.Q ;
  assign n725gat = \DFF_40.Q ;
  assign n726gat = \DFF_40.Q ;
  assign n733gat = \DFF_40.Q ;
  assign n734gat = \DFF_45.Q ;
  assign n735gat = \DFF_41.Q ;
  assign n736gat = \DFF_164.D ;
  assign n748gat = \DFF_9.D ;
  assign n776gat = \DFF_85.Q ;
  assign n777gat = \DFF_85.Q ;
  assign n784gat = \DFF_83.Q ;
  assign n785gat = \DFF_84.Q ;
  assign n786gat = \DFF_85.Q ;
  assign n808gat = \DFF_48.Q ;
  assign n809gat = \DFF_49.Q ;
  assign n810gat = \DFF_50.Q ;
  assign n815gat = \DFF_49.Q ;
  assign n816gat = \DFF_49.Q ;
  assign n818gat = \DFF_160.D ;
  assign n819gat = \DFF_52.Q ;
  assign n820gat = \DFF_52.Q ;
  assign n822gat = \DFF_158.D ;
  assign n823gat = \DFF_51.Q ;
  assign n824gat = \DFF_51.Q ;
  assign n827gat = \DFF_139.D ;
  assign n828gat = \DFF_164.D ;
  assign n829gat = \DFF_45.Q ;
  assign n830gat = \DFF_45.Q ;
  assign n832gat = \DFF_165.D ;
  assign n833gat = \DFF_42.Q ;
  assign n834gat = \DFF_42.Q ;
  assign n836gat = \DFF_163.D ;
  assign n837gat = \DFF_44.Q ;
  assign n838gat = \DFF_44.Q ;
  assign n841gat = \DFF_25.Q ;
  assign n842gat = \DFF_25.Q ;
  assign n845gat = \DFF_40.Q ;
  assign n846gat = \DFF_40.Q ;
  assign n850gat = \DFF_77.Q ;
  assign n860gat = \DFF_30.Q ;
  assign n861gat = \DFF_30.Q ;
  assign n864gat = \DFF_34.Q ;
  assign n865gat = \DFF_34.Q ;
  assign n873gat = \DFF_89.Q ;
  assign n875gat = \DFF_86.Q ;
  assign n881gat = \DFF_159.D ;
  assign n882gat = \DFF_53.Q ;
  assign n883gat = \DFF_53.Q ;
  assign n911gat = \DFF_40.Q ;
  assign n912gat = \DFF_25.Q ;
  assign n913gat = \DFF_41.Q ;
  assign n918gat = \DFF_41.Q ;
  assign n919gat = \DFF_41.Q ;
  assign n922gat = \DFF_73.Q ;
  assign n923gat = \DFF_79.Q ;
  assign n924gat = \DFF_74.Q ;
  assign n927gat = \DFF_78.Q ;
  assign n930gat = \DFF_77.Q ;
  assign n931gat = \DFF_77.Q ;
  assign n933gat = \DFF_37.D ;
  assign n949gat = \DFF_28.Q ;
  assign n950gat = \DFF_29.Q ;
  assign n951gat = \DFF_30.Q ;
  assign n956gat = \DFF_29.Q ;
  assign n957gat = \DFF_29.Q ;
  assign n983gat = \DFF_88.Q ;
  assign n985gat = \DFF_85.Q ;
endmodule
