
module c880(L1, L8, L13, L17, L26, L29, L36, L42, L51, L55, L59, L68, L72, L73, L74, L75, L80, L85, L86, L87, L88, L89, L90, L91, L96, L101, L106, L111, L116, L121, L126, L130, L135, L138, L143, L146, L149, L152, L153, L156, L159, L165, L171, L177, L183, L189, L195, L201, L207, L210, L219, L228, L237, L246, L255, L259, L260, L261, L267, L268, L388, L389, L390, L391, L418, L419, L420, L421, L422, L423, L446, L447, L448, L449, L450, L767, L768, L850, L863, L864, L865, L866, L874, L878, L879, L880);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  input L1;
  input L101;
  input L106;
  input L111;
  input L116;
  input L121;
  input L126;
  input L13;
  input L130;
  input L135;
  input L138;
  input L143;
  input L146;
  input L149;
  input L152;
  input L153;
  input L156;
  input L159;
  input L165;
  input L17;
  input L171;
  input L177;
  input L183;
  input L189;
  input L195;
  input L201;
  input L207;
  input L210;
  input L219;
  input L228;
  input L237;
  input L246;
  input L255;
  input L259;
  input L26;
  input L260;
  input L261;
  input L267;
  input L268;
  wire L273;
  wire L276;
  input L29;
  wire L290;
  wire L291;
  wire L292;
  wire L297;
  wire L342;
  wire L344;
  wire L351;
  wire L353;
  wire L354;
  wire L356;
  input L36;
  wire L369;
  output L388;
  output L389;
  output L390;
  output L391;
  wire L392;
  wire L393;
  wire L399;
  wire L401;
  wire L402;
  wire L403;
  output L418;
  output L419;
  input L42;
  output L420;
  output L421;
  output L422;
  output L423;
  output L446;
  output L447;
  output L448;
  output L449;
  output L450;
  input L51;
  input L55;
  input L59;
  wire L660;
  wire L661;
  input L68;
  input L72;
  input L73;
  input L74;
  input L75;
  output L767;
  output L768;
  input L8;
  input L80;
  wire L811;
  wire L837;
  wire L838;
  wire L839;
  wire L840;
  input L85;
  output L850;
  wire L854;
  wire L855;
  wire L856;
  wire L857;
  wire L858;
  input L86;
  output L863;
  output L864;
  output L865;
  output L866;
  wire L867;
  wire L868;
  wire L869;
  input L87;
  wire L870;
  output L874;
  wire L875;
  wire L876;
  wire L877;
  output L878;
  output L879;
  input L88;
  output L880;
  input L89;
  input L90;
  input L91;
  input L96;
  al_and3 _196_ (
    .a(L1),
    .b(L26),
    .c(L51),
    .y(L447)
  );
  al_nand2 _197_ (
    .a(L59),
    .b(L156),
    .y(_184_)
  );
  al_nand3 _198_ (
    .a(L17),
    .b(_184_),
    .c(L447),
    .y(_185_)
  );
  al_nand2 _199_ (
    .a(L1),
    .b(_185_),
    .y(_186_)
  );
  al_nand3 _200_ (
    .a(L59),
    .b(L42),
    .c(L75),
    .y(_187_)
  );
  al_and2 _201_ (
    .a(L17),
    .b(L51),
    .y(_188_)
  );
  al_nand2 _202_ (
    .a(L1),
    .b(L8),
    .y(_189_)
  );
  al_and3ftt _203_ (
    .a(_189_),
    .b(_187_),
    .c(_188_),
    .y(_190_)
  );
  al_nor2 _204_ (
    .a(L17),
    .b(L42),
    .y(_191_)
  );
  al_nand2 _205_ (
    .a(L17),
    .b(L42),
    .y(_192_)
  );
  al_and3fft _206_ (
    .a(_191_),
    .b(_184_),
    .c(_192_),
    .y(_193_)
  );
  al_ao21 _207_ (
    .a(L447),
    .b(_193_),
    .c(_190_),
    .y(_194_)
  );
  al_and3 _208_ (
    .a(L29),
    .b(L80),
    .c(L75),
    .y(_195_)
  );
  al_nand2ft _209_ (
    .a(L268),
    .b(L55),
    .y(_000_)
  );
  al_and3ftt _210_ (
    .a(_000_),
    .b(L447),
    .c(_195_),
    .y(_001_)
  );
  al_aoi21 _211_ (
    .a(L111),
    .b(_194_),
    .c(_001_),
    .y(_002_)
  );
  al_ao21ttf _212_ (
    .a(L143),
    .b(_186_),
    .c(_002_),
    .y(_003_)
  );
  al_and2 _213_ (
    .a(L183),
    .b(_003_),
    .y(_004_)
  );
  al_nor2 _214_ (
    .a(L183),
    .b(_003_),
    .y(_005_)
  );
  al_nor2 _215_ (
    .a(_004_),
    .b(_005_),
    .y(_006_)
  );
  al_aoi21 _216_ (
    .a(L146),
    .b(_186_),
    .c(_001_),
    .y(_007_)
  );
  al_ao21ttf _217_ (
    .a(L116),
    .b(_194_),
    .c(_007_),
    .y(_008_)
  );
  al_nor2 _218_ (
    .a(L189),
    .b(_008_),
    .y(_009_)
  );
  al_and2 _219_ (
    .a(L189),
    .b(_008_),
    .y(_010_)
  );
  al_inv _220_ (
    .a(L195),
    .y(_011_)
  );
  al_nand2 _221_ (
    .a(L121),
    .b(_194_),
    .y(_012_)
  );
  al_aoi21 _222_ (
    .a(L149),
    .b(_186_),
    .c(_001_),
    .y(_013_)
  );
  al_aoi21 _223_ (
    .a(_013_),
    .b(_012_),
    .c(_011_),
    .y(_014_)
  );
  al_and3 _224_ (
    .a(_011_),
    .b(_013_),
    .c(_012_),
    .y(_015_)
  );
  al_inv _225_ (
    .a(L201),
    .y(_016_)
  );
  al_nand2 _226_ (
    .a(L126),
    .b(_194_),
    .y(_017_)
  );
  al_aoi21 _227_ (
    .a(L153),
    .b(_186_),
    .c(_001_),
    .y(_018_)
  );
  al_and3 _228_ (
    .a(_016_),
    .b(_018_),
    .c(_017_),
    .y(_019_)
  );
  al_inv _229_ (
    .a(L126),
    .y(_020_)
  );
  al_ao21ftf _230_ (
    .a(_020_),
    .b(_194_),
    .c(_018_),
    .y(_021_)
  );
  al_ao21 _231_ (
    .a(L201),
    .b(_021_),
    .c(L261),
    .y(_022_)
  );
  al_nand3fft _232_ (
    .a(_015_),
    .b(_019_),
    .c(_022_),
    .y(_023_)
  );
  al_nand3fft _233_ (
    .a(_010_),
    .b(_014_),
    .c(_023_),
    .y(_024_)
  );
  al_ao21ftt _234_ (
    .a(_009_),
    .b(_024_),
    .c(_006_),
    .y(_025_)
  );
  al_nand3ftt _235_ (
    .a(_009_),
    .b(_006_),
    .c(_024_),
    .y(_026_)
  );
  al_nand3 _236_ (
    .a(L219),
    .b(_026_),
    .c(_025_),
    .y(_027_)
  );
  al_inv _237_ (
    .a(L237),
    .y(_028_)
  );
  al_nand2 _238_ (
    .a(L106),
    .b(L210),
    .y(_029_)
  );
  al_or3fft _239_ (
    .a(L13),
    .b(L55),
    .c(_189_),
    .y(_030_)
  );
  al_nand2 _240_ (
    .a(L59),
    .b(L68),
    .y(_031_)
  );
  al_and3 _241_ (
    .a(L42),
    .b(L72),
    .c(L73),
    .y(_032_)
  );
  al_and3fft _242_ (
    .a(_031_),
    .b(_030_),
    .c(_032_),
    .y(_033_)
  );
  al_ao21ttf _243_ (
    .a(L183),
    .b(_033_),
    .c(_029_),
    .y(_034_)
  );
  al_aoi21 _244_ (
    .a(L246),
    .b(_003_),
    .c(_034_),
    .y(_035_)
  );
  al_ao21ftf _245_ (
    .a(_028_),
    .b(_004_),
    .c(_035_),
    .y(_036_)
  );
  al_aoi21 _246_ (
    .a(L228),
    .b(_006_),
    .c(_036_),
    .y(_037_)
  );
  al_nand2 _247_ (
    .a(_037_),
    .b(_027_),
    .y(L863)
  );
  al_or2 _248_ (
    .a(_010_),
    .b(_009_),
    .y(_038_)
  );
  al_nand3ftt _249_ (
    .a(_014_),
    .b(_023_),
    .c(_038_),
    .y(_039_)
  );
  al_ao21ftt _250_ (
    .a(_014_),
    .b(_023_),
    .c(_038_),
    .y(_040_)
  );
  al_nand3 _251_ (
    .a(L219),
    .b(_039_),
    .c(_040_),
    .y(_041_)
  );
  al_nand2 _252_ (
    .a(L255),
    .b(L259),
    .y(_042_)
  );
  al_aoi21ttf _253_ (
    .a(L111),
    .b(L210),
    .c(_042_),
    .y(_043_)
  );
  al_ao21ttf _254_ (
    .a(L189),
    .b(_033_),
    .c(_043_),
    .y(_044_)
  );
  al_aoi21 _255_ (
    .a(L246),
    .b(_008_),
    .c(_044_),
    .y(_045_)
  );
  al_ao21ftf _256_ (
    .a(_028_),
    .b(_010_),
    .c(_045_),
    .y(_046_)
  );
  al_oa21ftf _257_ (
    .a(L228),
    .b(_038_),
    .c(_046_),
    .y(_047_)
  );
  al_nand2 _258_ (
    .a(_047_),
    .b(_041_),
    .y(L864)
  );
  al_ao21 _259_ (
    .a(_018_),
    .b(_017_),
    .c(_016_),
    .y(_048_)
  );
  al_ao21ftt _260_ (
    .a(L261),
    .b(_048_),
    .c(_019_),
    .y(_049_)
  );
  al_nor2 _261_ (
    .a(_015_),
    .b(_014_),
    .y(_050_)
  );
  al_oa21ftt _262_ (
    .a(_049_),
    .b(_050_),
    .c(L219),
    .y(_051_)
  );
  al_ao21ftf _263_ (
    .a(_049_),
    .b(_050_),
    .c(_051_),
    .y(_052_)
  );
  al_ao21ttf _264_ (
    .a(_013_),
    .b(_012_),
    .c(L246),
    .y(_053_)
  );
  al_nand2 _265_ (
    .a(L255),
    .b(L260),
    .y(_054_)
  );
  al_aoi21ttf _266_ (
    .a(L116),
    .b(L210),
    .c(_054_),
    .y(_055_)
  );
  al_ao21ttf _267_ (
    .a(L195),
    .b(_033_),
    .c(_055_),
    .y(_056_)
  );
  al_aoi21 _268_ (
    .a(L237),
    .b(_014_),
    .c(_056_),
    .y(_057_)
  );
  al_aoi21ttf _269_ (
    .a(L228),
    .b(_050_),
    .c(_057_),
    .y(_058_)
  );
  al_nand3 _270_ (
    .a(_053_),
    .b(_058_),
    .c(_052_),
    .y(L865)
  );
  al_or3fft _271_ (
    .a(L261),
    .b(_048_),
    .c(_019_),
    .y(_059_)
  );
  al_ao21ftt _272_ (
    .a(_019_),
    .b(_048_),
    .c(L261),
    .y(_060_)
  );
  al_nand3 _273_ (
    .a(L219),
    .b(_059_),
    .c(_060_),
    .y(_061_)
  );
  al_inv _274_ (
    .a(L228),
    .y(_062_)
  );
  al_nand3fft _275_ (
    .a(_062_),
    .b(_019_),
    .c(_048_),
    .y(_063_)
  );
  al_nand2 _276_ (
    .a(L255),
    .b(L267),
    .y(_064_)
  );
  al_ao21ttf _277_ (
    .a(L121),
    .b(L210),
    .c(_064_),
    .y(_065_)
  );
  al_ao21 _278_ (
    .a(L201),
    .b(_033_),
    .c(_065_),
    .y(_066_)
  );
  al_aoi21 _279_ (
    .a(L246),
    .b(_021_),
    .c(_066_),
    .y(_067_)
  );
  al_aoi21ftf _280_ (
    .a(_048_),
    .b(L237),
    .c(_067_),
    .y(_068_)
  );
  al_nand3 _281_ (
    .a(_063_),
    .b(_068_),
    .c(_061_),
    .y(L850)
  );
  al_aoi21ttf _282_ (
    .a(L59),
    .b(L156),
    .c(L447),
    .y(_069_)
  );
  al_nand3 _283_ (
    .a(L55),
    .b(L153),
    .c(_069_),
    .y(_070_)
  );
  al_nand2 _284_ (
    .a(L138),
    .b(L152),
    .y(_071_)
  );
  al_nand2ft _285_ (
    .a(L268),
    .b(L17),
    .y(_072_)
  );
  al_nand3ftt _286_ (
    .a(_072_),
    .b(L447),
    .c(_195_),
    .y(_073_)
  );
  al_and3 _287_ (
    .a(_071_),
    .b(_073_),
    .c(_070_),
    .y(_074_)
  );
  al_ao21ttf _288_ (
    .a(L106),
    .b(_194_),
    .c(_074_),
    .y(_075_)
  );
  al_and2 _289_ (
    .a(L177),
    .b(_075_),
    .y(_076_)
  );
  al_nor2 _290_ (
    .a(L177),
    .b(_075_),
    .y(_077_)
  );
  al_or2 _291_ (
    .a(_076_),
    .b(_077_),
    .y(_078_)
  );
  al_inv _292_ (
    .a(_004_),
    .y(_079_)
  );
  al_nand3fft _293_ (
    .a(_005_),
    .b(_009_),
    .c(_024_),
    .y(_080_)
  );
  al_nand3 _294_ (
    .a(L219),
    .b(_079_),
    .c(_080_),
    .y(_081_)
  );
  al_ao21 _295_ (
    .a(_062_),
    .b(_081_),
    .c(_078_),
    .y(_082_)
  );
  al_oai21 _296_ (
    .a(_076_),
    .b(_077_),
    .c(L219),
    .y(_083_)
  );
  al_ao21 _297_ (
    .a(_079_),
    .b(_080_),
    .c(_083_),
    .y(_084_)
  );
  al_nand2 _298_ (
    .a(L101),
    .b(L210),
    .y(_085_)
  );
  al_ao21ttf _299_ (
    .a(L177),
    .b(_033_),
    .c(_085_),
    .y(_086_)
  );
  al_aoi21 _300_ (
    .a(L246),
    .b(_075_),
    .c(_086_),
    .y(_087_)
  );
  al_aoi21ftf _301_ (
    .a(_028_),
    .b(_076_),
    .c(_087_),
    .y(_088_)
  );
  al_nand3 _302_ (
    .a(_088_),
    .b(_084_),
    .c(_082_),
    .y(L874)
  );
  al_nand3 _303_ (
    .a(L55),
    .b(L143),
    .c(_069_),
    .y(_089_)
  );
  al_nand2 _304_ (
    .a(L8),
    .b(L138),
    .y(_090_)
  );
  al_and3 _305_ (
    .a(_073_),
    .b(_090_),
    .c(_089_),
    .y(_091_)
  );
  al_ao21ttf _306_ (
    .a(L91),
    .b(_194_),
    .c(_091_),
    .y(_092_)
  );
  al_nand2 _307_ (
    .a(L159),
    .b(_092_),
    .y(_093_)
  );
  al_nor2 _308_ (
    .a(L159),
    .b(_092_),
    .y(_094_)
  );
  al_nand3 _309_ (
    .a(L55),
    .b(L146),
    .c(_069_),
    .y(_095_)
  );
  al_nand2 _310_ (
    .a(L51),
    .b(L138),
    .y(_096_)
  );
  al_and3 _311_ (
    .a(_073_),
    .b(_096_),
    .c(_095_),
    .y(_097_)
  );
  al_ao21ttf _312_ (
    .a(L96),
    .b(_194_),
    .c(_097_),
    .y(_098_)
  );
  al_or2 _313_ (
    .a(L165),
    .b(_098_),
    .y(_099_)
  );
  al_and2 _314_ (
    .a(L165),
    .b(_098_),
    .y(_100_)
  );
  al_nand3 _315_ (
    .a(L55),
    .b(L149),
    .c(_069_),
    .y(_101_)
  );
  al_nand2 _316_ (
    .a(L17),
    .b(L138),
    .y(_102_)
  );
  al_and3 _317_ (
    .a(_073_),
    .b(_102_),
    .c(_101_),
    .y(_103_)
  );
  al_ao21ttf _318_ (
    .a(L101),
    .b(_194_),
    .c(_103_),
    .y(_104_)
  );
  al_and2 _319_ (
    .a(L171),
    .b(_104_),
    .y(_105_)
  );
  al_nor2 _320_ (
    .a(L171),
    .b(_104_),
    .y(_106_)
  );
  al_nand3fft _321_ (
    .a(_004_),
    .b(_076_),
    .c(_080_),
    .y(_107_)
  );
  al_nand3fft _322_ (
    .a(_077_),
    .b(_106_),
    .c(_107_),
    .y(_108_)
  );
  al_nand3fft _323_ (
    .a(_100_),
    .b(_105_),
    .c(_108_),
    .y(_109_)
  );
  al_nand3ftt _324_ (
    .a(_094_),
    .b(_099_),
    .c(_109_),
    .y(_110_)
  );
  al_nand2 _325_ (
    .a(_093_),
    .b(_110_),
    .y(L866)
  );
  al_nor2ft _326_ (
    .a(_093_),
    .b(_094_),
    .y(_111_)
  );
  al_nand3 _327_ (
    .a(_099_),
    .b(_111_),
    .c(_109_),
    .y(_112_)
  );
  al_ao21 _328_ (
    .a(_099_),
    .b(_109_),
    .c(_111_),
    .y(_113_)
  );
  al_nand3 _329_ (
    .a(L219),
    .b(_112_),
    .c(_113_),
    .y(_114_)
  );
  al_nand2 _330_ (
    .a(L268),
    .b(L210),
    .y(_115_)
  );
  al_ao21ttf _331_ (
    .a(L159),
    .b(_033_),
    .c(_115_),
    .y(_116_)
  );
  al_aoi21 _332_ (
    .a(L246),
    .b(_092_),
    .c(_116_),
    .y(_117_)
  );
  al_oai21 _333_ (
    .a(_028_),
    .b(_093_),
    .c(_117_),
    .y(_118_)
  );
  al_aoi21 _334_ (
    .a(L228),
    .b(_111_),
    .c(_118_),
    .y(_119_)
  );
  al_nand2 _335_ (
    .a(_119_),
    .b(_114_),
    .y(L878)
  );
  al_inv _336_ (
    .a(_105_),
    .y(_120_)
  );
  al_nand2ft _337_ (
    .a(_100_),
    .b(_099_),
    .y(_121_)
  );
  al_ao21 _338_ (
    .a(_120_),
    .b(_108_),
    .c(_121_),
    .y(_122_)
  );
  al_nand3 _339_ (
    .a(_120_),
    .b(_121_),
    .c(_108_),
    .y(_123_)
  );
  al_nand3 _340_ (
    .a(L219),
    .b(_123_),
    .c(_122_),
    .y(_124_)
  );
  al_nand2 _341_ (
    .a(L91),
    .b(L210),
    .y(_125_)
  );
  al_ao21ttf _342_ (
    .a(L165),
    .b(_033_),
    .c(_125_),
    .y(_126_)
  );
  al_aoi21 _343_ (
    .a(L246),
    .b(_098_),
    .c(_126_),
    .y(_127_)
  );
  al_ao21ftf _344_ (
    .a(_028_),
    .b(_100_),
    .c(_127_),
    .y(_128_)
  );
  al_oa21ftf _345_ (
    .a(L228),
    .b(_121_),
    .c(_128_),
    .y(_129_)
  );
  al_nand2 _346_ (
    .a(_129_),
    .b(_124_),
    .y(L879)
  );
  al_inv _347_ (
    .a(_077_),
    .y(_130_)
  );
  al_nor2 _348_ (
    .a(_105_),
    .b(_106_),
    .y(_131_)
  );
  al_nand3 _349_ (
    .a(_130_),
    .b(_131_),
    .c(_107_),
    .y(_132_)
  );
  al_ao21 _350_ (
    .a(_130_),
    .b(_107_),
    .c(_131_),
    .y(_133_)
  );
  al_nand3 _351_ (
    .a(L219),
    .b(_132_),
    .c(_133_),
    .y(_134_)
  );
  al_nand2 _352_ (
    .a(L96),
    .b(L210),
    .y(_135_)
  );
  al_ao21ttf _353_ (
    .a(L171),
    .b(_033_),
    .c(_135_),
    .y(_136_)
  );
  al_aoi21 _354_ (
    .a(L246),
    .b(_104_),
    .c(_136_),
    .y(_137_)
  );
  al_ao21ftf _355_ (
    .a(_028_),
    .b(_105_),
    .c(_137_),
    .y(_138_)
  );
  al_aoi21 _356_ (
    .a(L228),
    .b(_131_),
    .c(_138_),
    .y(_139_)
  );
  al_nand2 _357_ (
    .a(_139_),
    .b(_134_),
    .y(L880)
  );
  al_and3 _358_ (
    .a(L42),
    .b(L29),
    .c(L36),
    .y(L390)
  );
  al_nand3 _359_ (
    .a(L59),
    .b(L80),
    .c(L75),
    .y(L420)
  );
  al_nand3 _360_ (
    .a(L59),
    .b(L80),
    .c(L36),
    .y(L421)
  );
  al_nand3 _361_ (
    .a(L59),
    .b(L42),
    .c(L36),
    .y(L422)
  );
  al_nor3fft _362_ (
    .a(L68),
    .b(L29),
    .c(_030_),
    .y(L448)
  );
  al_and3fft _363_ (
    .a(_031_),
    .b(_030_),
    .c(L74),
    .y(L449)
  );
  al_inv _364_ (
    .a(L130),
    .y(_140_)
  );
  al_nand2 _365_ (
    .a(L91),
    .b(L96),
    .y(_141_)
  );
  al_or2 _366_ (
    .a(L91),
    .b(L96),
    .y(_142_)
  );
  al_ao21 _367_ (
    .a(_142_),
    .b(_141_),
    .c(_140_),
    .y(_143_)
  );
  al_and3ftt _368_ (
    .a(L130),
    .b(_142_),
    .c(_141_),
    .y(_144_)
  );
  al_nand2ft _369_ (
    .a(_144_),
    .b(_143_),
    .y(_145_)
  );
  al_nand2ft _370_ (
    .a(L116),
    .b(L135),
    .y(_146_)
  );
  al_and2ft _371_ (
    .a(L135),
    .b(L116),
    .y(_147_)
  );
  al_nor3fft _372_ (
    .a(L111),
    .b(_146_),
    .c(_147_),
    .y(_148_)
  );
  al_oai21ftf _373_ (
    .a(_146_),
    .b(_147_),
    .c(L111),
    .y(_149_)
  );
  al_nand2ft _374_ (
    .a(_148_),
    .b(_149_),
    .y(_150_)
  );
  al_and2ft _375_ (
    .a(L106),
    .b(L101),
    .y(_151_)
  );
  al_nand2ft _376_ (
    .a(L101),
    .b(L106),
    .y(_152_)
  );
  al_nand2ft _377_ (
    .a(_151_),
    .b(_152_),
    .y(_153_)
  );
  al_and2ft _378_ (
    .a(L121),
    .b(L126),
    .y(_154_)
  );
  al_nand2ft _379_ (
    .a(L126),
    .b(L121),
    .y(_155_)
  );
  al_nand3ftt _380_ (
    .a(_154_),
    .b(_155_),
    .c(_153_),
    .y(_156_)
  );
  al_ao21ftt _381_ (
    .a(_154_),
    .b(_155_),
    .c(_153_),
    .y(_157_)
  );
  al_nand3 _382_ (
    .a(_156_),
    .b(_150_),
    .c(_157_),
    .y(_158_)
  );
  al_ao21 _383_ (
    .a(_156_),
    .b(_157_),
    .c(_150_),
    .y(_159_)
  );
  al_ao21 _384_ (
    .a(_159_),
    .b(_158_),
    .c(_145_),
    .y(_160_)
  );
  al_and3 _385_ (
    .a(_145_),
    .b(_159_),
    .c(_158_),
    .y(_161_)
  );
  al_nand2ft _386_ (
    .a(_161_),
    .b(_160_),
    .y(L767)
  );
  al_nand2 _387_ (
    .a(L159),
    .b(L165),
    .y(_162_)
  );
  al_or2 _388_ (
    .a(L159),
    .b(L165),
    .y(_163_)
  );
  al_ao21 _389_ (
    .a(_163_),
    .b(_162_),
    .c(_140_),
    .y(_164_)
  );
  al_and3ftt _390_ (
    .a(L130),
    .b(_163_),
    .c(_162_),
    .y(_165_)
  );
  al_nand2ft _391_ (
    .a(_165_),
    .b(_164_),
    .y(_166_)
  );
  al_nand2ft _392_ (
    .a(L189),
    .b(L207),
    .y(_167_)
  );
  al_and2ft _393_ (
    .a(L207),
    .b(L189),
    .y(_168_)
  );
  al_nor3fft _394_ (
    .a(L183),
    .b(_167_),
    .c(_168_),
    .y(_169_)
  );
  al_oai21ftf _395_ (
    .a(_167_),
    .b(_168_),
    .c(L183),
    .y(_170_)
  );
  al_nand2ft _396_ (
    .a(_169_),
    .b(_170_),
    .y(_171_)
  );
  al_and2ft _397_ (
    .a(L177),
    .b(L171),
    .y(_172_)
  );
  al_nand2ft _398_ (
    .a(L171),
    .b(L177),
    .y(_173_)
  );
  al_nand2ft _399_ (
    .a(_172_),
    .b(_173_),
    .y(_174_)
  );
  al_and2ft _400_ (
    .a(L195),
    .b(L201),
    .y(_175_)
  );
  al_nand2ft _401_ (
    .a(L201),
    .b(L195),
    .y(_176_)
  );
  al_nand3ftt _402_ (
    .a(_175_),
    .b(_176_),
    .c(_174_),
    .y(_177_)
  );
  al_ao21ftt _403_ (
    .a(_175_),
    .b(_176_),
    .c(_174_),
    .y(_178_)
  );
  al_nand3 _404_ (
    .a(_177_),
    .b(_171_),
    .c(_178_),
    .y(_179_)
  );
  al_ao21 _405_ (
    .a(_177_),
    .b(_178_),
    .c(_171_),
    .y(_180_)
  );
  al_ao21 _406_ (
    .a(_180_),
    .b(_179_),
    .c(_166_),
    .y(_181_)
  );
  al_and3 _407_ (
    .a(_166_),
    .b(_180_),
    .c(_179_),
    .y(_182_)
  );
  al_nand2ft _408_ (
    .a(_182_),
    .b(_181_),
    .y(L768)
  );
  al_nor3fft _409_ (
    .a(L17),
    .b(L13),
    .c(_189_),
    .y(L418)
  );
  al_and3 _410_ (
    .a(L42),
    .b(L29),
    .c(L75),
    .y(L388)
  );
  al_and3 _411_ (
    .a(L29),
    .b(L80),
    .c(L36),
    .y(L389)
  );
  al_and2 _412_ (
    .a(L85),
    .b(L86),
    .y(L391)
  );
  al_and3 _413_ (
    .a(L17),
    .b(L1),
    .c(L26),
    .y(_183_)
  );
  al_or3fft _414_ (
    .a(L13),
    .b(_183_),
    .c(L390),
    .y(L419)
  );
  al_oa21 _415_ (
    .a(L87),
    .b(L88),
    .c(L89),
    .y(L450)
  );
  al_oa21 _416_ (
    .a(L87),
    .b(L88),
    .c(L90),
    .y(L423)
  );
  al_nand3 _417_ (
    .a(L13),
    .b(L390),
    .c(_183_),
    .y(L446)
  );
  assign L273 = L390;
  assign L276 = L447;
  assign L290 = L388;
  assign L291 = L389;
  assign L292 = L390;
  assign L297 = L391;
  assign L342 = L418;
  assign L344 = L419;
  assign L351 = L420;
  assign L353 = L421;
  assign L354 = L422;
  assign L356 = L423;
  assign L369 = L268;
  assign L392 = L446;
  assign L393 = L447;
  assign L399 = L447;
  assign L401 = L448;
  assign L402 = L449;
  assign L403 = L450;
  assign L660 = L767;
  assign L661 = L768;
  assign L811 = L850;
  assign L837 = L863;
  assign L838 = L864;
  assign L839 = L865;
  assign L840 = L850;
  assign L854 = L874;
  assign L855 = L863;
  assign L856 = L864;
  assign L857 = L865;
  assign L858 = L866;
  assign L867 = L878;
  assign L868 = L879;
  assign L869 = L880;
  assign L870 = L874;
  assign L875 = L878;
  assign L876 = L879;
  assign L877 = L880;
endmodule
