
module c1908(N1, N4, N7, N10, N13, N16, N19, N22, N25, N28, N31, N34, N37, N40, N43, N46, N49, N53, N56, N60, N63, N66, N69, N72, N76, N79, N82, N85, N88, N91, N94, N99, N104, N2753, N2754, N2755, N2756, N2762, N2767, N2768, N2779, N2780, N2781, N2782, N2783, N2784, N2785, N2786, N2787, N2811, N2886, N2887, N2888, N2889, N2890, N2891, N2892, N2899);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  input N1;
  input N10;
  wire N1001;
  wire N1002;
  wire N1003;
  wire N1004;
  wire N1005;
  wire N1006;
  wire N1007;
  wire N1008;
  wire N1009;
  input N104;
  wire N1148;
  wire N1149;
  wire N1151;
  wire N1152;
  wire N1153;
  wire N1154;
  wire N1156;
  wire N1161;
  wire N1205;
  wire N1207;
  wire N1209;
  wire N1211;
  wire N1213;
  wire N1215;
  wire N1217;
  wire N1219;
  wire N1220;
  wire N1222;
  wire N1223;
  wire N1225;
  wire N1228;
  wire N1238;
  wire N1240;
  wire N1241;
  input N13;
  input N16;
  input N19;
  input N22;
  input N25;
  wire N257;
  wire N260;
  output N2753;
  output N2754;
  output N2755;
  output N2756;
  output N2762;
  output N2767;
  output N2768;
  output N2779;
  output N2780;
  output N2781;
  output N2782;
  output N2783;
  output N2784;
  output N2785;
  output N2786;
  output N2787;
  input N28;
  output N2811;
  wire N283;
  output N2886;
  output N2887;
  output N2888;
  output N2889;
  output N2890;
  output N2891;
  output N2892;
  output N2899;
  wire N297;
  wire N303;
  input N31;
  wire N316;
  wire N326;
  wire N331;
  input N34;
  wire N343;
  wire N346;
  wire N349;
  wire N352;
  wire N355;
  wire N358;
  wire N361;
  wire N364;
  wire N367;
  input N37;
  wire N370;
  wire N373;
  wire N376;
  wire N379;
  wire N382;
  wire N385;
  wire N388;
  input N4;
  input N40;
  input N43;
  input N46;
  input N49;
  input N53;
  input N56;
  input N60;
  input N63;
  input N66;
  input N69;
  input N7;
  input N72;
  input N76;
  input N79;
  input N82;
  input N85;
  input N88;
  wire N888;
  wire N889;
  wire N890;
  wire N891;
  wire N892;
  wire N894;
  wire N895;
  input N91;
  wire N913;
  wire N914;
  wire N915;
  wire N916;
  wire N917;
  wire N918;
  wire N919;
  wire N920;
  wire N938;
  input N94;
  wire N942;
  wire N946;
  wire N950;
  wire N954;
  wire N958;
  wire N968;
  wire N972;
  wire N976;
  wire N980;
  wire N984;
  wire N988;
  wire N989;
  input N99;
  wire N990;
  wire N992;
  wire N993;
  wire N997;
  al_inv _283_ (
    .a(N94),
    .y(_242_)
  );
  al_nand3ftt _284_ (
    .a(N104),
    .b(N69),
    .c(N60),
    .y(_243_)
  );
  al_nand2 _285_ (
    .a(N10),
    .b(N19),
    .y(_244_)
  );
  al_or2 _286_ (
    .a(N10),
    .b(N19),
    .y(_245_)
  );
  al_aoi21 _287_ (
    .a(_245_),
    .b(_244_),
    .c(_243_),
    .y(_246_)
  );
  al_nand3 _288_ (
    .a(_243_),
    .b(_244_),
    .c(_245_),
    .y(_247_)
  );
  al_nand2ft _289_ (
    .a(_246_),
    .b(_247_),
    .y(_248_)
  );
  al_inv _290_ (
    .a(N46),
    .y(_249_)
  );
  al_nand2ft _291_ (
    .a(N40),
    .b(N25),
    .y(_250_)
  );
  al_nand2ft _292_ (
    .a(N25),
    .b(N40),
    .y(_251_)
  );
  al_ao21 _293_ (
    .a(_250_),
    .b(_251_),
    .c(_249_),
    .y(_252_)
  );
  al_nand3ftt _294_ (
    .a(N46),
    .b(_250_),
    .c(_251_),
    .y(_253_)
  );
  al_nand2 _295_ (
    .a(N28),
    .b(N37),
    .y(_254_)
  );
  al_nor2 _296_ (
    .a(N28),
    .b(N37),
    .y(_255_)
  );
  al_nand2ft _297_ (
    .a(_255_),
    .b(_254_),
    .y(_256_)
  );
  al_nand3 _298_ (
    .a(_253_),
    .b(_252_),
    .c(_256_),
    .y(_257_)
  );
  al_ao21 _299_ (
    .a(_253_),
    .b(_252_),
    .c(_256_),
    .y(_258_)
  );
  al_ao21ttf _300_ (
    .a(_258_),
    .b(_257_),
    .c(_248_),
    .y(_259_)
  );
  al_or3fft _301_ (
    .a(_258_),
    .b(_257_),
    .c(_248_),
    .y(_260_)
  );
  al_nand3 _302_ (
    .a(_242_),
    .b(_259_),
    .c(_260_),
    .y(_261_)
  );
  al_oa21ftt _303_ (
    .a(N69),
    .b(N94),
    .c(N56),
    .y(_262_)
  );
  al_inv _304_ (
    .a(_262_),
    .y(_263_)
  );
  al_or2 _305_ (
    .a(_263_),
    .b(_261_),
    .y(_264_)
  );
  al_and2 _306_ (
    .a(_263_),
    .b(_261_),
    .y(_265_)
  );
  al_nand2ft _307_ (
    .a(_265_),
    .b(_264_),
    .y(_266_)
  );
  al_inv _308_ (
    .a(N79),
    .y(_267_)
  );
  al_inv _309_ (
    .a(N34),
    .y(_268_)
  );
  al_nand2ft _310_ (
    .a(N31),
    .b(N37),
    .y(_269_)
  );
  al_nand2ft _311_ (
    .a(N37),
    .b(N31),
    .y(_270_)
  );
  al_ao21 _312_ (
    .a(_269_),
    .b(_270_),
    .c(_268_),
    .y(_271_)
  );
  al_nand3ftt _313_ (
    .a(N34),
    .b(_269_),
    .c(_270_),
    .y(_272_)
  );
  al_nand2ft _314_ (
    .a(N43),
    .b(N28),
    .y(_273_)
  );
  al_and2ft _315_ (
    .a(N28),
    .b(N43),
    .y(_274_)
  );
  al_nor3fft _316_ (
    .a(N46),
    .b(_273_),
    .c(_274_),
    .y(_275_)
  );
  al_oai21ftf _317_ (
    .a(_273_),
    .b(_274_),
    .c(N46),
    .y(_276_)
  );
  al_nand2ft _318_ (
    .a(_275_),
    .b(_276_),
    .y(_277_)
  );
  al_nand3 _319_ (
    .a(_271_),
    .b(_272_),
    .c(_277_),
    .y(_278_)
  );
  al_nand2 _320_ (
    .a(_272_),
    .b(_271_),
    .y(_279_)
  );
  al_or3fft _321_ (
    .a(N46),
    .b(_273_),
    .c(_274_),
    .y(_280_)
  );
  al_nand3 _322_ (
    .a(_280_),
    .b(_276_),
    .c(_279_),
    .y(_281_)
  );
  al_nand2ft _323_ (
    .a(N13),
    .b(N19),
    .y(_282_)
  );
  al_nand2ft _324_ (
    .a(N19),
    .b(N13),
    .y(_000_)
  );
  al_ao21ttf _325_ (
    .a(_282_),
    .b(_000_),
    .c(N16),
    .y(_001_)
  );
  al_nand3ftt _326_ (
    .a(N16),
    .b(_282_),
    .c(_000_),
    .y(_002_)
  );
  al_nand3fft _327_ (
    .a(N72),
    .b(N104),
    .c(N49),
    .y(_003_)
  );
  al_or2 _328_ (
    .a(N1),
    .b(_003_),
    .y(_004_)
  );
  al_and2 _329_ (
    .a(N1),
    .b(_003_),
    .y(_005_)
  );
  al_nand2ft _330_ (
    .a(_005_),
    .b(_004_),
    .y(_006_)
  );
  al_ao21 _331_ (
    .a(_001_),
    .b(_002_),
    .c(_006_),
    .y(_007_)
  );
  al_and3 _332_ (
    .a(_001_),
    .b(_002_),
    .c(_006_),
    .y(_008_)
  );
  al_nand2ft _333_ (
    .a(_008_),
    .b(_007_),
    .y(_009_)
  );
  al_nand3 _334_ (
    .a(_278_),
    .b(_281_),
    .c(_009_),
    .y(_010_)
  );
  al_and3 _335_ (
    .a(_271_),
    .b(_272_),
    .c(_277_),
    .y(_011_)
  );
  al_ao21ftt _336_ (
    .a(_011_),
    .b(_281_),
    .c(_009_),
    .y(_012_)
  );
  al_nand2 _337_ (
    .a(_010_),
    .b(_012_),
    .y(_013_)
  );
  al_nand3fft _338_ (
    .a(_267_),
    .b(N94),
    .c(_013_),
    .y(_014_)
  );
  al_ao21 _339_ (
    .a(_010_),
    .b(_012_),
    .c(N94),
    .y(_015_)
  );
  al_nand2 _340_ (
    .a(_267_),
    .b(_015_),
    .y(_016_)
  );
  al_and3 _341_ (
    .a(_266_),
    .b(_016_),
    .c(_014_),
    .y(_017_)
  );
  al_oa21 _342_ (
    .a(N72),
    .b(N94),
    .c(N53),
    .y(_018_)
  );
  al_inv _343_ (
    .a(_018_),
    .y(_019_)
  );
  al_and2 _344_ (
    .a(_002_),
    .b(_001_),
    .y(_020_)
  );
  al_and2ft _345_ (
    .a(N10),
    .b(N22),
    .y(_021_)
  );
  al_nand2ft _346_ (
    .a(N22),
    .b(N10),
    .y(_022_)
  );
  al_nand2ft _347_ (
    .a(_021_),
    .b(_022_),
    .y(_023_)
  );
  al_or2 _348_ (
    .a(N4),
    .b(N7),
    .y(_024_)
  );
  al_nand2 _349_ (
    .a(N4),
    .b(N7),
    .y(_025_)
  );
  al_nand3 _350_ (
    .a(N1),
    .b(_024_),
    .c(_025_),
    .y(_026_)
  );
  al_nand2ft _351_ (
    .a(N4),
    .b(N7),
    .y(_027_)
  );
  al_nand2ft _352_ (
    .a(N7),
    .b(N4),
    .y(_028_)
  );
  al_nand3ftt _353_ (
    .a(N1),
    .b(_027_),
    .c(_028_),
    .y(_029_)
  );
  al_or3fft _354_ (
    .a(_029_),
    .b(_026_),
    .c(_023_),
    .y(_030_)
  );
  al_ao21ttf _355_ (
    .a(_029_),
    .b(_026_),
    .c(_023_),
    .y(_031_)
  );
  al_nand3 _356_ (
    .a(_031_),
    .b(_020_),
    .c(_030_),
    .y(_032_)
  );
  al_ao21 _357_ (
    .a(_031_),
    .b(_030_),
    .c(_020_),
    .y(_033_)
  );
  al_and3fft _358_ (
    .a(N104),
    .b(N25),
    .c(N63),
    .y(_034_)
  );
  al_oai21ftt _359_ (
    .a(N63),
    .b(N104),
    .c(N25),
    .y(_035_)
  );
  al_nand2ft _360_ (
    .a(_034_),
    .b(_035_),
    .y(_036_)
  );
  al_ao21 _361_ (
    .a(_280_),
    .b(_276_),
    .c(_036_),
    .y(_037_)
  );
  al_and3ftt _362_ (
    .a(_275_),
    .b(_276_),
    .c(_036_),
    .y(_038_)
  );
  al_and2ft _363_ (
    .a(_038_),
    .b(_037_),
    .y(_039_)
  );
  al_ao21 _364_ (
    .a(_033_),
    .b(_032_),
    .c(_039_),
    .y(_040_)
  );
  al_nand3 _365_ (
    .a(_033_),
    .b(_032_),
    .c(_039_),
    .y(_041_)
  );
  al_nand3 _366_ (
    .a(_242_),
    .b(_040_),
    .c(_041_),
    .y(_042_)
  );
  al_oai21 _367_ (
    .a(N72),
    .b(N94),
    .c(N49),
    .y(_043_)
  );
  al_nand2 _368_ (
    .a(_043_),
    .b(_042_),
    .y(_044_)
  );
  al_or2 _369_ (
    .a(_043_),
    .b(_042_),
    .y(_045_)
  );
  al_and3 _370_ (
    .a(_019_),
    .b(_044_),
    .c(_045_),
    .y(_046_)
  );
  al_oa21ftt _371_ (
    .a(N69),
    .b(N94),
    .c(N60),
    .y(_047_)
  );
  al_inv _372_ (
    .a(_047_),
    .y(_048_)
  );
  al_nand2ft _373_ (
    .a(_011_),
    .b(_281_),
    .y(_049_)
  );
  al_and3ftt _374_ (
    .a(N1),
    .b(_027_),
    .c(_028_),
    .y(_050_)
  );
  al_and2ft _375_ (
    .a(_050_),
    .b(_026_),
    .y(_051_)
  );
  al_inv _376_ (
    .a(N104),
    .y(_052_)
  );
  al_and2ft _377_ (
    .a(N40),
    .b(N10),
    .y(_053_)
  );
  al_nand2ft _378_ (
    .a(N10),
    .b(N40),
    .y(_054_)
  );
  al_nand2ft _379_ (
    .a(_053_),
    .b(_054_),
    .y(_055_)
  );
  al_or3fft _380_ (
    .a(_052_),
    .b(N66),
    .c(_055_),
    .y(_056_)
  );
  al_aoi21ftf _381_ (
    .a(N104),
    .b(N66),
    .c(_055_),
    .y(_057_)
  );
  al_oai21ftf _382_ (
    .a(_056_),
    .b(_057_),
    .c(_051_),
    .y(_058_)
  );
  al_nand3ftt _383_ (
    .a(_057_),
    .b(_051_),
    .c(_056_),
    .y(_059_)
  );
  al_nand3 _384_ (
    .a(_058_),
    .b(_059_),
    .c(_049_),
    .y(_060_)
  );
  al_ao21 _385_ (
    .a(_058_),
    .b(_059_),
    .c(_049_),
    .y(_061_)
  );
  al_and3 _386_ (
    .a(_242_),
    .b(_060_),
    .c(_061_),
    .y(_062_)
  );
  al_nand2 _387_ (
    .a(N76),
    .b(_062_),
    .y(_063_)
  );
  al_inv _388_ (
    .a(N76),
    .y(_064_)
  );
  al_nand3 _389_ (
    .a(_242_),
    .b(_060_),
    .c(_061_),
    .y(_065_)
  );
  al_nand2 _390_ (
    .a(_064_),
    .b(_065_),
    .y(_066_)
  );
  al_and3 _391_ (
    .a(_048_),
    .b(_066_),
    .c(_063_),
    .y(_067_)
  );
  al_and3ftt _392_ (
    .a(N104),
    .b(N69),
    .c(N56),
    .y(_068_)
  );
  al_inv _393_ (
    .a(N7),
    .y(_069_)
  );
  al_nand2ft _394_ (
    .a(N16),
    .b(N22),
    .y(_070_)
  );
  al_nand2ft _395_ (
    .a(N22),
    .b(N16),
    .y(_071_)
  );
  al_ao21 _396_ (
    .a(_070_),
    .b(_071_),
    .c(_069_),
    .y(_072_)
  );
  al_nand3ftt _397_ (
    .a(N7),
    .b(_070_),
    .c(_071_),
    .y(_073_)
  );
  al_nand3 _398_ (
    .a(_068_),
    .b(_073_),
    .c(_072_),
    .y(_074_)
  );
  al_ao21 _399_ (
    .a(_073_),
    .b(_072_),
    .c(_068_),
    .y(_075_)
  );
  al_nor3fft _400_ (
    .a(N34),
    .b(_273_),
    .c(_274_),
    .y(_076_)
  );
  al_oai21ftf _401_ (
    .a(_273_),
    .b(_274_),
    .c(N34),
    .y(_077_)
  );
  al_nand2ft _402_ (
    .a(_076_),
    .b(_077_),
    .y(_078_)
  );
  al_ao21 _403_ (
    .a(_074_),
    .b(_075_),
    .c(_078_),
    .y(_079_)
  );
  al_and3 _404_ (
    .a(_074_),
    .b(_075_),
    .c(_078_),
    .y(_080_)
  );
  al_or3fft _405_ (
    .a(_242_),
    .b(_079_),
    .c(_080_),
    .y(_081_)
  );
  al_and2 _406_ (
    .a(N85),
    .b(_081_),
    .y(_082_)
  );
  al_or2 _407_ (
    .a(N85),
    .b(_081_),
    .y(_083_)
  );
  al_and2ft _408_ (
    .a(_082_),
    .b(_083_),
    .y(_084_)
  );
  al_inv _409_ (
    .a(N82),
    .y(_085_)
  );
  al_inv _410_ (
    .a(N4),
    .y(_086_)
  );
  al_nand2ft _411_ (
    .a(N13),
    .b(N22),
    .y(_087_)
  );
  al_and2ft _412_ (
    .a(N22),
    .b(N13),
    .y(_088_)
  );
  al_oai21ftf _413_ (
    .a(_087_),
    .b(_088_),
    .c(_086_),
    .y(_089_)
  );
  al_and3fft _414_ (
    .a(N4),
    .b(_088_),
    .c(_087_),
    .y(_090_)
  );
  al_nand2ft _415_ (
    .a(_090_),
    .b(_089_),
    .y(_091_)
  );
  al_inv _416_ (
    .a(_091_),
    .y(_092_)
  );
  al_nand2 _417_ (
    .a(_253_),
    .b(_252_),
    .y(_093_)
  );
  al_and3fft _418_ (
    .a(N72),
    .b(N104),
    .c(N53),
    .y(_094_)
  );
  al_and2ft _419_ (
    .a(N43),
    .b(N31),
    .y(_095_)
  );
  al_nand2ft _420_ (
    .a(N31),
    .b(N43),
    .y(_096_)
  );
  al_nand3fft _421_ (
    .a(_094_),
    .b(_095_),
    .c(_096_),
    .y(_097_)
  );
  al_oai21ftt _422_ (
    .a(_096_),
    .b(_095_),
    .c(_094_),
    .y(_098_)
  );
  al_or3fft _423_ (
    .a(_097_),
    .b(_098_),
    .c(_093_),
    .y(_099_)
  );
  al_oai21ftf _424_ (
    .a(_096_),
    .b(_095_),
    .c(_094_),
    .y(_100_)
  );
  al_nand3ftt _425_ (
    .a(_095_),
    .b(_094_),
    .c(_096_),
    .y(_101_)
  );
  al_and3 _426_ (
    .a(_100_),
    .b(_101_),
    .c(_093_),
    .y(_102_)
  );
  al_oai21ftf _427_ (
    .a(_099_),
    .b(_102_),
    .c(_092_),
    .y(_103_)
  );
  al_nand3ftt _428_ (
    .a(_102_),
    .b(_099_),
    .c(_092_),
    .y(_104_)
  );
  al_nand3 _429_ (
    .a(_242_),
    .b(_104_),
    .c(_103_),
    .y(_105_)
  );
  al_or2 _430_ (
    .a(_085_),
    .b(_105_),
    .y(_106_)
  );
  al_and2 _431_ (
    .a(_085_),
    .b(_105_),
    .y(_107_)
  );
  al_nand2ft _432_ (
    .a(_107_),
    .b(_106_),
    .y(_108_)
  );
  al_nand2ft _433_ (
    .a(N88),
    .b(N104),
    .y(_109_)
  );
  al_aoi21ttf _434_ (
    .a(N72),
    .b(N69),
    .c(N94),
    .y(_110_)
  );
  al_nand2 _435_ (
    .a(N72),
    .b(N69),
    .y(_111_)
  );
  al_nand3ftt _436_ (
    .a(N104),
    .b(N99),
    .c(_111_),
    .y(_112_)
  );
  al_ao21ftf _437_ (
    .a(_109_),
    .b(_110_),
    .c(_112_),
    .y(_113_)
  );
  al_and3 _438_ (
    .a(_084_),
    .b(_113_),
    .c(_108_),
    .y(_114_)
  );
  al_nand3 _439_ (
    .a(_046_),
    .b(_067_),
    .c(_114_),
    .y(_115_)
  );
  al_oai21ftt _440_ (
    .a(_017_),
    .b(_115_),
    .c(N1),
    .y(_116_)
  );
  al_and3fft _441_ (
    .a(N1),
    .b(_115_),
    .c(_017_),
    .y(_117_)
  );
  al_nand2ft _442_ (
    .a(_117_),
    .b(_116_),
    .y(N2753)
  );
  al_nand3fft _443_ (
    .a(N79),
    .b(N94),
    .c(_013_),
    .y(_118_)
  );
  al_nand2 _444_ (
    .a(N79),
    .b(_015_),
    .y(_119_)
  );
  al_and3 _445_ (
    .a(_266_),
    .b(_119_),
    .c(_118_),
    .y(_120_)
  );
  al_and3 _446_ (
    .a(_046_),
    .b(_067_),
    .c(_120_),
    .y(_121_)
  );
  al_nor3fft _447_ (
    .a(_084_),
    .b(_113_),
    .c(_108_),
    .y(_122_)
  );
  al_ao21 _448_ (
    .a(_122_),
    .b(_121_),
    .c(_086_),
    .y(_123_)
  );
  al_and3 _449_ (
    .a(_086_),
    .b(_122_),
    .c(_121_),
    .y(_124_)
  );
  al_nand2ft _450_ (
    .a(_124_),
    .b(_123_),
    .y(N2754)
  );
  al_and3ftt _451_ (
    .a(_084_),
    .b(_113_),
    .c(_108_),
    .y(_125_)
  );
  al_ao21 _452_ (
    .a(_125_),
    .b(_121_),
    .c(_069_),
    .y(_126_)
  );
  al_and3 _453_ (
    .a(_069_),
    .b(_125_),
    .c(_121_),
    .y(_127_)
  );
  al_nand2ft _454_ (
    .a(_127_),
    .b(_126_),
    .y(N2755)
  );
  al_and3ftt _455_ (
    .a(_266_),
    .b(_119_),
    .c(_118_),
    .y(_128_)
  );
  al_oai21ftt _456_ (
    .a(_128_),
    .b(_115_),
    .c(N10),
    .y(_129_)
  );
  al_and3fft _457_ (
    .a(N10),
    .b(_115_),
    .c(_128_),
    .y(_130_)
  );
  al_nand2ft _458_ (
    .a(_130_),
    .b(_129_),
    .y(N2756)
  );
  al_and3ftt _459_ (
    .a(_266_),
    .b(_016_),
    .c(_014_),
    .y(_131_)
  );
  al_and3 _460_ (
    .a(_046_),
    .b(_067_),
    .c(_131_),
    .y(_132_)
  );
  al_nand2ft _461_ (
    .a(N91),
    .b(N104),
    .y(_133_)
  );
  al_ao21ftf _462_ (
    .a(_133_),
    .b(_110_),
    .c(_112_),
    .y(_134_)
  );
  al_and3ftt _463_ (
    .a(_084_),
    .b(_134_),
    .c(_108_),
    .y(_135_)
  );
  al_ao21ttf _464_ (
    .a(_135_),
    .b(_132_),
    .c(N28),
    .y(_136_)
  );
  al_and3ftt _465_ (
    .a(N28),
    .b(_135_),
    .c(_132_),
    .y(_137_)
  );
  al_nand2ft _466_ (
    .a(_137_),
    .b(_136_),
    .y(N2762)
  );
  al_and2 _467_ (
    .a(_046_),
    .b(_067_),
    .y(_138_)
  );
  al_and3fft _468_ (
    .a(_107_),
    .b(_084_),
    .c(_106_),
    .y(_139_)
  );
  al_nand3 _469_ (
    .a(_134_),
    .b(_139_),
    .c(_017_),
    .y(_140_)
  );
  al_ao21ftf _470_ (
    .a(_140_),
    .b(_138_),
    .c(N43),
    .y(_141_)
  );
  al_and3fft _471_ (
    .a(N43),
    .b(_140_),
    .c(_138_),
    .y(_142_)
  );
  al_nand2ft _472_ (
    .a(_142_),
    .b(_141_),
    .y(N2767)
  );
  al_nor3fft _473_ (
    .a(_084_),
    .b(_134_),
    .c(_108_),
    .y(_143_)
  );
  al_ao21 _474_ (
    .a(_143_),
    .b(_132_),
    .c(_249_),
    .y(_144_)
  );
  al_and3 _475_ (
    .a(_249_),
    .b(_143_),
    .c(_132_),
    .y(_145_)
  );
  al_nand2ft _476_ (
    .a(_145_),
    .b(_144_),
    .y(N2768)
  );
  al_nand2 _477_ (
    .a(N76),
    .b(_065_),
    .y(_146_)
  );
  al_nand2 _478_ (
    .a(_064_),
    .b(_062_),
    .y(_147_)
  );
  al_and3 _479_ (
    .a(_048_),
    .b(_146_),
    .c(_147_),
    .y(_148_)
  );
  al_and3 _480_ (
    .a(_046_),
    .b(_148_),
    .c(_017_),
    .y(_149_)
  );
  al_ao21ttf _481_ (
    .a(_122_),
    .b(_149_),
    .c(N13),
    .y(_150_)
  );
  al_and3ftt _482_ (
    .a(N13),
    .b(_122_),
    .c(_149_),
    .y(_151_)
  );
  al_nand2ft _483_ (
    .a(_151_),
    .b(_150_),
    .y(N2779)
  );
  al_ao21ttf _484_ (
    .a(_125_),
    .b(_149_),
    .c(N16),
    .y(_152_)
  );
  al_and3ftt _485_ (
    .a(N16),
    .b(_125_),
    .c(_149_),
    .y(_153_)
  );
  al_nand2ft _486_ (
    .a(_153_),
    .b(_152_),
    .y(N2780)
  );
  al_and2 _487_ (
    .a(_046_),
    .b(_148_),
    .y(_154_)
  );
  al_oa21ftt _488_ (
    .a(_106_),
    .b(_107_),
    .c(_084_),
    .y(_155_)
  );
  al_nand3 _489_ (
    .a(_155_),
    .b(_113_),
    .c(_131_),
    .y(_156_)
  );
  al_ao21ftf _490_ (
    .a(_156_),
    .b(_154_),
    .c(N19),
    .y(_157_)
  );
  al_and3fft _491_ (
    .a(N19),
    .b(_156_),
    .c(_154_),
    .y(_158_)
  );
  al_nand2ft _492_ (
    .a(_158_),
    .b(_157_),
    .y(N2781)
  );
  al_nand3 _493_ (
    .a(_113_),
    .b(_139_),
    .c(_120_),
    .y(_159_)
  );
  al_ao21ftf _494_ (
    .a(_159_),
    .b(_154_),
    .c(N22),
    .y(_160_)
  );
  al_and3fft _495_ (
    .a(N22),
    .b(_159_),
    .c(_154_),
    .y(_161_)
  );
  al_nand2ft _496_ (
    .a(_161_),
    .b(_160_),
    .y(N2782)
  );
  al_nand2 _497_ (
    .a(_128_),
    .b(_143_),
    .y(_162_)
  );
  al_oai21ftt _498_ (
    .a(_154_),
    .b(_162_),
    .c(N25),
    .y(_163_)
  );
  al_and3fft _499_ (
    .a(N25),
    .b(_162_),
    .c(_154_),
    .y(_164_)
  );
  al_nand2ft _500_ (
    .a(_164_),
    .b(_163_),
    .y(N2783)
  );
  al_aoi21 _501_ (
    .a(_044_),
    .b(_045_),
    .c(_018_),
    .y(_165_)
  );
  al_and3 _502_ (
    .a(_165_),
    .b(_067_),
    .c(_017_),
    .y(_166_)
  );
  al_ao21ttf _503_ (
    .a(_143_),
    .b(_166_),
    .c(N31),
    .y(_167_)
  );
  al_and3ftt _504_ (
    .a(N31),
    .b(_143_),
    .c(_166_),
    .y(_168_)
  );
  al_nand2ft _505_ (
    .a(_168_),
    .b(_167_),
    .y(N2784)
  );
  al_ao21 _506_ (
    .a(_135_),
    .b(_166_),
    .c(_268_),
    .y(_169_)
  );
  al_and3 _507_ (
    .a(_268_),
    .b(_135_),
    .c(_166_),
    .y(_170_)
  );
  al_nand2ft _508_ (
    .a(_170_),
    .b(_169_),
    .y(N2785)
  );
  al_nand2 _509_ (
    .a(_044_),
    .b(_045_),
    .y(_171_)
  );
  al_nand3 _510_ (
    .a(_019_),
    .b(_171_),
    .c(_067_),
    .y(_172_)
  );
  al_nand3 _511_ (
    .a(_155_),
    .b(_134_),
    .c(_131_),
    .y(_173_)
  );
  al_oa21 _512_ (
    .a(_172_),
    .b(_173_),
    .c(N37),
    .y(_174_)
  );
  al_or3 _513_ (
    .a(N37),
    .b(_172_),
    .c(_173_),
    .y(_175_)
  );
  al_or2ft _514_ (
    .a(_175_),
    .b(_174_),
    .y(N2786)
  );
  al_oa21 _515_ (
    .a(_172_),
    .b(_162_),
    .c(N40),
    .y(_176_)
  );
  al_or3 _516_ (
    .a(N40),
    .b(_172_),
    .c(_162_),
    .y(_177_)
  );
  al_or2ft _517_ (
    .a(_177_),
    .b(_176_),
    .y(N2787)
  );
  al_nand3 _518_ (
    .a(_017_),
    .b(_125_),
    .c(_154_),
    .y(_178_)
  );
  al_nand3 _519_ (
    .a(_017_),
    .b(_122_),
    .c(_154_),
    .y(_179_)
  );
  al_aoi21ftf _520_ (
    .a(_115_),
    .b(_128_),
    .c(_179_),
    .y(_180_)
  );
  al_and3 _521_ (
    .a(_017_),
    .b(_114_),
    .c(_138_),
    .y(_181_)
  );
  al_ao21ttf _522_ (
    .a(_159_),
    .b(_156_),
    .c(_154_),
    .y(_182_)
  );
  al_oai21 _523_ (
    .a(_122_),
    .b(_125_),
    .c(_121_),
    .y(_183_)
  );
  al_and3ftt _524_ (
    .a(_181_),
    .b(_183_),
    .c(_182_),
    .y(_184_)
  );
  al_and3 _525_ (
    .a(_178_),
    .b(_180_),
    .c(_184_),
    .y(_185_)
  );
  al_nand3 _526_ (
    .a(_128_),
    .b(_143_),
    .c(_154_),
    .y(_186_)
  );
  al_aoi21ftf _527_ (
    .a(_140_),
    .b(_138_),
    .c(_186_),
    .y(_187_)
  );
  al_ao21 _528_ (
    .a(_173_),
    .b(_162_),
    .c(_172_),
    .y(_188_)
  );
  al_nand3 _529_ (
    .a(_131_),
    .b(_135_),
    .c(_138_),
    .y(_189_)
  );
  al_and3 _530_ (
    .a(_131_),
    .b(_143_),
    .c(_138_),
    .y(_190_)
  );
  al_oai21 _531_ (
    .a(_135_),
    .b(_143_),
    .c(_166_),
    .y(_191_)
  );
  al_and3ftt _532_ (
    .a(_190_),
    .b(_189_),
    .c(_191_),
    .y(_192_)
  );
  al_and3 _533_ (
    .a(_188_),
    .b(_187_),
    .c(_192_),
    .y(_193_)
  );
  al_nand2 _534_ (
    .a(_047_),
    .b(_018_),
    .y(_194_)
  );
  al_nor2 _535_ (
    .a(_047_),
    .b(_018_),
    .y(_195_)
  );
  al_nand2ft _536_ (
    .a(_195_),
    .b(_194_),
    .y(_196_)
  );
  al_and3 _537_ (
    .a(_146_),
    .b(_147_),
    .c(_171_),
    .y(_197_)
  );
  al_aoi21ftt _538_ (
    .a(_196_),
    .b(_197_),
    .c(_154_),
    .y(_198_)
  );
  al_nand3ftt _539_ (
    .a(_112_),
    .b(_155_),
    .c(_120_),
    .y(_199_)
  );
  al_ao21 _540_ (
    .a(_172_),
    .b(_198_),
    .c(_199_),
    .y(_200_)
  );
  al_nand3 _541_ (
    .a(_200_),
    .b(_185_),
    .c(_193_),
    .y(_201_)
  );
  al_nand2 _542_ (
    .a(_155_),
    .b(_120_),
    .y(_202_)
  );
  al_nand3 _543_ (
    .a(_019_),
    .b(_171_),
    .c(_148_),
    .y(_203_)
  );
  al_or2 _544_ (
    .a(_155_),
    .b(_120_),
    .y(_204_)
  );
  al_nor2 _545_ (
    .a(_139_),
    .b(_131_),
    .y(_205_)
  );
  al_nand3ftt _546_ (
    .a(_112_),
    .b(_204_),
    .c(_205_),
    .y(_206_)
  );
  al_ao21 _547_ (
    .a(_202_),
    .b(_206_),
    .c(_203_),
    .y(_207_)
  );
  al_nand2 _548_ (
    .a(_052_),
    .b(_207_),
    .y(_208_)
  );
  al_ao21 _549_ (
    .a(N99),
    .b(_201_),
    .c(_208_),
    .y(N2811)
  );
  al_and3 _550_ (
    .a(_109_),
    .b(_033_),
    .c(_032_),
    .y(_209_)
  );
  al_or2 _551_ (
    .a(N104),
    .b(_185_),
    .y(_210_)
  );
  al_ao21ttf _552_ (
    .a(N88),
    .b(N63),
    .c(N104),
    .y(_211_)
  );
  al_ao21 _553_ (
    .a(_211_),
    .b(_210_),
    .c(_209_),
    .y(_212_)
  );
  al_and3 _554_ (
    .a(_209_),
    .b(_211_),
    .c(_210_),
    .y(_213_)
  );
  al_nand2ft _555_ (
    .a(_213_),
    .b(_212_),
    .y(N2891)
  );
  al_or2 _556_ (
    .a(N104),
    .b(_193_),
    .y(_214_)
  );
  al_ao21ttf _557_ (
    .a(N91),
    .b(N66),
    .c(N104),
    .y(_215_)
  );
  al_and2 _558_ (
    .a(_250_),
    .b(_251_),
    .y(_216_)
  );
  al_nand3 _559_ (
    .a(_216_),
    .b(_278_),
    .c(_281_),
    .y(_217_)
  );
  al_ao21 _560_ (
    .a(_278_),
    .b(_281_),
    .c(_216_),
    .y(_218_)
  );
  al_and3 _561_ (
    .a(_133_),
    .b(_217_),
    .c(_218_),
    .y(_219_)
  );
  al_and3 _562_ (
    .a(_215_),
    .b(_219_),
    .c(_214_),
    .y(_220_)
  );
  al_ao21 _563_ (
    .a(_215_),
    .b(_214_),
    .c(_219_),
    .y(_221_)
  );
  al_nand2ft _564_ (
    .a(_220_),
    .b(_221_),
    .y(N2892)
  );
  al_and2 _565_ (
    .a(_040_),
    .b(_041_),
    .y(_222_)
  );
  al_aoi21 _566_ (
    .a(_185_),
    .b(_193_),
    .c(_242_),
    .y(_223_)
  );
  al_nand3 _567_ (
    .a(N49),
    .b(_222_),
    .c(_223_),
    .y(_224_)
  );
  al_nand2ft _568_ (
    .a(N99),
    .b(N104),
    .y(_225_)
  );
  al_ao21 _569_ (
    .a(N49),
    .b(_223_),
    .c(_222_),
    .y(_226_)
  );
  al_and3 _570_ (
    .a(_225_),
    .b(_224_),
    .c(_226_),
    .y(N2886)
  );
  al_nand2 _571_ (
    .a(_060_),
    .b(_061_),
    .y(_227_)
  );
  al_nand3fft _572_ (
    .a(_064_),
    .b(_227_),
    .c(_223_),
    .y(_228_)
  );
  al_ao21ttf _573_ (
    .a(N76),
    .b(_223_),
    .c(_227_),
    .y(_229_)
  );
  al_and3 _574_ (
    .a(_225_),
    .b(_228_),
    .c(_229_),
    .y(N2887)
  );
  al_nand2 _575_ (
    .a(_104_),
    .b(_103_),
    .y(_230_)
  );
  al_nand3fft _576_ (
    .a(_085_),
    .b(_230_),
    .c(_223_),
    .y(_231_)
  );
  al_ao21ttf _577_ (
    .a(N82),
    .b(_223_),
    .c(_230_),
    .y(_232_)
  );
  al_and3 _578_ (
    .a(_225_),
    .b(_231_),
    .c(_232_),
    .y(N2888)
  );
  al_and2ft _579_ (
    .a(_080_),
    .b(_079_),
    .y(_233_)
  );
  al_nand3 _580_ (
    .a(N85),
    .b(_233_),
    .c(_223_),
    .y(_234_)
  );
  al_ao21 _581_ (
    .a(N85),
    .b(_223_),
    .c(_233_),
    .y(_235_)
  );
  al_and3 _582_ (
    .a(_225_),
    .b(_234_),
    .c(_235_),
    .y(N2889)
  );
  al_nand2 _583_ (
    .a(_259_),
    .b(_260_),
    .y(_236_)
  );
  al_inv _584_ (
    .a(_236_),
    .y(_237_)
  );
  al_nand3 _585_ (
    .a(N56),
    .b(_237_),
    .c(_223_),
    .y(_238_)
  );
  al_ao21 _586_ (
    .a(N56),
    .b(_223_),
    .c(_237_),
    .y(_239_)
  );
  al_and3 _587_ (
    .a(_225_),
    .b(_238_),
    .c(_239_),
    .y(N2890)
  );
  al_nand3 _588_ (
    .a(N79),
    .b(_013_),
    .c(_223_),
    .y(_240_)
  );
  al_ao21 _589_ (
    .a(N79),
    .b(_223_),
    .c(_013_),
    .y(_241_)
  );
  al_and3 _590_ (
    .a(_225_),
    .b(_240_),
    .c(_241_),
    .y(N2899)
  );
  assign N1001 = N25;
  assign N1002 = N16;
  assign N1003 = N22;
  assign N1004 = N7;
  assign N1005 = N28;
  assign N1006 = N43;
  assign N1007 = N34;
  assign N1008 = N19;
  assign N1009 = N28;
  assign N1148 = N1;
  assign N1149 = N1;
  assign N1151 = N13;
  assign N1152 = N13;
  assign N1153 = N28;
  assign N1154 = N28;
  assign N1156 = N31;
  assign N1161 = N46;
  assign N1205 = N4;
  assign N1207 = N4;
  assign N1209 = N16;
  assign N1211 = N16;
  assign N1213 = N43;
  assign N1215 = N43;
  assign N1217 = N25;
  assign N1219 = N25;
  assign N1220 = N34;
  assign N1222 = N31;
  assign N1223 = N34;
  assign N1225 = N40;
  assign N1228 = N40;
  assign N1238 = N40;
  assign N1240 = N46;
  assign N1241 = N40;
  assign N257 = N69;
  assign N260 = N69;
  assign N283 = N94;
  assign N297 = N94;
  assign N303 = N99;
  assign N316 = N104;
  assign N326 = N104;
  assign N331 = N104;
  assign N343 = N1;
  assign N346 = N4;
  assign N349 = N7;
  assign N352 = N10;
  assign N355 = N13;
  assign N358 = N16;
  assign N361 = N19;
  assign N364 = N22;
  assign N367 = N25;
  assign N370 = N28;
  assign N373 = N31;
  assign N376 = N34;
  assign N379 = N37;
  assign N382 = N40;
  assign N385 = N43;
  assign N388 = N46;
  assign N888 = N10;
  assign N889 = N22;
  assign N890 = N25;
  assign N891 = N40;
  assign N892 = N1;
  assign N894 = N10;
  assign N895 = N37;
  assign N913 = N76;
  assign N914 = N76;
  assign N915 = N79;
  assign N916 = N79;
  assign N917 = N82;
  assign N918 = N82;
  assign N919 = N85;
  assign N920 = N85;
  assign N938 = N7;
  assign N942 = N7;
  assign N946 = N19;
  assign N950 = N19;
  assign N954 = N46;
  assign N958 = N46;
  assign N968 = N37;
  assign N972 = N37;
  assign N976 = N10;
  assign N980 = N10;
  assign N984 = N1;
  assign N988 = N13;
  assign N989 = N22;
  assign N990 = N4;
  assign N992 = N43;
  assign N993 = N31;
  assign N997 = N25;
endmodule
