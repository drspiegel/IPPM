
module c7552(N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N242, N245, N248, N251, N254, N257, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N358, N361, N364, N367, N382, N241_I, N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884, N885, N889, N945, N1110, N1111, N1112, N1113, N1114, N1489, N1490, N1781, N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908, N11333, N11334, N11340, N11342, N241_O);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  input N1;
  input N100;
  output N10025;
  output N10101;
  output N10102;
  output N10103;
  output N10104;
  output N10109;
  output N10110;
  output N10111;
  output N10112;
  input N103;
  output N10350;
  output N10351;
  output N10352;
  output N10353;
  output N10574;
  output N10575;
  output N10576;
  input N106;
  output N10628;
  output N10632;
  output N10641;
  output N10704;
  output N10706;
  output N10711;
  output N10712;
  output N10713;
  output N10714;
  output N10715;
  output N10716;
  output N10717;
  output N10718;
  output N10729;
  output N10759;
  output N10760;
  output N10761;
  output N10762;
  output N10763;
  wire N10778;
  wire N10781;
  output N10827;
  output N10837;
  output N10838;
  output N10839;
  output N10840;
  output N10868;
  output N10869;
  output N10870;
  output N10871;
  input N109;
  output N10905;
  output N10906;
  output N10907;
  output N10908;
  input N110;
  input N111;
  output N1110;
  output N1111;
  output N1112;
  output N1113;
  output N1114;
  wire N1116;
  input N112;
  wire N1125;
  input N113;
  output N11333;
  output N11334;
  output N11340;
  output N11342;
  wire N1136;
  input N114;
  wire N1147;
  input N115;
  wire N1160;
  wire N1175;
  input N118;
  wire N1182;
  input N12;
  input N121;
  wire N1233;
  input N124;
  wire N1244;
  wire N1249;
  wire N1256;
  input N127;
  wire N1270;
  wire N1277;
  wire N1287;
  wire N1299;
  input N130;
  wire N1308;
  wire N1311;
  input N133;
  input N134;
  input N135;
  input N138;
  input N141;
  wire N1428;
  wire N1431;
  input N144;
  input N147;
  output N1489;
  output N1490;
  input N15;
  input N150;
  input N151;
  input N152;
  input N153;
  input N154;
  input N155;
  input N156;
  input N157;
  input N158;
  input N159;
  input N160;
  input N161;
  input N162;
  input N163;
  input N164;
  input N165;
  input N166;
  input N167;
  input N168;
  input N169;
  input N170;
  input N171;
  input N172;
  input N173;
  input N174;
  input N175;
  input N176;
  input N177;
  input N178;
  output N1781;
  input N179;
  input N18;
  input N180;
  input N181;
  input N182;
  wire N1828;
  wire N1829;
  input N183;
  wire N1830;
  wire N1833;
  input N184;
  wire N1840;
  wire N1841;
  wire N1842;
  wire N1843;
  input N185;
  input N186;
  wire N1867;
  wire N1868;
  wire N1869;
  input N187;
  wire N1870;
  wire N1871;
  wire N1872;
  wire N1873;
  wire N1874;
  wire N1875;
  wire N1876;
  wire N1877;
  wire N1878;
  wire N1879;
  input N188;
  wire N1880;
  wire N1881;
  wire N1882;
  wire N1883;
  wire N1884;
  input N189;
  input N190;
  input N191;
  wire N1913;
  input N192;
  input N193;
  wire N1931;
  wire N1932;
  wire N1933;
  wire N1934;
  wire N1935;
  wire N1936;
  wire N1937;
  wire N1938;
  wire N1939;
  input N194;
  wire N1940;
  wire N1941;
  wire N1942;
  wire N1943;
  wire N1944;
  wire N1945;
  wire N1946;
  input N195;
  input N196;
  wire N1968;
  wire N1969;
  input N197;
  wire N1970;
  wire N1971;
  wire N1972;
  wire N1973;
  wire N1974;
  wire N1975;
  wire N1976;
  input N198;
  input N199;
  wire N1997;
  input N200;
  input N201;
  wire N2015;
  wire N2016;
  wire N2017;
  wire N2018;
  wire N2019;
  input N202;
  wire N2020;
  wire N2021;
  wire N2022;
  wire N2023;
  input N203;
  input N204;
  input N205;
  input N206;
  input N207;
  input N208;
  input N209;
  input N210;
  input N211;
  input N212;
  input N213;
  input N214;
  input N215;
  input N216;
  input N217;
  input N218;
  input N219;
  input N220;
  input N221;
  input N222;
  input N223;
  input N224;
  input N225;
  input N226;
  wire N2267;
  input N227;
  wire N2275;
  input N228;
  wire N2287;
  input N229;
  wire N2293;
  input N23;
  input N230;
  wire N2309;
  input N231;
  wire N2315;
  input N232;
  input N233;
  wire N2331;
  input N234;
  input N235;
  input N236;
  wire N2368;
  input N237;
  input N238;
  wire N2384;
  input N239;
  wire N2390;
  input N240;
  wire N2406;
  wire N2412;
  input N241_I;
  output N241_O;
  input N242;
  input N245;
  input N248;
  input N251;
  input N254;
  input N257;
  input N26;
  input N260;
  input N263;
  input N267;
  input N271;
  input N274;
  input N277;
  input N280;
  input N283;
  input N286;
  input N289;
  input N29;
  input N293;
  input N296;
  input N299;
  input N303;
  input N307;
  input N310;
  input N313;
  input N316;
  input N319;
  input N32;
  input N322;
  input N325;
  input N328;
  input N331;
  input N334;
  input N337;
  input N340;
  input N343;
  input N346;
  input N349;
  input N35;
  input N352;
  input N355;
  input N358;
  input N361;
  input N364;
  input N367;
  input N38;
  input N382;
  output N387;
  output N388;
  input N41;
  input N44;
  input N47;
  output N478;
  output N482;
  output N484;
  output N486;
  output N489;
  output N492;
  input N5;
  input N50;
  output N501;
  output N505;
  output N507;
  output N509;
  output N511;
  output N513;
  output N515;
  output N517;
  output N519;
  input N53;
  output N535;
  output N537;
  output N539;
  input N54;
  output N541;
  output N543;
  output N545;
  output N547;
  output N549;
  input N55;
  output N551;
  output N553;
  output N556;
  output N559;
  input N56;
  output N561;
  output N563;
  output N565;
  output N567;
  output N569;
  input N57;
  output N571;
  output N573;
  input N58;
  output N582;
  input N59;
  wire N590;
  input N60;
  input N61;
  wire N614;
  input N62;
  wire N625;
  input N63;
  wire N636;
  input N64;
  output N643;
  input N65;
  wire N657;
  input N66;
  wire N676;
  wire N682;
  wire N689;
  input N69;
  input N70;
  output N707;
  input N73;
  input N74;
  input N75;
  wire N750;
  input N76;
  input N77;
  input N78;
  input N79;
  input N80;
  input N81;
  output N813;
  input N82;
  input N83;
  input N84;
  input N85;
  input N86;
  input N87;
  wire N871;
  input N88;
  output N881;
  output N882;
  output N883;
  output N884;
  output N885;
  output N889;
  input N89;
  input N9;
  input N94;
  output N945;
  input N97;
  al_or2 _0971_ (
    .a(N57),
    .b(N5),
    .y(N881)
  );
  al_and2 _0972_ (
    .a(N150),
    .b(N184),
    .y(_0270_)
  );
  al_and3 _0973_ (
    .a(N228),
    .b(N240),
    .c(_0270_),
    .y(_0271_)
  );
  al_inv _0974_ (
    .a(_0271_),
    .y(N882)
  );
  al_and2 _0975_ (
    .a(N152),
    .b(N218),
    .y(_0272_)
  );
  al_nand3 _0976_ (
    .a(N210),
    .b(N230),
    .c(_0272_),
    .y(N883)
  );
  al_and2 _0977_ (
    .a(N183),
    .b(N182),
    .y(_0273_)
  );
  al_and3 _0978_ (
    .a(N185),
    .b(N186),
    .c(_0273_),
    .y(_0274_)
  );
  al_inv _0979_ (
    .a(_0274_),
    .y(N884)
  );
  al_and2 _0980_ (
    .a(N162),
    .b(N172),
    .y(_0275_)
  );
  al_and3 _0981_ (
    .a(N188),
    .b(N199),
    .c(_0275_),
    .y(_0276_)
  );
  al_inv _0982_ (
    .a(_0276_),
    .y(N885)
  );
  al_nand2ft _0983_ (
    .a(N5),
    .b(N242),
    .y(N1110)
  );
  al_inv _0984_ (
    .a(N15),
    .y(N1111)
  );
  al_nand3ftt _0985_ (
    .a(N5),
    .b(N134),
    .c(N133),
    .y(N1113)
  );
  al_nand3fft _0986_ (
    .a(N310),
    .b(N18),
    .c(N41),
    .y(_0277_)
  );
  al_and3fft _0987_ (
    .a(N18),
    .b(N41),
    .c(N310),
    .y(_0278_)
  );
  al_nor3fft _0988_ (
    .a(N367),
    .b(_0277_),
    .c(_0278_),
    .y(_0279_)
  );
  al_oai21ftf _0989_ (
    .a(_0277_),
    .b(_0278_),
    .c(N367),
    .y(_0280_)
  );
  al_and2ft _0990_ (
    .a(_0279_),
    .b(_0280_),
    .y(N10025)
  );
  al_mux2l _0991_ (
    .a(N235),
    .b(N103),
    .s(N18),
    .y(_0281_)
  );
  al_and2ft _0992_ (
    .a(N322),
    .b(_0281_),
    .y(_0282_)
  );
  al_or2ft _0993_ (
    .a(N322),
    .b(_0281_),
    .y(_0283_)
  );
  al_mux2l _0994_ (
    .a(N236),
    .b(N23),
    .s(N18),
    .y(_0284_)
  );
  al_nor2ft _0995_ (
    .a(N319),
    .b(_0284_),
    .y(_0285_)
  );
  al_and2ft _0996_ (
    .a(N319),
    .b(_0284_),
    .y(_0286_)
  );
  al_inv _0997_ (
    .a(_0286_),
    .y(_0287_)
  );
  al_mux2l _0998_ (
    .a(N237),
    .b(N26),
    .s(N18),
    .y(_0288_)
  );
  al_nor2ft _0999_ (
    .a(N316),
    .b(_0288_),
    .y(_0289_)
  );
  al_and2ft _1000_ (
    .a(N316),
    .b(_0288_),
    .y(_0290_)
  );
  al_mux2l _1001_ (
    .a(N238),
    .b(N29),
    .s(N18),
    .y(_0291_)
  );
  al_or2ft _1002_ (
    .a(N313),
    .b(_0291_),
    .y(_0292_)
  );
  al_aoi21ftf _1003_ (
    .a(N313),
    .b(_0291_),
    .c(_0277_),
    .y(_0293_)
  );
  al_nand3ftt _1004_ (
    .a(_0278_),
    .b(_0292_),
    .c(_0293_),
    .y(_0294_)
  );
  al_or3 _1005_ (
    .a(_0289_),
    .b(_0290_),
    .c(_0294_),
    .y(_0295_)
  );
  al_or2ft _1006_ (
    .a(N316),
    .b(_0288_),
    .y(_0296_)
  );
  al_nand2ft _1007_ (
    .a(N313),
    .b(_0291_),
    .y(_0297_)
  );
  al_oai21ftf _1008_ (
    .a(N313),
    .b(_0291_),
    .c(_0277_),
    .y(_0298_)
  );
  al_nand3ftt _1009_ (
    .a(_0290_),
    .b(_0297_),
    .c(_0298_),
    .y(_0299_)
  );
  al_nand2 _1010_ (
    .a(_0296_),
    .b(_0299_),
    .y(_0300_)
  );
  al_oai21ftt _1011_ (
    .a(N367),
    .b(_0295_),
    .c(_0300_),
    .y(_0301_)
  );
  al_oa21ftf _1012_ (
    .a(_0287_),
    .b(_0301_),
    .c(_0285_),
    .y(_0302_)
  );
  al_or3ftt _1013_ (
    .a(_0283_),
    .b(_0282_),
    .c(_0302_),
    .y(_0303_)
  );
  al_nand2ft _1014_ (
    .a(_0282_),
    .b(_0283_),
    .y(_0304_)
  );
  al_and2 _1015_ (
    .a(_0304_),
    .b(_0302_),
    .y(_0305_)
  );
  al_nand2ft _1016_ (
    .a(_0305_),
    .b(_0303_),
    .y(N10109)
  );
  al_or2ft _1017_ (
    .a(N319),
    .b(_0284_),
    .y(_0306_)
  );
  al_and2ft _1018_ (
    .a(_0286_),
    .b(_0306_),
    .y(_0307_)
  );
  al_and2ft _1019_ (
    .a(_0307_),
    .b(_0301_),
    .y(_0308_)
  );
  al_or3fft _1020_ (
    .a(_0306_),
    .b(_0287_),
    .c(_0301_),
    .y(_0309_)
  );
  al_nand2ft _1021_ (
    .a(_0308_),
    .b(_0309_),
    .y(N10110)
  );
  al_aoi21ftf _1022_ (
    .a(_0279_),
    .b(_0293_),
    .c(_0292_),
    .y(_0310_)
  );
  al_aoi21ftf _1023_ (
    .a(_0290_),
    .b(_0296_),
    .c(_0310_),
    .y(_0311_)
  );
  al_or3 _1024_ (
    .a(_0289_),
    .b(_0290_),
    .c(_0310_),
    .y(_0312_)
  );
  al_nand2ft _1025_ (
    .a(_0311_),
    .b(_0312_),
    .y(N10111)
  );
  al_oa21ftt _1026_ (
    .a(N367),
    .b(_0278_),
    .c(_0277_),
    .y(_0313_)
  );
  al_and3 _1027_ (
    .a(_0297_),
    .b(_0292_),
    .c(_0313_),
    .y(_0314_)
  );
  al_ao21 _1028_ (
    .a(_0292_),
    .b(_0297_),
    .c(_0313_),
    .y(_0315_)
  );
  al_nand2ft _1029_ (
    .a(_0314_),
    .b(_0315_),
    .y(N10112)
  );
  al_mux2l _1030_ (
    .a(N232),
    .b(N124),
    .s(N18),
    .y(_0316_)
  );
  al_mux2l _1031_ (
    .a(N229),
    .b(N41),
    .s(N18),
    .y(_0317_)
  );
  al_and2ft _1032_ (
    .a(_0316_),
    .b(_0317_),
    .y(_0318_)
  );
  al_nand2ft _1033_ (
    .a(_0317_),
    .b(_0316_),
    .y(_0319_)
  );
  al_mux2l _1034_ (
    .a(N231),
    .b(N100),
    .s(N18),
    .y(_0320_)
  );
  al_and2ft _1035_ (
    .a(_0284_),
    .b(_0320_),
    .y(_0321_)
  );
  al_nand2ft _1036_ (
    .a(_0320_),
    .b(_0284_),
    .y(_0322_)
  );
  al_nand2ft _1037_ (
    .a(_0321_),
    .b(_0322_),
    .y(_0323_)
  );
  al_and3ftt _1038_ (
    .a(_0318_),
    .b(_0319_),
    .c(_0323_),
    .y(_0324_)
  );
  al_ao21ftt _1039_ (
    .a(_0318_),
    .b(_0319_),
    .c(_0323_),
    .y(_0325_)
  );
  al_nand2ft _1040_ (
    .a(_0324_),
    .b(_0325_),
    .y(_0326_)
  );
  al_nor2 _1041_ (
    .a(_0281_),
    .b(_0288_),
    .y(_0327_)
  );
  al_nand2 _1042_ (
    .a(_0281_),
    .b(_0288_),
    .y(_0328_)
  );
  al_nand2ft _1043_ (
    .a(_0327_),
    .b(_0328_),
    .y(_0329_)
  );
  al_mux2l _1044_ (
    .a(N234),
    .b(N130),
    .s(N18),
    .y(_0330_)
  );
  al_mux2l _1045_ (
    .a(N233),
    .b(N127),
    .s(N18),
    .y(_0331_)
  );
  al_nor2 _1046_ (
    .a(_0330_),
    .b(_0331_),
    .y(_0332_)
  );
  al_nand2 _1047_ (
    .a(_0330_),
    .b(_0331_),
    .y(_0333_)
  );
  al_mux2l _1048_ (
    .a(N239),
    .b(N44),
    .s(N18),
    .y(_0334_)
  );
  al_nor2 _1049_ (
    .a(_0291_),
    .b(_0334_),
    .y(_0335_)
  );
  al_nand2 _1050_ (
    .a(_0291_),
    .b(_0334_),
    .y(_0336_)
  );
  al_nand2ft _1051_ (
    .a(_0335_),
    .b(_0336_),
    .y(_0337_)
  );
  al_nand3ftt _1052_ (
    .a(_0332_),
    .b(_0333_),
    .c(_0337_),
    .y(_0338_)
  );
  al_ao21ftt _1053_ (
    .a(_0332_),
    .b(_0333_),
    .c(_0337_),
    .y(_0339_)
  );
  al_nand3 _1054_ (
    .a(_0329_),
    .b(_0338_),
    .c(_0339_),
    .y(_0340_)
  );
  al_ao21 _1055_ (
    .a(_0338_),
    .b(_0339_),
    .c(_0329_),
    .y(_0341_)
  );
  al_or3fft _1056_ (
    .a(_0340_),
    .b(_0341_),
    .c(_0326_),
    .y(_0342_)
  );
  al_aoi21ttf _1057_ (
    .a(_0340_),
    .b(_0341_),
    .c(_0326_),
    .y(_0343_)
  );
  al_nand2ft _1058_ (
    .a(_0343_),
    .b(_0342_),
    .y(_0344_)
  );
  al_nand2ft _1059_ (
    .a(N156),
    .b(N18),
    .y(_0345_)
  );
  al_nand2 _1060_ (
    .a(N12),
    .b(N9),
    .y(_0346_)
  );
  al_nand2ft _1061_ (
    .a(N155),
    .b(N18),
    .y(_0347_)
  );
  al_nand3ftt _1062_ (
    .a(_0347_),
    .b(_0346_),
    .c(_0345_),
    .y(_0348_)
  );
  al_aoi21ttf _1063_ (
    .a(N12),
    .b(N9),
    .c(_0347_),
    .y(_0349_)
  );
  al_ao21ftf _1064_ (
    .a(_0345_),
    .b(_0349_),
    .c(_0348_),
    .y(_0350_)
  );
  al_nand2ft _1065_ (
    .a(N154),
    .b(N18),
    .y(_0351_)
  );
  al_aoi21ttf _1066_ (
    .a(N12),
    .b(N9),
    .c(_0351_),
    .y(_0352_)
  );
  al_nand2ft _1067_ (
    .a(N153),
    .b(N18),
    .y(_0353_)
  );
  al_nand3ftt _1068_ (
    .a(_0351_),
    .b(_0346_),
    .c(_0353_),
    .y(_0354_)
  );
  al_ao21ftf _1069_ (
    .a(_0353_),
    .b(_0352_),
    .c(_0354_),
    .y(_0355_)
  );
  al_mux2l _1070_ (
    .a(N161),
    .b(N141),
    .s(N18),
    .y(_0356_)
  );
  al_mux2l _1071_ (
    .a(N151),
    .b(N147),
    .s(N18),
    .y(_0357_)
  );
  al_and2ft _1072_ (
    .a(_0357_),
    .b(_0356_),
    .y(_0358_)
  );
  al_nand2ft _1073_ (
    .a(_0356_),
    .b(_0357_),
    .y(_0359_)
  );
  al_nand3ftt _1074_ (
    .a(_0358_),
    .b(_0359_),
    .c(_0355_),
    .y(_0360_)
  );
  al_ao21ftt _1075_ (
    .a(_0358_),
    .b(_0359_),
    .c(_0355_),
    .y(_0361_)
  );
  al_aoi21 _1076_ (
    .a(_0360_),
    .b(_0361_),
    .c(_0350_),
    .y(_0362_)
  );
  al_and3 _1077_ (
    .a(_0350_),
    .b(_0360_),
    .c(_0361_),
    .y(_0363_)
  );
  al_mux2l _1078_ (
    .a(N158),
    .b(N135),
    .s(N18),
    .y(_0364_)
  );
  al_aoi21ftf _1079_ (
    .a(N157),
    .b(N18),
    .c(_0346_),
    .y(_0365_)
  );
  al_nor2 _1080_ (
    .a(_0364_),
    .b(_0365_),
    .y(_0366_)
  );
  al_nand2 _1081_ (
    .a(_0364_),
    .b(_0365_),
    .y(_0367_)
  );
  al_mux2l _1082_ (
    .a(N160),
    .b(N138),
    .s(N18),
    .y(_0368_)
  );
  al_mux2l _1083_ (
    .a(N159),
    .b(N144),
    .s(N18),
    .y(_0369_)
  );
  al_nand2 _1084_ (
    .a(_0368_),
    .b(_0369_),
    .y(_0370_)
  );
  al_nor2 _1085_ (
    .a(_0368_),
    .b(_0369_),
    .y(_0371_)
  );
  al_nand2ft _1086_ (
    .a(_0371_),
    .b(_0370_),
    .y(_0372_)
  );
  al_ao21ftt _1087_ (
    .a(_0366_),
    .b(_0367_),
    .c(_0372_),
    .y(_0373_)
  );
  al_and3ftt _1088_ (
    .a(_0366_),
    .b(_0367_),
    .c(_0372_),
    .y(_0374_)
  );
  al_and2ft _1089_ (
    .a(_0374_),
    .b(_0373_),
    .y(_0375_)
  );
  al_nand3fft _1090_ (
    .a(_0362_),
    .b(_0363_),
    .c(_0375_),
    .y(_0376_)
  );
  al_nand2ft _1091_ (
    .a(N209),
    .b(N18),
    .y(_0377_)
  );
  al_nand2ft _1092_ (
    .a(N214),
    .b(N18),
    .y(_0378_)
  );
  al_aoi21ttf _1093_ (
    .a(N12),
    .b(N9),
    .c(_0378_),
    .y(_0379_)
  );
  al_nand2ft _1094_ (
    .a(N213),
    .b(N18),
    .y(_0380_)
  );
  al_nand3ftt _1095_ (
    .a(_0378_),
    .b(_0346_),
    .c(_0380_),
    .y(_0381_)
  );
  al_aoi21ftf _1096_ (
    .a(_0380_),
    .b(_0379_),
    .c(_0381_),
    .y(_0382_)
  );
  al_ao21ftt _1097_ (
    .a(_0377_),
    .b(_0346_),
    .c(_0382_),
    .y(_0383_)
  );
  al_and3ftt _1098_ (
    .a(_0377_),
    .b(_0346_),
    .c(_0382_),
    .y(_0384_)
  );
  al_nand2ft _1099_ (
    .a(_0384_),
    .b(_0383_),
    .y(_0385_)
  );
  al_nand2ft _1100_ (
    .a(N216),
    .b(N18),
    .y(_0386_)
  );
  al_aoi21ttf _1101_ (
    .a(N12),
    .b(N9),
    .c(_0386_),
    .y(_0387_)
  );
  al_nand2ft _1102_ (
    .a(N215),
    .b(N18),
    .y(_0388_)
  );
  al_nand3ftt _1103_ (
    .a(_0386_),
    .b(_0346_),
    .c(_0388_),
    .y(_0389_)
  );
  al_ao21ftf _1104_ (
    .a(_0388_),
    .b(_0387_),
    .c(_0389_),
    .y(_0390_)
  );
  al_ao21ttf _1105_ (
    .a(N12),
    .b(N9),
    .c(N18),
    .y(_0391_)
  );
  al_aoi21 _1106_ (
    .a(N212),
    .b(N211),
    .c(_0391_),
    .y(_0392_)
  );
  al_oai21 _1107_ (
    .a(N212),
    .b(N211),
    .c(_0392_),
    .y(_0393_)
  );
  al_or2ft _1108_ (
    .a(_0393_),
    .b(_0390_),
    .y(_0394_)
  );
  al_nand2ft _1109_ (
    .a(_0393_),
    .b(_0390_),
    .y(_0395_)
  );
  al_ao21 _1110_ (
    .a(_0394_),
    .b(_0395_),
    .c(_0385_),
    .y(_0396_)
  );
  al_and3 _1111_ (
    .a(_0394_),
    .b(_0395_),
    .c(_0385_),
    .y(_0397_)
  );
  al_oai21ttf _1112_ (
    .a(_0362_),
    .b(_0363_),
    .c(_0375_),
    .y(_0398_)
  );
  al_aoi21ftf _1113_ (
    .a(_0397_),
    .b(_0396_),
    .c(_0398_),
    .y(_0399_)
  );
  al_mux2l _1114_ (
    .a(N224),
    .b(N121),
    .s(N18),
    .y(_0400_)
  );
  al_mux2l _1115_ (
    .a(N223),
    .b(N47),
    .s(N18),
    .y(_0401_)
  );
  al_and2ft _1116_ (
    .a(_0400_),
    .b(_0401_),
    .y(_0402_)
  );
  al_nand2ft _1117_ (
    .a(_0401_),
    .b(_0400_),
    .y(_0403_)
  );
  al_nand2ft _1118_ (
    .a(_0402_),
    .b(_0403_),
    .y(_0404_)
  );
  al_mux2l _1119_ (
    .a(N226),
    .b(N97),
    .s(N18),
    .y(_0405_)
  );
  al_mux2l _1120_ (
    .a(N225),
    .b(N94),
    .s(N18),
    .y(_0406_)
  );
  al_nand2 _1121_ (
    .a(_0405_),
    .b(_0406_),
    .y(_0407_)
  );
  al_nor2 _1122_ (
    .a(_0405_),
    .b(_0406_),
    .y(_0408_)
  );
  al_and3ftt _1123_ (
    .a(_0408_),
    .b(_0407_),
    .c(_0404_),
    .y(_0409_)
  );
  al_ao21ftt _1124_ (
    .a(_0408_),
    .b(_0407_),
    .c(_0404_),
    .y(_0410_)
  );
  al_nand2ft _1125_ (
    .a(_0409_),
    .b(_0410_),
    .y(_0411_)
  );
  al_mux2l _1126_ (
    .a(N227),
    .b(N115),
    .s(N18),
    .y(_0412_)
  );
  al_mux2l _1127_ (
    .a(N217),
    .b(N118),
    .s(N18),
    .y(_0413_)
  );
  al_and2ft _1128_ (
    .a(_0412_),
    .b(_0413_),
    .y(_0414_)
  );
  al_nand2ft _1129_ (
    .a(_0413_),
    .b(_0412_),
    .y(_0415_)
  );
  al_nand2ft _1130_ (
    .a(_0414_),
    .b(_0415_),
    .y(_0416_)
  );
  al_mux2l _1131_ (
    .a(N220),
    .b(N50),
    .s(N18),
    .y(_0417_)
  );
  al_mux2l _1132_ (
    .a(N219),
    .b(N66),
    .s(N18),
    .y(_0418_)
  );
  al_nor2 _1133_ (
    .a(_0417_),
    .b(_0418_),
    .y(_0419_)
  );
  al_nand2 _1134_ (
    .a(_0417_),
    .b(_0418_),
    .y(_0420_)
  );
  al_mux2l _1135_ (
    .a(N222),
    .b(N35),
    .s(N18),
    .y(_0421_)
  );
  al_mux2l _1136_ (
    .a(N221),
    .b(N32),
    .s(N18),
    .y(_0422_)
  );
  al_nand2 _1137_ (
    .a(_0421_),
    .b(_0422_),
    .y(_0423_)
  );
  al_nor2 _1138_ (
    .a(_0421_),
    .b(_0422_),
    .y(_0424_)
  );
  al_nand2ft _1139_ (
    .a(_0424_),
    .b(_0423_),
    .y(_0425_)
  );
  al_ao21ftt _1140_ (
    .a(_0419_),
    .b(_0420_),
    .c(_0425_),
    .y(_0426_)
  );
  al_nand3ftt _1141_ (
    .a(_0419_),
    .b(_0420_),
    .c(_0425_),
    .y(_0427_)
  );
  al_ao21ttf _1142_ (
    .a(_0427_),
    .b(_0426_),
    .c(_0416_),
    .y(_0428_)
  );
  al_nand3ftt _1143_ (
    .a(_0416_),
    .b(_0427_),
    .c(_0426_),
    .y(_0429_)
  );
  al_aoi21 _1144_ (
    .a(_0429_),
    .b(_0428_),
    .c(_0411_),
    .y(_0430_)
  );
  al_nand3 _1145_ (
    .a(_0429_),
    .b(_0428_),
    .c(_0411_),
    .y(_0431_)
  );
  al_nand2ft _1146_ (
    .a(_0430_),
    .b(_0431_),
    .y(_0432_)
  );
  al_and3 _1147_ (
    .a(_0376_),
    .b(_0399_),
    .c(_0432_),
    .y(_0433_)
  );
  al_nand2 _1148_ (
    .a(_0344_),
    .b(_0433_),
    .y(N10574)
  );
  al_nand2ft _1149_ (
    .a(N18),
    .b(N76),
    .y(_0434_)
  );
  al_ao21ftf _1150_ (
    .a(N316),
    .b(N18),
    .c(_0434_),
    .y(_0435_)
  );
  al_or2 _1151_ (
    .a(N18),
    .b(N70),
    .y(_0436_)
  );
  al_ao21ttf _1152_ (
    .a(N310),
    .b(N18),
    .c(_0436_),
    .y(_0437_)
  );
  al_nand2ft _1153_ (
    .a(N18),
    .b(N69),
    .y(_0438_)
  );
  al_ao21ftf _1154_ (
    .a(N307),
    .b(N18),
    .c(_0438_),
    .y(_0439_)
  );
  al_nand2ft _1155_ (
    .a(_0437_),
    .b(_0439_),
    .y(_0440_)
  );
  al_and2ft _1156_ (
    .a(_0439_),
    .b(_0437_),
    .y(_0441_)
  );
  al_nand2ft _1157_ (
    .a(N18),
    .b(N74),
    .y(_0442_)
  );
  al_ao21ftf _1158_ (
    .a(N313),
    .b(N18),
    .c(_0442_),
    .y(_0443_)
  );
  al_nor3fft _1159_ (
    .a(_0443_),
    .b(_0440_),
    .c(_0441_),
    .y(_0444_)
  );
  al_oai21ftf _1160_ (
    .a(_0440_),
    .b(_0441_),
    .c(_0443_),
    .y(_0445_)
  );
  al_nor3fft _1161_ (
    .a(_0435_),
    .b(_0445_),
    .c(_0444_),
    .y(_0446_)
  );
  al_ao21ftt _1162_ (
    .a(_0444_),
    .b(_0445_),
    .c(_0435_),
    .y(_0447_)
  );
  al_nand2ft _1163_ (
    .a(_0446_),
    .b(_0447_),
    .y(_0448_)
  );
  al_nand2ft _1164_ (
    .a(N18),
    .b(N55),
    .y(_0449_)
  );
  al_ao21ftf _1165_ (
    .a(N331),
    .b(N18),
    .c(_0449_),
    .y(_0450_)
  );
  al_nand2ft _1166_ (
    .a(N18),
    .b(N56),
    .y(_0451_)
  );
  al_ao21ftf _1167_ (
    .a(N334),
    .b(N18),
    .c(_0451_),
    .y(_0452_)
  );
  al_nand2ft _1168_ (
    .a(_0450_),
    .b(_0452_),
    .y(_0453_)
  );
  al_and2ft _1169_ (
    .a(_0452_),
    .b(_0450_),
    .y(_0454_)
  );
  al_or2 _1170_ (
    .a(N18),
    .b(N54),
    .y(_0455_)
  );
  al_ao21ttf _1171_ (
    .a(N328),
    .b(N18),
    .c(_0455_),
    .y(_0456_)
  );
  al_and3fft _1172_ (
    .a(_0456_),
    .b(_0454_),
    .c(_0453_),
    .y(_0457_)
  );
  al_oai21ftt _1173_ (
    .a(_0453_),
    .b(_0454_),
    .c(_0456_),
    .y(_0458_)
  );
  al_nand2ft _1174_ (
    .a(_0457_),
    .b(_0458_),
    .y(_0459_)
  );
  al_nand2ft _1175_ (
    .a(N18),
    .b(N53),
    .y(_0460_)
  );
  al_ao21ftf _1176_ (
    .a(N325),
    .b(N18),
    .c(_0460_),
    .y(_0461_)
  );
  al_nand2ft _1177_ (
    .a(N18),
    .b(N75),
    .y(_0462_)
  );
  al_ao21ftf _1178_ (
    .a(N319),
    .b(N18),
    .c(_0462_),
    .y(_0463_)
  );
  al_nand2ft _1179_ (
    .a(N18),
    .b(N73),
    .y(_0464_)
  );
  al_ao21ftf _1180_ (
    .a(N322),
    .b(N18),
    .c(_0464_),
    .y(_0465_)
  );
  al_nand2ft _1181_ (
    .a(_0465_),
    .b(_0463_),
    .y(_0466_)
  );
  al_nand2ft _1182_ (
    .a(_0463_),
    .b(_0465_),
    .y(_0467_)
  );
  al_aoi21 _1183_ (
    .a(_0466_),
    .b(_0467_),
    .c(_0461_),
    .y(_0468_)
  );
  al_nand3 _1184_ (
    .a(_0461_),
    .b(_0466_),
    .c(_0467_),
    .y(_0469_)
  );
  al_or3ftt _1185_ (
    .a(_0469_),
    .b(_0468_),
    .c(_0459_),
    .y(_0470_)
  );
  al_ao21ftf _1186_ (
    .a(_0468_),
    .b(_0469_),
    .c(_0459_),
    .y(_0471_)
  );
  al_or3fft _1187_ (
    .a(_0471_),
    .b(_0470_),
    .c(_0448_),
    .y(_0472_)
  );
  al_nand2ft _1188_ (
    .a(N18),
    .b(N85),
    .y(_0473_)
  );
  al_ao21ftf _1189_ (
    .a(N286),
    .b(N18),
    .c(_0473_),
    .y(_0474_)
  );
  al_or2 _1190_ (
    .a(N18),
    .b(N64),
    .y(_0475_)
  );
  al_ao21ttf _1191_ (
    .a(N289),
    .b(N18),
    .c(_0475_),
    .y(_0476_)
  );
  al_nand2ft _1192_ (
    .a(_0476_),
    .b(_0474_),
    .y(_0477_)
  );
  al_and2ft _1193_ (
    .a(_0474_),
    .b(_0476_),
    .y(_0478_)
  );
  al_nand2ft _1194_ (
    .a(_0478_),
    .b(_0477_),
    .y(_0479_)
  );
  al_inv _1195_ (
    .a(N299),
    .y(_0480_)
  );
  al_mux2h _1196_ (
    .a(N109),
    .b(_0480_),
    .s(N18),
    .y(_0481_)
  );
  al_inv _1197_ (
    .a(N303),
    .y(_0482_)
  );
  al_mux2h _1198_ (
    .a(N110),
    .b(_0482_),
    .s(N18),
    .y(_0483_)
  );
  al_nor2 _1199_ (
    .a(_0481_),
    .b(_0483_),
    .y(_0484_)
  );
  al_nand2 _1200_ (
    .a(_0481_),
    .b(_0483_),
    .y(_0485_)
  );
  al_and3ftt _1201_ (
    .a(_0484_),
    .b(_0485_),
    .c(_0479_),
    .y(_0486_)
  );
  al_ao21ftt _1202_ (
    .a(_0484_),
    .b(_0485_),
    .c(_0479_),
    .y(_0487_)
  );
  al_nand2ft _1203_ (
    .a(_0486_),
    .b(_0487_),
    .y(_0488_)
  );
  al_nand2ft _1204_ (
    .a(N18),
    .b(N82),
    .y(_0489_)
  );
  al_ao21ftf _1205_ (
    .a(N274),
    .b(N18),
    .c(_0489_),
    .y(_0490_)
  );
  al_nand2ft _1206_ (
    .a(N18),
    .b(N65),
    .y(_0491_)
  );
  al_ao21ftf _1207_ (
    .a(N277),
    .b(N18),
    .c(_0491_),
    .y(_0492_)
  );
  al_nand2 _1208_ (
    .a(_0490_),
    .b(_0492_),
    .y(_0493_)
  );
  al_nor2 _1209_ (
    .a(_0490_),
    .b(_0492_),
    .y(_0494_)
  );
  al_nand2ft _1210_ (
    .a(N18),
    .b(N84),
    .y(_0495_)
  );
  al_ao21ftf _1211_ (
    .a(N283),
    .b(N18),
    .c(_0495_),
    .y(_0496_)
  );
  al_oai21ftf _1212_ (
    .a(_0493_),
    .b(_0494_),
    .c(_0496_),
    .y(_0497_)
  );
  al_nor3fft _1213_ (
    .a(_0496_),
    .b(_0493_),
    .c(_0494_),
    .y(_0498_)
  );
  al_nand2ft _1214_ (
    .a(_0498_),
    .b(_0497_),
    .y(_0499_)
  );
  al_inv _1215_ (
    .a(N293),
    .y(_0500_)
  );
  al_mux2h _1216_ (
    .a(N63),
    .b(_0500_),
    .s(N18),
    .y(_0501_)
  );
  al_inv _1217_ (
    .a(N296),
    .y(_0502_)
  );
  al_mux2h _1218_ (
    .a(N86),
    .b(_0502_),
    .s(N18),
    .y(_0503_)
  );
  al_nand2 _1219_ (
    .a(_0501_),
    .b(_0503_),
    .y(_0504_)
  );
  al_nor2 _1220_ (
    .a(_0501_),
    .b(_0503_),
    .y(_0505_)
  );
  al_or2 _1221_ (
    .a(N18),
    .b(N83),
    .y(_0506_)
  );
  al_ao21ttf _1222_ (
    .a(N280),
    .b(N18),
    .c(_0506_),
    .y(_0507_)
  );
  al_and3fft _1223_ (
    .a(_0507_),
    .b(_0505_),
    .c(_0504_),
    .y(_0508_)
  );
  al_oai21ftt _1224_ (
    .a(_0504_),
    .b(_0505_),
    .c(_0507_),
    .y(_0509_)
  );
  al_or3ftt _1225_ (
    .a(_0509_),
    .b(_0508_),
    .c(_0499_),
    .y(_0510_)
  );
  al_ao21ftf _1226_ (
    .a(_0508_),
    .b(_0509_),
    .c(_0499_),
    .y(_0511_)
  );
  al_nand3 _1227_ (
    .a(_0511_),
    .b(_0488_),
    .c(_0510_),
    .y(_0512_)
  );
  al_aoi21ttf _1228_ (
    .a(_0471_),
    .b(_0470_),
    .c(_0448_),
    .y(_0513_)
  );
  al_and3ftt _1229_ (
    .a(_0513_),
    .b(_0472_),
    .c(_0512_),
    .y(_0514_)
  );
  al_nand2ft _1230_ (
    .a(N18),
    .b(N81),
    .y(_0515_)
  );
  al_ao21ftf _1231_ (
    .a(N349),
    .b(N18),
    .c(_0515_),
    .y(_0516_)
  );
  al_nand2ft _1232_ (
    .a(N18),
    .b(N80),
    .y(_0517_)
  );
  al_ao21ftf _1233_ (
    .a(N352),
    .b(N18),
    .c(_0517_),
    .y(_0518_)
  );
  al_and2ft _1234_ (
    .a(_0518_),
    .b(_0516_),
    .y(_0519_)
  );
  al_and2ft _1235_ (
    .a(_0516_),
    .b(_0518_),
    .y(_0520_)
  );
  al_nand2ft _1236_ (
    .a(N18),
    .b(N61),
    .y(_0521_)
  );
  al_ao21ftf _1237_ (
    .a(N361),
    .b(N18),
    .c(_0521_),
    .y(_0522_)
  );
  al_nand2ft _1238_ (
    .a(N18),
    .b(N62),
    .y(_0523_)
  );
  al_ao21ftf _1239_ (
    .a(N364),
    .b(N18),
    .c(_0523_),
    .y(_0524_)
  );
  al_and2ft _1240_ (
    .a(_0522_),
    .b(_0524_),
    .y(_0525_)
  );
  al_nand2ft _1241_ (
    .a(_0524_),
    .b(_0522_),
    .y(_0526_)
  );
  al_nand2ft _1242_ (
    .a(_0525_),
    .b(_0526_),
    .y(_0527_)
  );
  al_nand3fft _1243_ (
    .a(_0519_),
    .b(_0520_),
    .c(_0527_),
    .y(_0528_)
  );
  al_oai21ttf _1244_ (
    .a(_0519_),
    .b(_0520_),
    .c(_0527_),
    .y(_0529_)
  );
  al_nand2ft _1245_ (
    .a(N18),
    .b(N78),
    .y(_0530_)
  );
  al_ao21ftf _1246_ (
    .a(N343),
    .b(N18),
    .c(_0530_),
    .y(_0531_)
  );
  al_nand2ft _1247_ (
    .a(N18),
    .b(N59),
    .y(_0532_)
  );
  al_ao21ftf _1248_ (
    .a(N346),
    .b(N18),
    .c(_0532_),
    .y(_0533_)
  );
  al_and2ft _1249_ (
    .a(_0531_),
    .b(_0533_),
    .y(_0534_)
  );
  al_nand2ft _1250_ (
    .a(_0533_),
    .b(_0531_),
    .y(_0535_)
  );
  al_nand2ft _1251_ (
    .a(_0534_),
    .b(_0535_),
    .y(_0536_)
  );
  al_ao21ttf _1252_ (
    .a(_0528_),
    .b(_0529_),
    .c(_0536_),
    .y(_0537_)
  );
  al_nand3ftt _1253_ (
    .a(_0536_),
    .b(_0528_),
    .c(_0529_),
    .y(_0538_)
  );
  al_nand2ft _1254_ (
    .a(N18),
    .b(N79),
    .y(_0539_)
  );
  al_ao21ftf _1255_ (
    .a(N355),
    .b(N18),
    .c(_0539_),
    .y(_0540_)
  );
  al_or2 _1256_ (
    .a(N18),
    .b(N60),
    .y(_0541_)
  );
  al_ao21ttf _1257_ (
    .a(N358),
    .b(N18),
    .c(_0541_),
    .y(_0542_)
  );
  al_nor2 _1258_ (
    .a(_0540_),
    .b(_0542_),
    .y(_0543_)
  );
  al_nand2 _1259_ (
    .a(_0540_),
    .b(_0542_),
    .y(_0544_)
  );
  al_nand2ft _1260_ (
    .a(_0543_),
    .b(_0544_),
    .y(_0545_)
  );
  al_or2 _1261_ (
    .a(N18),
    .b(N58),
    .y(_0546_)
  );
  al_ao21ttf _1262_ (
    .a(N337),
    .b(N18),
    .c(_0546_),
    .y(_0547_)
  );
  al_inv _1263_ (
    .a(N340),
    .y(_0548_)
  );
  al_mux2h _1264_ (
    .a(N77),
    .b(_0548_),
    .s(N18),
    .y(_0549_)
  );
  al_and2ft _1265_ (
    .a(_0547_),
    .b(_0549_),
    .y(_0550_)
  );
  al_or2ft _1266_ (
    .a(_0547_),
    .b(_0549_),
    .y(_0551_)
  );
  al_or3ftt _1267_ (
    .a(_0551_),
    .b(_0550_),
    .c(_0545_),
    .y(_0552_)
  );
  al_aoi21ftf _1268_ (
    .a(_0550_),
    .b(_0551_),
    .c(_0545_),
    .y(_0553_)
  );
  al_nand2ft _1269_ (
    .a(_0553_),
    .b(_0552_),
    .y(_0554_)
  );
  al_or3fft _1270_ (
    .a(_0538_),
    .b(_0537_),
    .c(_0554_),
    .y(_0555_)
  );
  al_aoi21ttf _1271_ (
    .a(_0538_),
    .b(_0537_),
    .c(_0554_),
    .y(_0556_)
  );
  al_nand2ft _1272_ (
    .a(_0556_),
    .b(_0555_),
    .y(_0557_)
  );
  al_nand2ft _1273_ (
    .a(N18),
    .b(N114),
    .y(_0558_)
  );
  al_ao21ftf _1274_ (
    .a(N248),
    .b(N18),
    .c(_0558_),
    .y(_0559_)
  );
  al_inv _1275_ (
    .a(N251),
    .y(_0560_)
  );
  al_mux2h _1276_ (
    .a(N113),
    .b(_0560_),
    .s(N18),
    .y(_0561_)
  );
  al_nand2 _1277_ (
    .a(_0559_),
    .b(_0561_),
    .y(_0562_)
  );
  al_nor2 _1278_ (
    .a(_0559_),
    .b(_0561_),
    .y(_0563_)
  );
  al_nand2ft _1279_ (
    .a(_0563_),
    .b(_0562_),
    .y(_0564_)
  );
  al_inv _1280_ (
    .a(N257),
    .y(_0565_)
  );
  al_mux2h _1281_ (
    .a(N112),
    .b(_0565_),
    .s(N18),
    .y(_0566_)
  );
  al_inv _1282_ (
    .a(N260),
    .y(_0567_)
  );
  al_mux2h _1283_ (
    .a(N88),
    .b(_0567_),
    .s(N18),
    .y(_0568_)
  );
  al_and2ft _1284_ (
    .a(_0566_),
    .b(_0568_),
    .y(_0569_)
  );
  al_nand2ft _1285_ (
    .a(_0568_),
    .b(_0566_),
    .y(_0570_)
  );
  al_nand3ftt _1286_ (
    .a(_0569_),
    .b(_0570_),
    .c(_0564_),
    .y(_0571_)
  );
  al_aoi21ftt _1287_ (
    .a(_0569_),
    .b(_0570_),
    .c(_0564_),
    .y(_0572_)
  );
  al_inv _1288_ (
    .a(N254),
    .y(_0573_)
  );
  al_mux2h _1289_ (
    .a(N111),
    .b(_0573_),
    .s(N18),
    .y(_0574_)
  );
  al_inv _1290_ (
    .a(N106),
    .y(_0575_)
  );
  al_mux2h _1291_ (
    .a(N87),
    .b(_0575_),
    .s(N18),
    .y(_0576_)
  );
  al_nand2ft _1292_ (
    .a(_0574_),
    .b(_0576_),
    .y(_0577_)
  );
  al_nand2ft _1293_ (
    .a(_0576_),
    .b(_0574_),
    .y(_0578_)
  );
  al_nand2 _1294_ (
    .a(N263),
    .b(N267),
    .y(_0579_)
  );
  al_or2 _1295_ (
    .a(N263),
    .b(N267),
    .y(_0580_)
  );
  al_nand3 _1296_ (
    .a(N18),
    .b(_0580_),
    .c(_0579_),
    .y(_0581_)
  );
  al_nor2 _1297_ (
    .a(N245),
    .b(N271),
    .y(_0582_)
  );
  al_aoi21 _1298_ (
    .a(N245),
    .b(N271),
    .c(N18),
    .y(_0583_)
  );
  al_aoi21ftf _1299_ (
    .a(_0582_),
    .b(_0583_),
    .c(_0581_),
    .y(_0584_)
  );
  al_and3ftt _1300_ (
    .a(_0584_),
    .b(_0577_),
    .c(_0578_),
    .y(_0585_)
  );
  al_ao21ttf _1301_ (
    .a(_0577_),
    .b(_0578_),
    .c(_0584_),
    .y(_0586_)
  );
  al_and2ft _1302_ (
    .a(_0585_),
    .b(_0586_),
    .y(_0587_)
  );
  al_oai21ftf _1303_ (
    .a(_0571_),
    .b(_0572_),
    .c(_0587_),
    .y(_0588_)
  );
  al_and3ftt _1304_ (
    .a(_0572_),
    .b(_0571_),
    .c(_0587_),
    .y(_0589_)
  );
  al_aoi21 _1305_ (
    .a(_0511_),
    .b(_0510_),
    .c(_0488_),
    .y(_0590_)
  );
  al_ao21ftt _1306_ (
    .a(_0589_),
    .b(_0588_),
    .c(_0590_),
    .y(_0591_)
  );
  al_nand3ftt _1307_ (
    .a(_0591_),
    .b(_0557_),
    .c(_0514_),
    .y(N10575)
  );
  al_mux2l _1308_ (
    .a(N196),
    .b(N97),
    .s(N18),
    .y(_0592_)
  );
  al_mux2l _1309_ (
    .a(N195),
    .b(N94),
    .s(N18),
    .y(_0593_)
  );
  al_nand2 _1310_ (
    .a(_0592_),
    .b(_0593_),
    .y(_0594_)
  );
  al_nor2 _1311_ (
    .a(_0592_),
    .b(_0593_),
    .y(_0595_)
  );
  al_nand2ft _1312_ (
    .a(_0595_),
    .b(_0594_),
    .y(_0596_)
  );
  al_mux2l _1313_ (
    .a(N190),
    .b(N50),
    .s(N18),
    .y(_0597_)
  );
  al_mux2l _1314_ (
    .a(N189),
    .b(N66),
    .s(N18),
    .y(_0598_)
  );
  al_nor2 _1315_ (
    .a(_0597_),
    .b(_0598_),
    .y(_0599_)
  );
  al_nand2 _1316_ (
    .a(_0597_),
    .b(_0598_),
    .y(_0600_)
  );
  al_nand2ft _1317_ (
    .a(_0599_),
    .b(_0600_),
    .y(_0601_)
  );
  al_mux2l _1318_ (
    .a(N192),
    .b(N35),
    .s(N18),
    .y(_0602_)
  );
  al_mux2l _1319_ (
    .a(N191),
    .b(N32),
    .s(N18),
    .y(_0603_)
  );
  al_nand2 _1320_ (
    .a(_0602_),
    .b(_0603_),
    .y(_0604_)
  );
  al_nor2 _1321_ (
    .a(_0602_),
    .b(_0603_),
    .y(_0605_)
  );
  al_nand3ftt _1322_ (
    .a(_0605_),
    .b(_0604_),
    .c(_0601_),
    .y(_0606_)
  );
  al_ao21ftt _1323_ (
    .a(_0605_),
    .b(_0604_),
    .c(_0601_),
    .y(_0607_)
  );
  al_ao21 _1324_ (
    .a(_0606_),
    .b(_0607_),
    .c(_0596_),
    .y(_0608_)
  );
  al_and3 _1325_ (
    .a(_0596_),
    .b(_0606_),
    .c(_0607_),
    .y(_0609_)
  );
  al_mux2l _1326_ (
    .a(N194),
    .b(N121),
    .s(N18),
    .y(_0610_)
  );
  al_mux2l _1327_ (
    .a(N193),
    .b(N47),
    .s(N18),
    .y(_0611_)
  );
  al_nand2 _1328_ (
    .a(_0610_),
    .b(_0611_),
    .y(_0612_)
  );
  al_nor2 _1329_ (
    .a(_0610_),
    .b(_0611_),
    .y(_0613_)
  );
  al_nand2ft _1330_ (
    .a(_0613_),
    .b(_0612_),
    .y(_0614_)
  );
  al_mux2l _1331_ (
    .a(N197),
    .b(N115),
    .s(N18),
    .y(_0615_)
  );
  al_mux2l _1332_ (
    .a(N187),
    .b(N118),
    .s(N18),
    .y(_0616_)
  );
  al_nor2 _1333_ (
    .a(_0615_),
    .b(_0616_),
    .y(_0617_)
  );
  al_nand2 _1334_ (
    .a(_0615_),
    .b(_0616_),
    .y(_0618_)
  );
  al_or3ftt _1335_ (
    .a(_0618_),
    .b(_0617_),
    .c(_0614_),
    .y(_0619_)
  );
  al_aoi21ftf _1336_ (
    .a(_0617_),
    .b(_0618_),
    .c(_0614_),
    .y(_0620_)
  );
  al_nand2ft _1337_ (
    .a(_0620_),
    .b(_0619_),
    .y(_0621_)
  );
  al_ao21ftf _1338_ (
    .a(_0609_),
    .b(_0608_),
    .c(_0621_),
    .y(_0622_)
  );
  al_and3fft _1339_ (
    .a(_0609_),
    .b(_0621_),
    .c(_0608_),
    .y(_0623_)
  );
  al_mux2l _1340_ (
    .a(N208),
    .b(N44),
    .s(N18),
    .y(_0624_)
  );
  al_mux2l _1341_ (
    .a(N198),
    .b(N41),
    .s(N18),
    .y(_0625_)
  );
  al_and2ft _1342_ (
    .a(_0624_),
    .b(_0625_),
    .y(_0626_)
  );
  al_nand2ft _1343_ (
    .a(_0625_),
    .b(_0624_),
    .y(_0627_)
  );
  al_nand2ft _1344_ (
    .a(_0626_),
    .b(_0627_),
    .y(_0628_)
  );
  al_mux2l _1345_ (
    .a(N207),
    .b(N29),
    .s(N18),
    .y(_0629_)
  );
  al_mux2l _1346_ (
    .a(N206),
    .b(N26),
    .s(N18),
    .y(_0630_)
  );
  al_nand2 _1347_ (
    .a(_0629_),
    .b(_0630_),
    .y(_0631_)
  );
  al_nor2 _1348_ (
    .a(_0629_),
    .b(_0630_),
    .y(_0632_)
  );
  al_mux2l _1349_ (
    .a(N205),
    .b(N23),
    .s(N18),
    .y(_0633_)
  );
  al_mux2l _1350_ (
    .a(N204),
    .b(N103),
    .s(N18),
    .y(_0634_)
  );
  al_and2ft _1351_ (
    .a(_0633_),
    .b(_0634_),
    .y(_0635_)
  );
  al_nand2ft _1352_ (
    .a(_0634_),
    .b(_0633_),
    .y(_0636_)
  );
  al_and2ft _1353_ (
    .a(_0635_),
    .b(_0636_),
    .y(_0637_)
  );
  al_nand3ftt _1354_ (
    .a(_0632_),
    .b(_0631_),
    .c(_0637_),
    .y(_0638_)
  );
  al_ao21ftt _1355_ (
    .a(_0632_),
    .b(_0631_),
    .c(_0637_),
    .y(_0639_)
  );
  al_ao21 _1356_ (
    .a(_0638_),
    .b(_0639_),
    .c(_0628_),
    .y(_0640_)
  );
  al_nand3 _1357_ (
    .a(_0628_),
    .b(_0638_),
    .c(_0639_),
    .y(_0641_)
  );
  al_mux2l _1358_ (
    .a(N201),
    .b(N124),
    .s(N18),
    .y(_0642_)
  );
  al_mux2l _1359_ (
    .a(N200),
    .b(N100),
    .s(N18),
    .y(_0643_)
  );
  al_nor2 _1360_ (
    .a(_0642_),
    .b(_0643_),
    .y(_0644_)
  );
  al_nand2 _1361_ (
    .a(_0642_),
    .b(_0643_),
    .y(_0645_)
  );
  al_mux2l _1362_ (
    .a(N203),
    .b(N130),
    .s(N18),
    .y(_0646_)
  );
  al_mux2l _1363_ (
    .a(N202),
    .b(N127),
    .s(N18),
    .y(_0647_)
  );
  al_nand2 _1364_ (
    .a(_0646_),
    .b(_0647_),
    .y(_0648_)
  );
  al_nor2 _1365_ (
    .a(_0646_),
    .b(_0647_),
    .y(_0649_)
  );
  al_nand2ft _1366_ (
    .a(_0649_),
    .b(_0648_),
    .y(_0650_)
  );
  al_aoi21ftt _1367_ (
    .a(_0644_),
    .b(_0645_),
    .c(_0650_),
    .y(_0651_)
  );
  al_and3ftt _1368_ (
    .a(_0644_),
    .b(_0645_),
    .c(_0650_),
    .y(_0652_)
  );
  al_or2 _1369_ (
    .a(_0652_),
    .b(_0651_),
    .y(_0653_)
  );
  al_ao21ttf _1370_ (
    .a(_0641_),
    .b(_0640_),
    .c(_0653_),
    .y(_0654_)
  );
  al_nand3ftt _1371_ (
    .a(_0623_),
    .b(_0622_),
    .c(_0654_),
    .y(_0655_)
  );
  al_aoi21ftf _1372_ (
    .a(N174),
    .b(N18),
    .c(_0346_),
    .y(_0656_)
  );
  al_nand2ft _1373_ (
    .a(N173),
    .b(N18),
    .y(_0657_)
  );
  al_nand2ft _1374_ (
    .a(N174),
    .b(N18),
    .y(_0658_)
  );
  al_nand3ftt _1375_ (
    .a(_0658_),
    .b(_0346_),
    .c(_0657_),
    .y(_0659_)
  );
  al_aoi21ftf _1376_ (
    .a(_0657_),
    .b(_0656_),
    .c(_0659_),
    .y(_0660_)
  );
  al_mux2l _1377_ (
    .a(N181),
    .b(N141),
    .s(N18),
    .y(_0661_)
  );
  al_mux2l _1378_ (
    .a(N171),
    .b(N147),
    .s(N18),
    .y(_0662_)
  );
  al_and2ft _1379_ (
    .a(_0661_),
    .b(_0662_),
    .y(_0663_)
  );
  al_nand2ft _1380_ (
    .a(_0662_),
    .b(_0661_),
    .y(_0664_)
  );
  al_aoi21ftf _1381_ (
    .a(N176),
    .b(N18),
    .c(_0346_),
    .y(_0665_)
  );
  al_nand2ft _1382_ (
    .a(N175),
    .b(N18),
    .y(_0666_)
  );
  al_nand2ft _1383_ (
    .a(N176),
    .b(N18),
    .y(_0667_)
  );
  al_nand3ftt _1384_ (
    .a(_0667_),
    .b(_0346_),
    .c(_0666_),
    .y(_0668_)
  );
  al_aoi21ftf _1385_ (
    .a(_0666_),
    .b(_0665_),
    .c(_0668_),
    .y(_0669_)
  );
  al_nand3ftt _1386_ (
    .a(_0663_),
    .b(_0664_),
    .c(_0669_),
    .y(_0670_)
  );
  al_ao21ftt _1387_ (
    .a(_0663_),
    .b(_0664_),
    .c(_0669_),
    .y(_0671_)
  );
  al_ao21 _1388_ (
    .a(_0670_),
    .b(_0671_),
    .c(_0660_),
    .y(_0672_)
  );
  al_and3 _1389_ (
    .a(_0660_),
    .b(_0670_),
    .c(_0671_),
    .y(_0673_)
  );
  al_mux2l _1390_ (
    .a(N178),
    .b(N135),
    .s(N18),
    .y(_0674_)
  );
  al_ao21ftf _1391_ (
    .a(N177),
    .b(N18),
    .c(_0346_),
    .y(_0675_)
  );
  al_and2 _1392_ (
    .a(_0674_),
    .b(_0675_),
    .y(_0676_)
  );
  al_or2 _1393_ (
    .a(_0674_),
    .b(_0675_),
    .y(_0677_)
  );
  al_mux2l _1394_ (
    .a(N180),
    .b(N138),
    .s(N18),
    .y(_0678_)
  );
  al_mux2l _1395_ (
    .a(N179),
    .b(N144),
    .s(N18),
    .y(_0679_)
  );
  al_and2ft _1396_ (
    .a(_0679_),
    .b(_0678_),
    .y(_0680_)
  );
  al_nand2ft _1397_ (
    .a(_0678_),
    .b(_0679_),
    .y(_0681_)
  );
  al_nand2ft _1398_ (
    .a(_0680_),
    .b(_0681_),
    .y(_0682_)
  );
  al_and3ftt _1399_ (
    .a(_0676_),
    .b(_0677_),
    .c(_0682_),
    .y(_0683_)
  );
  al_ao21ftt _1400_ (
    .a(_0676_),
    .b(_0677_),
    .c(_0682_),
    .y(_0684_)
  );
  al_nand2ft _1401_ (
    .a(_0683_),
    .b(_0684_),
    .y(_0685_)
  );
  al_and3fft _1402_ (
    .a(_0673_),
    .b(_0685_),
    .c(_0672_),
    .y(_0686_)
  );
  al_aoi21ftf _1403_ (
    .a(_0673_),
    .b(_0672_),
    .c(_0685_),
    .y(_0687_)
  );
  al_or2 _1404_ (
    .a(_0687_),
    .b(_0686_),
    .y(_0688_)
  );
  al_nand2ft _1405_ (
    .a(N167),
    .b(N18),
    .y(_0689_)
  );
  al_ao21ttf _1406_ (
    .a(N12),
    .b(N9),
    .c(_0689_),
    .y(_0690_)
  );
  al_nand2ft _1407_ (
    .a(N166),
    .b(N18),
    .y(_0691_)
  );
  al_nand3ftt _1408_ (
    .a(_0689_),
    .b(_0346_),
    .c(_0691_),
    .y(_0692_)
  );
  al_oa21 _1409_ (
    .a(_0691_),
    .b(_0690_),
    .c(_0692_),
    .y(_0693_)
  );
  al_oa21 _1410_ (
    .a(N170),
    .b(_0391_),
    .c(_0693_),
    .y(_0694_)
  );
  al_or3 _1411_ (
    .a(N170),
    .b(_0391_),
    .c(_0693_),
    .y(_0695_)
  );
  al_nand2ft _1412_ (
    .a(_0694_),
    .b(_0695_),
    .y(_0696_)
  );
  al_nand2ft _1413_ (
    .a(N169),
    .b(N18),
    .y(_0697_)
  );
  al_aoi21ttf _1414_ (
    .a(N12),
    .b(N9),
    .c(_0697_),
    .y(_0698_)
  );
  al_nand2ft _1415_ (
    .a(N168),
    .b(N18),
    .y(_0699_)
  );
  al_nand3ftt _1416_ (
    .a(_0697_),
    .b(_0346_),
    .c(_0699_),
    .y(_0700_)
  );
  al_aoi21ftf _1417_ (
    .a(_0699_),
    .b(_0698_),
    .c(_0700_),
    .y(_0701_)
  );
  al_nor2 _1418_ (
    .a(N165),
    .b(N164),
    .y(_0702_)
  );
  al_nand2 _1419_ (
    .a(N165),
    .b(N164),
    .y(_0703_)
  );
  al_nand3fft _1420_ (
    .a(_0391_),
    .b(_0702_),
    .c(_0703_),
    .y(_0704_)
  );
  al_nand2ft _1421_ (
    .a(_0704_),
    .b(_0701_),
    .y(_0705_)
  );
  al_or2ft _1422_ (
    .a(_0704_),
    .b(_0701_),
    .y(_0706_)
  );
  al_and3 _1423_ (
    .a(_0705_),
    .b(_0706_),
    .c(_0696_),
    .y(_0707_)
  );
  al_aoi21 _1424_ (
    .a(_0705_),
    .b(_0706_),
    .c(_0696_),
    .y(_0708_)
  );
  al_or3fft _1425_ (
    .a(_0641_),
    .b(_0640_),
    .c(_0653_),
    .y(_0709_)
  );
  al_oai21 _1426_ (
    .a(_0707_),
    .b(_0708_),
    .c(_0709_),
    .y(_0710_)
  );
  al_or3 _1427_ (
    .a(_0710_),
    .b(_0688_),
    .c(_0655_),
    .y(N10576)
  );
  al_and2ft _1428_ (
    .a(N277),
    .b(_0357_),
    .y(_0711_)
  );
  al_or2ft _1429_ (
    .a(N277),
    .b(_0357_),
    .y(_0712_)
  );
  al_nand2ft _1430_ (
    .a(_0711_),
    .b(_0712_),
    .y(_0713_)
  );
  al_nand2ft _1431_ (
    .a(N364),
    .b(_0418_),
    .y(_0714_)
  );
  al_or2ft _1432_ (
    .a(N364),
    .b(_0418_),
    .y(_0715_)
  );
  al_inv _1433_ (
    .a(_0715_),
    .y(_0716_)
  );
  al_or2ft _1434_ (
    .a(N361),
    .b(_0417_),
    .y(_0717_)
  );
  al_and2ft _1435_ (
    .a(N361),
    .b(_0417_),
    .y(_0718_)
  );
  al_or2ft _1436_ (
    .a(N358),
    .b(_0422_),
    .y(_0719_)
  );
  al_and2ft _1437_ (
    .a(N358),
    .b(_0422_),
    .y(_0720_)
  );
  al_nand2ft _1438_ (
    .a(N355),
    .b(_0421_),
    .y(_0721_)
  );
  al_oai21ftt _1439_ (
    .a(_0721_),
    .b(_0720_),
    .c(_0719_),
    .y(_0722_)
  );
  al_oa21ftf _1440_ (
    .a(_0717_),
    .b(_0722_),
    .c(_0718_),
    .y(_0723_)
  );
  al_and2ft _1441_ (
    .a(_0720_),
    .b(_0719_),
    .y(_0724_)
  );
  al_nor2ft _1442_ (
    .a(N355),
    .b(_0421_),
    .y(_0725_)
  );
  al_and3ftt _1443_ (
    .a(_0725_),
    .b(_0721_),
    .c(_0724_),
    .y(_0726_)
  );
  al_aoi21ttf _1444_ (
    .a(_0717_),
    .b(_0726_),
    .c(_0723_),
    .y(_0727_)
  );
  al_or2ft _1445_ (
    .a(N349),
    .b(_0400_),
    .y(_0728_)
  );
  al_and2ft _1446_ (
    .a(N349),
    .b(_0400_),
    .y(_0729_)
  );
  al_nand2ft _1447_ (
    .a(_0729_),
    .b(_0728_),
    .y(_0730_)
  );
  al_nand2ft _1448_ (
    .a(N340),
    .b(_0413_),
    .y(_0731_)
  );
  al_aoi21ftf _1449_ (
    .a(_0405_),
    .b(N343),
    .c(_0731_),
    .y(_0732_)
  );
  al_nand2ft _1450_ (
    .a(N343),
    .b(_0405_),
    .y(_0733_)
  );
  al_ao21ftf _1451_ (
    .a(_0413_),
    .b(N340),
    .c(_0733_),
    .y(_0734_)
  );
  al_nor2ft _1452_ (
    .a(N346),
    .b(_0406_),
    .y(_0735_)
  );
  al_and2ft _1453_ (
    .a(N346),
    .b(_0406_),
    .y(_0736_)
  );
  al_nor2 _1454_ (
    .a(_0736_),
    .b(_0735_),
    .y(_0737_)
  );
  al_nand3ftt _1455_ (
    .a(_0734_),
    .b(_0732_),
    .c(_0737_),
    .y(_0738_)
  );
  al_nand2ft _1456_ (
    .a(N352),
    .b(_0401_),
    .y(_0739_)
  );
  al_or2ft _1457_ (
    .a(N352),
    .b(_0401_),
    .y(_0740_)
  );
  al_and2 _1458_ (
    .a(_0739_),
    .b(_0740_),
    .y(_0741_)
  );
  al_or3ftt _1459_ (
    .a(_0741_),
    .b(_0730_),
    .c(_0738_),
    .y(_0742_)
  );
  al_or2ft _1460_ (
    .a(N334),
    .b(_0320_),
    .y(_0743_)
  );
  al_and2ft _1461_ (
    .a(N334),
    .b(_0320_),
    .y(_0744_)
  );
  al_nor2ft _1462_ (
    .a(N331),
    .b(_0316_),
    .y(_0745_)
  );
  al_and2ft _1463_ (
    .a(N331),
    .b(_0316_),
    .y(_0746_)
  );
  al_or2ft _1464_ (
    .a(N328),
    .b(_0331_),
    .y(_0747_)
  );
  al_and2ft _1465_ (
    .a(N328),
    .b(_0331_),
    .y(_0748_)
  );
  al_and2ft _1466_ (
    .a(N325),
    .b(_0330_),
    .y(_0749_)
  );
  al_oa21 _1467_ (
    .a(_0748_),
    .b(_0749_),
    .c(_0747_),
    .y(_0750_)
  );
  al_oai21ttf _1468_ (
    .a(_0746_),
    .b(_0750_),
    .c(_0745_),
    .y(_0751_)
  );
  al_ao21ftf _1469_ (
    .a(_0744_),
    .b(_0751_),
    .c(_0743_),
    .y(_0752_)
  );
  al_nand3fft _1470_ (
    .a(_0285_),
    .b(_0289_),
    .c(_0299_),
    .y(_0753_)
  );
  al_ao21ttf _1471_ (
    .a(_0287_),
    .b(_0753_),
    .c(_0283_),
    .y(_0754_)
  );
  al_nand3fft _1472_ (
    .a(N367),
    .b(_0282_),
    .c(_0754_),
    .y(_0755_)
  );
  al_nand2ft _1473_ (
    .a(_0290_),
    .b(_0296_),
    .y(_0756_)
  );
  al_nand3fft _1474_ (
    .a(_0294_),
    .b(_0756_),
    .c(_0307_),
    .y(_0757_)
  );
  al_nand3 _1475_ (
    .a(_0287_),
    .b(_0753_),
    .c(_0757_),
    .y(_0758_)
  );
  al_ao21 _1476_ (
    .a(_0283_),
    .b(_0758_),
    .c(_0282_),
    .y(_0759_)
  );
  al_and2ft _1477_ (
    .a(_0748_),
    .b(_0747_),
    .y(_0760_)
  );
  al_or2ft _1478_ (
    .a(N325),
    .b(_0330_),
    .y(_0761_)
  );
  al_and3ftt _1479_ (
    .a(_0749_),
    .b(_0761_),
    .c(_0760_),
    .y(_0762_)
  );
  al_nor2 _1480_ (
    .a(_0746_),
    .b(_0745_),
    .y(_0763_)
  );
  al_and2ft _1481_ (
    .a(_0744_),
    .b(_0743_),
    .y(_0764_)
  );
  al_and3 _1482_ (
    .a(_0763_),
    .b(_0764_),
    .c(_0762_),
    .y(_0765_)
  );
  al_nand3 _1483_ (
    .a(_0765_),
    .b(_0755_),
    .c(_0759_),
    .y(_0766_)
  );
  al_ao21 _1484_ (
    .a(_0752_),
    .b(_0766_),
    .c(_0742_),
    .y(_0767_)
  );
  al_or2ft _1485_ (
    .a(N343),
    .b(_0405_),
    .y(_0768_)
  );
  al_ao21ttf _1486_ (
    .a(_0731_),
    .b(_0733_),
    .c(_0768_),
    .y(_0769_)
  );
  al_oa21ttf _1487_ (
    .a(_0735_),
    .b(_0769_),
    .c(_0736_),
    .y(_0770_)
  );
  al_oa21ftf _1488_ (
    .a(_0728_),
    .b(_0770_),
    .c(_0729_),
    .y(_0771_)
  );
  al_oa21ftt _1489_ (
    .a(_0740_),
    .b(_0771_),
    .c(_0739_),
    .y(_0772_)
  );
  al_nand3 _1490_ (
    .a(_0723_),
    .b(_0772_),
    .c(_0767_),
    .y(_0773_)
  );
  al_nand3fft _1491_ (
    .a(_0716_),
    .b(_0727_),
    .c(_0773_),
    .y(_0774_)
  );
  al_ao21 _1492_ (
    .a(_0714_),
    .b(_0774_),
    .c(_0713_),
    .y(_0775_)
  );
  al_and3 _1493_ (
    .a(_0713_),
    .b(_0714_),
    .c(_0774_),
    .y(_0776_)
  );
  al_and2ft _1494_ (
    .a(_0776_),
    .b(_0775_),
    .y(N10632)
  );
  al_nand3ftt _1495_ (
    .a(N251),
    .b(_0377_),
    .c(_0346_),
    .y(_0777_)
  );
  al_ao21 _1496_ (
    .a(_0377_),
    .b(_0346_),
    .c(_0560_),
    .y(_0778_)
  );
  al_and2 _1497_ (
    .a(_0777_),
    .b(_0778_),
    .y(_0779_)
  );
  al_inv _1498_ (
    .a(_0779_),
    .y(_0780_)
  );
  al_aoi21 _1499_ (
    .a(_0351_),
    .b(_0346_),
    .c(_0480_),
    .y(_0781_)
  );
  al_and3ftt _1500_ (
    .a(N299),
    .b(_0351_),
    .c(_0346_),
    .y(_0782_)
  );
  al_nor2 _1501_ (
    .a(_0782_),
    .b(_0781_),
    .y(_0783_)
  );
  al_nand3ftt _1502_ (
    .a(N293),
    .b(_0345_),
    .c(_0346_),
    .y(_0784_)
  );
  al_ao21 _1503_ (
    .a(_0347_),
    .b(_0346_),
    .c(_0502_),
    .y(_0785_)
  );
  al_ao21 _1504_ (
    .a(_0345_),
    .b(_0346_),
    .c(_0500_),
    .y(_0786_)
  );
  al_nand3ftt _1505_ (
    .a(N296),
    .b(_0347_),
    .c(_0346_),
    .y(_0787_)
  );
  al_and3 _1506_ (
    .a(_0787_),
    .b(_0785_),
    .c(_0786_),
    .y(_0788_)
  );
  al_nand2 _1507_ (
    .a(_0784_),
    .b(_0788_),
    .y(_0789_)
  );
  al_inv _1508_ (
    .a(_0789_),
    .y(_0790_)
  );
  al_nor2ft _1509_ (
    .a(N289),
    .b(_0365_),
    .y(_0791_)
  );
  al_and2ft _1510_ (
    .a(N289),
    .b(_0365_),
    .y(_0792_)
  );
  al_or2ft _1511_ (
    .a(N286),
    .b(_0364_),
    .y(_0793_)
  );
  al_and2ft _1512_ (
    .a(N286),
    .b(_0364_),
    .y(_0794_)
  );
  al_and2ft _1513_ (
    .a(N283),
    .b(_0369_),
    .y(_0795_)
  );
  al_or2ft _1514_ (
    .a(N283),
    .b(_0369_),
    .y(_0796_)
  );
  al_and2ft _1515_ (
    .a(N280),
    .b(_0368_),
    .y(_0797_)
  );
  al_nor2ft _1516_ (
    .a(N280),
    .b(_0368_),
    .y(_0798_)
  );
  al_oai21ftf _1517_ (
    .a(_0711_),
    .b(_0798_),
    .c(_0797_),
    .y(_0799_)
  );
  al_ao21 _1518_ (
    .a(_0796_),
    .b(_0799_),
    .c(_0795_),
    .y(_0800_)
  );
  al_oai21 _1519_ (
    .a(_0794_),
    .b(_0800_),
    .c(_0793_),
    .y(_0801_)
  );
  al_and2ft _1520_ (
    .a(_0792_),
    .b(_0801_),
    .y(_0802_)
  );
  al_nor2 _1521_ (
    .a(_0797_),
    .b(_0798_),
    .y(_0803_)
  );
  al_and2ft _1522_ (
    .a(_0794_),
    .b(_0793_),
    .y(_0804_)
  );
  al_and3ftt _1523_ (
    .a(_0795_),
    .b(_0796_),
    .c(_0804_),
    .y(_0805_)
  );
  al_nand3ftt _1524_ (
    .a(_0713_),
    .b(_0803_),
    .c(_0805_),
    .y(_0806_)
  );
  al_aoi21 _1525_ (
    .a(_0806_),
    .b(_0802_),
    .c(_0791_),
    .y(_0807_)
  );
  al_nand3 _1526_ (
    .a(_0714_),
    .b(_0802_),
    .c(_0774_),
    .y(_0808_)
  );
  al_and3 _1527_ (
    .a(_0790_),
    .b(_0807_),
    .c(_0808_),
    .y(_0809_)
  );
  al_ao21 _1528_ (
    .a(_0353_),
    .b(_0346_),
    .c(_0482_),
    .y(_0810_)
  );
  al_and3ftt _1529_ (
    .a(N303),
    .b(_0353_),
    .c(_0346_),
    .y(_0811_)
  );
  al_and2ft _1530_ (
    .a(_0811_),
    .b(_0810_),
    .y(_0812_)
  );
  al_nand3 _1531_ (
    .a(_0783_),
    .b(_0812_),
    .c(_0809_),
    .y(_0813_)
  );
  al_ao21ttf _1532_ (
    .a(_0787_),
    .b(_0784_),
    .c(_0785_),
    .y(_0814_)
  );
  al_aoi21ftt _1533_ (
    .a(_0782_),
    .b(_0814_),
    .c(_0781_),
    .y(_0815_)
  );
  al_aoi21 _1534_ (
    .a(_0810_),
    .b(_0815_),
    .c(_0811_),
    .y(_0816_)
  );
  al_ao21 _1535_ (
    .a(_0816_),
    .b(_0813_),
    .c(_0780_),
    .y(_0817_)
  );
  al_and3 _1536_ (
    .a(_0780_),
    .b(_0816_),
    .c(_0813_),
    .y(_0818_)
  );
  al_and2ft _1537_ (
    .a(_0818_),
    .b(_0817_),
    .y(N10641)
  );
  al_or2 _1538_ (
    .a(_0792_),
    .b(_0791_),
    .y(_0819_)
  );
  al_nand3ftt _1539_ (
    .a(_0711_),
    .b(_0712_),
    .c(_0803_),
    .y(_0820_)
  );
  al_ao21 _1540_ (
    .a(_0714_),
    .b(_0774_),
    .c(_0820_),
    .y(_0821_)
  );
  al_oai21ftt _1541_ (
    .a(_0805_),
    .b(_0821_),
    .c(_0801_),
    .y(_0822_)
  );
  al_or2 _1542_ (
    .a(_0819_),
    .b(_0822_),
    .y(_0823_)
  );
  al_and2 _1543_ (
    .a(_0819_),
    .b(_0822_),
    .y(_0824_)
  );
  al_nand2ft _1544_ (
    .a(_0824_),
    .b(_0823_),
    .y(N10711)
  );
  al_nand2 _1545_ (
    .a(_0714_),
    .b(_0774_),
    .y(_0825_)
  );
  al_and2ft _1546_ (
    .a(_0795_),
    .b(_0796_),
    .y(_0826_)
  );
  al_nand3ftt _1547_ (
    .a(_0820_),
    .b(_0826_),
    .c(_0825_),
    .y(_0827_)
  );
  al_and3ftt _1548_ (
    .a(_0800_),
    .b(_0804_),
    .c(_0827_),
    .y(_0828_)
  );
  al_ao21ftt _1549_ (
    .a(_0800_),
    .b(_0827_),
    .c(_0804_),
    .y(_0829_)
  );
  al_nand2ft _1550_ (
    .a(_0828_),
    .b(_0829_),
    .y(N10712)
  );
  al_inv _1551_ (
    .a(_0799_),
    .y(_0830_)
  );
  al_ao21 _1552_ (
    .a(_0830_),
    .b(_0821_),
    .c(_0826_),
    .y(_0831_)
  );
  al_and3 _1553_ (
    .a(_0830_),
    .b(_0826_),
    .c(_0821_),
    .y(_0832_)
  );
  al_nand2ft _1554_ (
    .a(_0832_),
    .b(_0831_),
    .y(N10713)
  );
  al_and3ftt _1555_ (
    .a(_0711_),
    .b(_0803_),
    .c(_0775_),
    .y(_0833_)
  );
  al_ao21ftt _1556_ (
    .a(_0711_),
    .b(_0775_),
    .c(_0803_),
    .y(_0834_)
  );
  al_nand2ft _1557_ (
    .a(_0833_),
    .b(_0834_),
    .y(N10714)
  );
  al_and3ftt _1558_ (
    .a(N257),
    .b(_0378_),
    .c(_0346_),
    .y(_0835_)
  );
  al_ao21 _1559_ (
    .a(_0378_),
    .b(_0346_),
    .c(_0565_),
    .y(_0836_)
  );
  al_and3ftt _1560_ (
    .a(N106),
    .b(_0388_),
    .c(_0346_),
    .y(_0837_)
  );
  al_ao21 _1561_ (
    .a(_0388_),
    .b(_0346_),
    .c(_0575_),
    .y(_0838_)
  );
  al_and3ftt _1562_ (
    .a(N254),
    .b(_0386_),
    .c(_0346_),
    .y(_0839_)
  );
  al_aoi21 _1563_ (
    .a(_0386_),
    .b(_0346_),
    .c(_0573_),
    .y(_0840_)
  );
  al_oai21ttf _1564_ (
    .a(_0777_),
    .b(_0840_),
    .c(_0839_),
    .y(_0841_)
  );
  al_ao21 _1565_ (
    .a(_0838_),
    .b(_0841_),
    .c(_0837_),
    .y(_0842_)
  );
  al_aoi21 _1566_ (
    .a(_0836_),
    .b(_0842_),
    .c(_0835_),
    .y(_0843_)
  );
  al_and2ft _1567_ (
    .a(_0837_),
    .b(_0838_),
    .y(_0844_)
  );
  al_nor2 _1568_ (
    .a(_0839_),
    .b(_0840_),
    .y(_0845_)
  );
  al_nand3 _1569_ (
    .a(_0844_),
    .b(_0779_),
    .c(_0845_),
    .y(_0846_)
  );
  al_ao21 _1570_ (
    .a(_0816_),
    .b(_0813_),
    .c(_0846_),
    .y(_0847_)
  );
  al_or3ftt _1571_ (
    .a(_0836_),
    .b(_0835_),
    .c(_0847_),
    .y(_0848_)
  );
  al_and3ftt _1572_ (
    .a(N260),
    .b(_0380_),
    .c(_0346_),
    .y(_0849_)
  );
  al_aoi21 _1573_ (
    .a(_0380_),
    .b(_0346_),
    .c(_0567_),
    .y(_0850_)
  );
  al_nor2 _1574_ (
    .a(_0849_),
    .b(_0850_),
    .y(_0851_)
  );
  al_and3 _1575_ (
    .a(_0843_),
    .b(_0851_),
    .c(_0848_),
    .y(_0852_)
  );
  al_ao21 _1576_ (
    .a(_0843_),
    .b(_0848_),
    .c(_0851_),
    .y(_0853_)
  );
  al_nand2ft _1577_ (
    .a(_0852_),
    .b(_0853_),
    .y(N10715)
  );
  al_and2ft _1578_ (
    .a(_0835_),
    .b(_0836_),
    .y(_0854_)
  );
  al_ao21ftt _1579_ (
    .a(_0842_),
    .b(_0847_),
    .c(_0854_),
    .y(_0855_)
  );
  al_and3ftt _1580_ (
    .a(_0842_),
    .b(_0854_),
    .c(_0847_),
    .y(_0856_)
  );
  al_nand2ft _1581_ (
    .a(_0856_),
    .b(_0855_),
    .y(N10716)
  );
  al_oa21ftf _1582_ (
    .a(_0845_),
    .b(_0817_),
    .c(_0841_),
    .y(_0857_)
  );
  al_or2 _1583_ (
    .a(_0844_),
    .b(_0857_),
    .y(_0858_)
  );
  al_and2 _1584_ (
    .a(_0844_),
    .b(_0857_),
    .y(_0859_)
  );
  al_nand2ft _1585_ (
    .a(_0859_),
    .b(_0858_),
    .y(N10717)
  );
  al_and3 _1586_ (
    .a(_0777_),
    .b(_0845_),
    .c(_0817_),
    .y(_0860_)
  );
  al_ao21 _1587_ (
    .a(_0777_),
    .b(_0817_),
    .c(_0845_),
    .y(_0861_)
  );
  al_nand2ft _1588_ (
    .a(_0860_),
    .b(_0861_),
    .y(N10718)
  );
  al_and2ft _1589_ (
    .a(N883),
    .b(_0271_),
    .y(_0862_)
  );
  al_and3 _1590_ (
    .a(_0274_),
    .b(_0276_),
    .c(_0862_),
    .y(_0863_)
  );
  al_nand3 _1591_ (
    .a(_0344_),
    .b(_0863_),
    .c(_0433_),
    .y(_0864_)
  );
  al_or3 _1592_ (
    .a(N10576),
    .b(_0864_),
    .c(N10575),
    .y(N10729)
  );
  al_or2ft _1593_ (
    .a(N340),
    .b(_0413_),
    .y(_0865_)
  );
  al_nand2 _1594_ (
    .a(_0752_),
    .b(_0766_),
    .y(_0866_)
  );
  al_nand3 _1595_ (
    .a(_0731_),
    .b(_0865_),
    .c(_0866_),
    .y(_0867_)
  );
  al_aoi21 _1596_ (
    .a(_0731_),
    .b(_0865_),
    .c(_0866_),
    .y(_0868_)
  );
  al_nor2ft _1597_ (
    .a(_0867_),
    .b(_0868_),
    .y(N10827)
  );
  al_nand3 _1598_ (
    .a(_0733_),
    .b(_0768_),
    .c(_0865_),
    .y(_0869_)
  );
  al_and3ftt _1599_ (
    .a(_0729_),
    .b(_0728_),
    .c(_0737_),
    .y(_0870_)
  );
  al_nand3ftt _1600_ (
    .a(_0869_),
    .b(_0731_),
    .c(_0870_),
    .y(_0871_)
  );
  al_ao21 _1601_ (
    .a(_0752_),
    .b(_0766_),
    .c(_0871_),
    .y(_0872_)
  );
  al_nor2ft _1602_ (
    .a(_0740_),
    .b(_0771_),
    .y(_0873_)
  );
  al_and2ft _1603_ (
    .a(_0741_),
    .b(_0771_),
    .y(_0874_)
  );
  al_ao21 _1604_ (
    .a(_0739_),
    .b(_0873_),
    .c(_0874_),
    .y(_0875_)
  );
  al_aoi21ttf _1605_ (
    .a(_0875_),
    .b(_0872_),
    .c(_0767_),
    .y(N10868)
  );
  al_aoi21ftf _1606_ (
    .a(_0738_),
    .b(_0866_),
    .c(_0770_),
    .y(_0876_)
  );
  al_and2ft _1607_ (
    .a(_0730_),
    .b(_0876_),
    .y(_0877_)
  );
  al_or2ft _1608_ (
    .a(_0730_),
    .b(_0876_),
    .y(_0878_)
  );
  al_nand2ft _1609_ (
    .a(_0877_),
    .b(_0878_),
    .y(N10869)
  );
  al_and2 _1610_ (
    .a(_0733_),
    .b(_0768_),
    .y(_0879_)
  );
  al_oai21ftt _1611_ (
    .a(_0879_),
    .b(_0867_),
    .c(_0769_),
    .y(_0880_)
  );
  al_and2ft _1612_ (
    .a(_0737_),
    .b(_0880_),
    .y(_0881_)
  );
  al_or3 _1613_ (
    .a(_0735_),
    .b(_0736_),
    .c(_0880_),
    .y(_0882_)
  );
  al_nand2ft _1614_ (
    .a(_0881_),
    .b(_0882_),
    .y(N10870)
  );
  al_and3 _1615_ (
    .a(_0731_),
    .b(_0879_),
    .c(_0867_),
    .y(_0883_)
  );
  al_ao21 _1616_ (
    .a(_0731_),
    .b(_0867_),
    .c(_0879_),
    .y(_0884_)
  );
  al_nand2ft _1617_ (
    .a(_0883_),
    .b(_0884_),
    .y(N10871)
  );
  al_and2 _1618_ (
    .a(N163),
    .b(N1),
    .y(N1781)
  );
  al_nand3ftt _1619_ (
    .a(N38),
    .b(N267),
    .c(N382),
    .y(_0885_)
  );
  al_aoi21ttf _1620_ (
    .a(N267),
    .b(N382),
    .c(N38),
    .y(_0886_)
  );
  al_aoi21ftt _1621_ (
    .a(N263),
    .b(N38),
    .c(_0886_),
    .y(_0887_)
  );
  al_nand3 _1622_ (
    .a(N263),
    .b(N38),
    .c(N382),
    .y(_0888_)
  );
  al_aoi21 _1623_ (
    .a(N263),
    .b(N382),
    .c(N38),
    .y(_0889_)
  );
  al_and3ftt _1624_ (
    .a(_0835_),
    .b(_0836_),
    .c(_0851_),
    .y(_0890_)
  );
  al_oai21ftf _1625_ (
    .a(_0835_),
    .b(_0850_),
    .c(_0849_),
    .y(_0891_)
  );
  al_aoi21 _1626_ (
    .a(_0890_),
    .b(_0842_),
    .c(_0891_),
    .y(_0892_)
  );
  al_oa21ftt _1627_ (
    .a(_0890_),
    .b(_0847_),
    .c(_0892_),
    .y(_0893_)
  );
  al_ao21ftt _1628_ (
    .a(_0889_),
    .b(_0888_),
    .c(_0893_),
    .y(_0894_)
  );
  al_aoi21ttf _1629_ (
    .a(_0887_),
    .b(_0894_),
    .c(_0885_),
    .y(N10101)
  );
  al_nand2 _1630_ (
    .a(N245),
    .b(N271),
    .y(_0895_)
  );
  al_and3ftt _1631_ (
    .a(N38),
    .b(N382),
    .c(_0895_),
    .y(_0896_)
  );
  al_or2 _1632_ (
    .a(_0646_),
    .b(_0461_),
    .y(_0897_)
  );
  al_and2 _1633_ (
    .a(_0634_),
    .b(_0465_),
    .y(_0898_)
  );
  al_or2 _1634_ (
    .a(N70),
    .b(N89),
    .y(_0899_)
  );
  al_nand3ftt _1635_ (
    .a(N18),
    .b(N41),
    .c(_0899_),
    .y(_0900_)
  );
  al_aoi21ttf _1636_ (
    .a(N89),
    .b(_0436_),
    .c(_0900_),
    .y(_0901_)
  );
  al_ao21ttf _1637_ (
    .a(_0443_),
    .b(_0629_),
    .c(_0901_),
    .y(_0902_)
  );
  al_or2 _1638_ (
    .a(_0629_),
    .b(_0443_),
    .y(_0903_)
  );
  al_oa21 _1639_ (
    .a(_0435_),
    .b(_0630_),
    .c(_0903_),
    .y(_0904_)
  );
  al_nand2 _1640_ (
    .a(_0630_),
    .b(_0435_),
    .y(_0905_)
  );
  al_ao21ttf _1641_ (
    .a(_0463_),
    .b(_0633_),
    .c(_0905_),
    .y(_0906_)
  );
  al_ao21 _1642_ (
    .a(_0902_),
    .b(_0904_),
    .c(_0906_),
    .y(_0907_)
  );
  al_or2 _1643_ (
    .a(_0634_),
    .b(_0465_),
    .y(_0908_)
  );
  al_oa21 _1644_ (
    .a(_0463_),
    .b(_0633_),
    .c(_0908_),
    .y(_0909_)
  );
  al_ao21 _1645_ (
    .a(_0909_),
    .b(_0907_),
    .c(_0898_),
    .y(_0910_)
  );
  al_nand2 _1646_ (
    .a(_0646_),
    .b(_0461_),
    .y(_0911_)
  );
  al_ao21ftf _1647_ (
    .a(_0456_),
    .b(_0647_),
    .c(_0911_),
    .y(_0912_)
  );
  al_ao21 _1648_ (
    .a(_0897_),
    .b(_0910_),
    .c(_0912_),
    .y(_0913_)
  );
  al_or2 _1649_ (
    .a(_0643_),
    .b(_0452_),
    .y(_0914_)
  );
  al_nand2 _1650_ (
    .a(_0642_),
    .b(_0450_),
    .y(_0915_)
  );
  al_nand2ft _1651_ (
    .a(_0647_),
    .b(_0456_),
    .y(_0916_)
  );
  al_oa21 _1652_ (
    .a(_0450_),
    .b(_0642_),
    .c(_0916_),
    .y(_0917_)
  );
  al_and3 _1653_ (
    .a(_0914_),
    .b(_0915_),
    .c(_0917_),
    .y(_0918_)
  );
  al_nand2 _1654_ (
    .a(_0643_),
    .b(_0452_),
    .y(_0919_)
  );
  al_aoi21ttf _1655_ (
    .a(_0549_),
    .b(_0616_),
    .c(_0919_),
    .y(_0920_)
  );
  al_ao21ftf _1656_ (
    .a(_0915_),
    .b(_0914_),
    .c(_0920_),
    .y(_0921_)
  );
  al_ao21 _1657_ (
    .a(_0918_),
    .b(_0913_),
    .c(_0921_),
    .y(_0922_)
  );
  al_nand2 _1658_ (
    .a(_0610_),
    .b(_0516_),
    .y(_0923_)
  );
  al_aoi21ttf _1659_ (
    .a(_0518_),
    .b(_0611_),
    .c(_0923_),
    .y(_0924_)
  );
  al_or2 _1660_ (
    .a(_0593_),
    .b(_0533_),
    .y(_0925_)
  );
  al_or2 _1661_ (
    .a(_0610_),
    .b(_0516_),
    .y(_0926_)
  );
  al_oa21 _1662_ (
    .a(_0518_),
    .b(_0611_),
    .c(_0926_),
    .y(_0927_)
  );
  al_and3 _1663_ (
    .a(_0925_),
    .b(_0924_),
    .c(_0927_),
    .y(_0928_)
  );
  al_nand2 _1664_ (
    .a(_0592_),
    .b(_0531_),
    .y(_0929_)
  );
  al_ao21ttf _1665_ (
    .a(_0533_),
    .b(_0593_),
    .c(_0929_),
    .y(_0930_)
  );
  al_nor2 _1666_ (
    .a(_0592_),
    .b(_0531_),
    .y(_0931_)
  );
  al_oai21ttf _1667_ (
    .a(_0549_),
    .b(_0616_),
    .c(_0931_),
    .y(_0932_)
  );
  al_and3fft _1668_ (
    .a(_0930_),
    .b(_0932_),
    .c(_0928_),
    .y(_0933_)
  );
  al_oai21ttf _1669_ (
    .a(_0518_),
    .b(_0611_),
    .c(_0924_),
    .y(_0934_)
  );
  al_ao21ttf _1670_ (
    .a(_0930_),
    .b(_0928_),
    .c(_0934_),
    .y(_0935_)
  );
  al_ao21 _1671_ (
    .a(_0933_),
    .b(_0922_),
    .c(_0935_),
    .y(_0936_)
  );
  al_or2 _1672_ (
    .a(_0598_),
    .b(_0524_),
    .y(_0937_)
  );
  al_nand2 _1673_ (
    .a(_0597_),
    .b(_0522_),
    .y(_0938_)
  );
  al_nand2 _1674_ (
    .a(_0598_),
    .b(_0524_),
    .y(_0939_)
  );
  al_oa21 _1675_ (
    .a(_0522_),
    .b(_0597_),
    .c(_0939_),
    .y(_0940_)
  );
  al_and3 _1676_ (
    .a(_0937_),
    .b(_0938_),
    .c(_0940_),
    .y(_0941_)
  );
  al_nand2 _1677_ (
    .a(_0602_),
    .b(_0540_),
    .y(_0942_)
  );
  al_ao21ftf _1678_ (
    .a(_0542_),
    .b(_0603_),
    .c(_0942_),
    .y(_0943_)
  );
  al_nand2ft _1679_ (
    .a(_0603_),
    .b(_0542_),
    .y(_0944_)
  );
  al_nor2 _1680_ (
    .a(_0602_),
    .b(_0540_),
    .y(_0945_)
  );
  al_and3fft _1681_ (
    .a(_0945_),
    .b(_0943_),
    .c(_0944_),
    .y(_0946_)
  );
  al_nand3 _1682_ (
    .a(_0941_),
    .b(_0946_),
    .c(_0936_),
    .y(_0947_)
  );
  al_and2 _1683_ (
    .a(_0944_),
    .b(_0943_),
    .y(_0948_)
  );
  al_aoi21ttf _1684_ (
    .a(_0938_),
    .b(_0939_),
    .c(_0937_),
    .y(_0949_)
  );
  al_aoi21 _1685_ (
    .a(_0948_),
    .b(_0941_),
    .c(_0949_),
    .y(_0950_)
  );
  al_nor2 _1686_ (
    .a(_0476_),
    .b(_0675_),
    .y(_0951_)
  );
  al_and2 _1687_ (
    .a(_0674_),
    .b(_0474_),
    .y(_0952_)
  );
  al_or2 _1688_ (
    .a(_0674_),
    .b(_0474_),
    .y(_0953_)
  );
  al_aoi21ttf _1689_ (
    .a(_0476_),
    .b(_0675_),
    .c(_0953_),
    .y(_0954_)
  );
  al_nand3fft _1690_ (
    .a(_0951_),
    .b(_0952_),
    .c(_0954_),
    .y(_0955_)
  );
  al_nand2 _1691_ (
    .a(_0679_),
    .b(_0496_),
    .y(_0956_)
  );
  al_ao21ftf _1692_ (
    .a(_0507_),
    .b(_0678_),
    .c(_0956_),
    .y(_0957_)
  );
  al_or2 _1693_ (
    .a(_0679_),
    .b(_0496_),
    .y(_0958_)
  );
  al_aoi21ftf _1694_ (
    .a(_0678_),
    .b(_0507_),
    .c(_0958_),
    .y(_0959_)
  );
  al_and3fft _1695_ (
    .a(_0957_),
    .b(_0955_),
    .c(_0959_),
    .y(_0960_)
  );
  al_nand2 _1696_ (
    .a(_0662_),
    .b(_0492_),
    .y(_0961_)
  );
  al_or2 _1697_ (
    .a(_0662_),
    .b(_0492_),
    .y(_0962_)
  );
  al_nand3 _1698_ (
    .a(_0961_),
    .b(_0962_),
    .c(_0960_),
    .y(_0963_)
  );
  al_ao21 _1699_ (
    .a(_0950_),
    .b(_0947_),
    .c(_0963_),
    .y(_0964_)
  );
  al_or3fft _1700_ (
    .a(_0957_),
    .b(_0958_),
    .c(_0955_),
    .y(_0965_)
  );
  al_ao21ttf _1701_ (
    .a(_0476_),
    .b(_0675_),
    .c(_0952_),
    .y(_0966_)
  );
  al_and3ftt _1702_ (
    .a(_0951_),
    .b(_0966_),
    .c(_0965_),
    .y(_0967_)
  );
  al_aoi21ftf _1703_ (
    .a(_0961_),
    .b(_0960_),
    .c(_0967_),
    .y(_0968_)
  );
  al_nand3 _1704_ (
    .a(_0346_),
    .b(_0658_),
    .c(_0481_),
    .y(_0969_)
  );
  al_nand3 _1705_ (
    .a(_0346_),
    .b(_0657_),
    .c(_0483_),
    .y(_0970_)
  );
  al_aoi21 _1706_ (
    .a(_0346_),
    .b(_0657_),
    .c(_0483_),
    .y(_0000_)
  );
  al_oa21ttf _1707_ (
    .a(_0481_),
    .b(_0656_),
    .c(_0000_),
    .y(_0001_)
  );
  al_and3 _1708_ (
    .a(_0969_),
    .b(_0970_),
    .c(_0001_),
    .y(_0002_)
  );
  al_nand3 _1709_ (
    .a(_0346_),
    .b(_0666_),
    .c(_0503_),
    .y(_0003_)
  );
  al_aoi21ttf _1710_ (
    .a(_0501_),
    .b(_0665_),
    .c(_0003_),
    .y(_0004_)
  );
  al_ao21 _1711_ (
    .a(_0346_),
    .b(_0666_),
    .c(_0503_),
    .y(_0005_)
  );
  al_oa21 _1712_ (
    .a(_0501_),
    .b(_0665_),
    .c(_0005_),
    .y(_0006_)
  );
  al_and3 _1713_ (
    .a(_0004_),
    .b(_0006_),
    .c(_0002_),
    .y(_0007_)
  );
  al_ao21ttf _1714_ (
    .a(_0968_),
    .b(_0964_),
    .c(_0007_),
    .y(_0008_)
  );
  al_nor2ft _1715_ (
    .a(_0005_),
    .b(_0004_),
    .y(_0009_)
  );
  al_aoi21 _1716_ (
    .a(_0970_),
    .b(_0969_),
    .c(_0000_),
    .y(_0010_)
  );
  al_aoi21 _1717_ (
    .a(_0009_),
    .b(_0002_),
    .c(_0010_),
    .y(_0011_)
  );
  al_ao21 _1718_ (
    .a(_0346_),
    .b(_0691_),
    .c(_0568_),
    .y(_0012_)
  );
  al_and3 _1719_ (
    .a(_0346_),
    .b(_0691_),
    .c(_0568_),
    .y(_0013_)
  );
  al_nand2ft _1720_ (
    .a(_0013_),
    .b(_0012_),
    .y(_0014_)
  );
  al_ao21 _1721_ (
    .a(_0346_),
    .b(_0699_),
    .c(_0576_),
    .y(_0015_)
  );
  al_and3 _1722_ (
    .a(_0346_),
    .b(_0689_),
    .c(_0566_),
    .y(_0016_)
  );
  al_ao21 _1723_ (
    .a(_0346_),
    .b(_0689_),
    .c(_0566_),
    .y(_0017_)
  );
  al_nand2ft _1724_ (
    .a(_0016_),
    .b(_0017_),
    .y(_0018_)
  );
  al_nor3ftt _1725_ (
    .a(_0015_),
    .b(_0014_),
    .c(_0018_),
    .y(_0019_)
  );
  al_nand2 _1726_ (
    .a(_0346_),
    .b(_0561_),
    .y(_0020_)
  );
  al_aoi21ttf _1727_ (
    .a(_0574_),
    .b(_0698_),
    .c(_0020_),
    .y(_0021_)
  );
  al_or3fft _1728_ (
    .a(N12),
    .b(N9),
    .c(_0561_),
    .y(_0022_)
  );
  al_and3 _1729_ (
    .a(_0346_),
    .b(_0699_),
    .c(_0576_),
    .y(_0023_)
  );
  al_ao21 _1730_ (
    .a(_0346_),
    .b(_0697_),
    .c(_0574_),
    .y(_0024_)
  );
  al_and3ftt _1731_ (
    .a(_0023_),
    .b(_0022_),
    .c(_0024_),
    .y(_0025_)
  );
  al_nand3 _1732_ (
    .a(_0021_),
    .b(_0025_),
    .c(_0019_),
    .y(_0026_)
  );
  al_ao21 _1733_ (
    .a(_0011_),
    .b(_0008_),
    .c(_0026_),
    .y(_0027_)
  );
  al_oai21ftf _1734_ (
    .a(_0024_),
    .b(_0021_),
    .c(_0023_),
    .y(_0028_)
  );
  al_aoi21ttf _1735_ (
    .a(N382),
    .b(_0582_),
    .c(N38),
    .y(_0029_)
  );
  al_nand3ftt _1736_ (
    .a(_0690_),
    .b(_0566_),
    .c(_0012_),
    .y(_0030_)
  );
  al_nand3fft _1737_ (
    .a(_0013_),
    .b(_0029_),
    .c(_0030_),
    .y(_0031_)
  );
  al_aoi21 _1738_ (
    .a(_0028_),
    .b(_0019_),
    .c(_0031_),
    .y(_0032_)
  );
  al_aoi21 _1739_ (
    .a(_0032_),
    .b(_0027_),
    .c(_0896_),
    .y(N10102)
  );
  al_and2ft _1740_ (
    .a(_0749_),
    .b(_0761_),
    .y(_0033_)
  );
  al_and3 _1741_ (
    .a(_0760_),
    .b(_0033_),
    .c(_0763_),
    .y(_0034_)
  );
  al_nand3 _1742_ (
    .a(_0034_),
    .b(_0755_),
    .c(_0759_),
    .y(_0035_)
  );
  al_and3 _1743_ (
    .a(_0751_),
    .b(_0764_),
    .c(_0035_),
    .y(_0036_)
  );
  al_ao21 _1744_ (
    .a(_0751_),
    .b(_0035_),
    .c(_0764_),
    .y(_0037_)
  );
  al_nand2ft _1745_ (
    .a(_0036_),
    .b(_0037_),
    .y(N10350)
  );
  al_nand3 _1746_ (
    .a(_0761_),
    .b(_0755_),
    .c(_0759_),
    .y(_0038_)
  );
  al_oa21ftf _1747_ (
    .a(_0760_),
    .b(_0038_),
    .c(_0750_),
    .y(_0039_)
  );
  al_and2 _1748_ (
    .a(_0763_),
    .b(_0039_),
    .y(_0040_)
  );
  al_or2 _1749_ (
    .a(_0763_),
    .b(_0039_),
    .y(_0041_)
  );
  al_nand2ft _1750_ (
    .a(_0040_),
    .b(_0041_),
    .y(N10351)
  );
  al_and3ftt _1751_ (
    .a(_0749_),
    .b(_0760_),
    .c(_0038_),
    .y(_0042_)
  );
  al_inv _1752_ (
    .a(_0760_),
    .y(_0043_)
  );
  al_ao21ftf _1753_ (
    .a(_0749_),
    .b(_0038_),
    .c(_0043_),
    .y(_0044_)
  );
  al_nand2ft _1754_ (
    .a(_0042_),
    .b(_0044_),
    .y(N10352)
  );
  al_and3ftt _1755_ (
    .a(_0033_),
    .b(_0755_),
    .c(_0759_),
    .y(_0045_)
  );
  al_ao21ttf _1756_ (
    .a(_0755_),
    .b(_0759_),
    .c(_0033_),
    .y(_0046_)
  );
  al_nand2ft _1757_ (
    .a(_0045_),
    .b(_0046_),
    .y(N10353)
  );
  al_nand2 _1758_ (
    .a(_0950_),
    .b(_0947_),
    .y(N10704)
  );
  al_oai21ftf _1759_ (
    .a(_0783_),
    .b(_0789_),
    .c(_0815_),
    .y(_0047_)
  );
  al_nand2 _1760_ (
    .a(_0807_),
    .b(_0808_),
    .y(_0048_)
  );
  al_ao21ftf _1761_ (
    .a(_0815_),
    .b(_0048_),
    .c(_0047_),
    .y(_0049_)
  );
  al_or2 _1762_ (
    .a(_0812_),
    .b(_0049_),
    .y(_0050_)
  );
  al_and2 _1763_ (
    .a(_0812_),
    .b(_0049_),
    .y(_0051_)
  );
  al_nand2ft _1764_ (
    .a(_0051_),
    .b(_0050_),
    .y(N10760)
  );
  al_inv _1765_ (
    .a(_0783_),
    .y(_0052_)
  );
  al_and3fft _1766_ (
    .a(_0052_),
    .b(_0809_),
    .c(_0814_),
    .y(_0053_)
  );
  al_oai21ftf _1767_ (
    .a(_0814_),
    .b(_0809_),
    .c(_0783_),
    .y(_0054_)
  );
  al_nand2ft _1768_ (
    .a(_0053_),
    .b(_0054_),
    .y(N10761)
  );
  al_and2 _1769_ (
    .a(_0787_),
    .b(_0785_),
    .y(_0055_)
  );
  al_nand3 _1770_ (
    .a(_0786_),
    .b(_0807_),
    .c(_0808_),
    .y(_0056_)
  );
  al_and3 _1771_ (
    .a(_0784_),
    .b(_0055_),
    .c(_0056_),
    .y(_0057_)
  );
  al_ao21 _1772_ (
    .a(_0784_),
    .b(_0056_),
    .c(_0055_),
    .y(_0058_)
  );
  al_nand2ft _1773_ (
    .a(_0057_),
    .b(_0058_),
    .y(N10762)
  );
  al_ao21ttf _1774_ (
    .a(_0786_),
    .b(_0784_),
    .c(_0048_),
    .y(_0059_)
  );
  al_aoi21ftf _1775_ (
    .a(_0056_),
    .b(_0784_),
    .c(_0059_),
    .y(N10763)
  );
  al_or2ft _1776_ (
    .a(_0885_),
    .b(_0886_),
    .y(_0060_)
  );
  al_nand3ftt _1777_ (
    .a(N38),
    .b(N263),
    .c(N382),
    .y(_0061_)
  );
  al_or3fft _1778_ (
    .a(_0854_),
    .b(_0851_),
    .c(_0847_),
    .y(_0062_)
  );
  al_ao21ttf _1779_ (
    .a(N263),
    .b(N382),
    .c(N38),
    .y(_0063_)
  );
  al_nand3 _1780_ (
    .a(_0892_),
    .b(_0063_),
    .c(_0062_),
    .y(_0064_)
  );
  al_and3 _1781_ (
    .a(_0060_),
    .b(_0061_),
    .c(_0064_),
    .y(_0065_)
  );
  al_ao21 _1782_ (
    .a(_0061_),
    .b(_0064_),
    .c(_0060_),
    .y(_0066_)
  );
  al_nand2ft _1783_ (
    .a(_0065_),
    .b(_0066_),
    .y(N10837)
  );
  al_and3ftt _1784_ (
    .a(_0889_),
    .b(_0888_),
    .c(_0893_),
    .y(_0067_)
  );
  al_and2ft _1785_ (
    .a(_0067_),
    .b(_0894_),
    .y(N10839)
  );
  al_nand2 _1786_ (
    .a(_0714_),
    .b(_0715_),
    .y(_0068_)
  );
  al_ao21ftf _1787_ (
    .a(_0727_),
    .b(_0773_),
    .c(_0068_),
    .y(_0069_)
  );
  al_oa21ftt _1788_ (
    .a(_0714_),
    .b(_0774_),
    .c(_0069_),
    .y(N10905)
  );
  al_nand2ft _1789_ (
    .a(_0718_),
    .b(_0717_),
    .y(_0070_)
  );
  al_nand2 _1790_ (
    .a(_0772_),
    .b(_0767_),
    .y(_0071_)
  );
  al_aoi21ttf _1791_ (
    .a(_0726_),
    .b(_0071_),
    .c(_0722_),
    .y(_0072_)
  );
  al_and2ft _1792_ (
    .a(_0070_),
    .b(_0072_),
    .y(_0073_)
  );
  al_or2ft _1793_ (
    .a(_0070_),
    .b(_0072_),
    .y(_0074_)
  );
  al_nand2ft _1794_ (
    .a(_0073_),
    .b(_0074_),
    .y(N10906)
  );
  al_inv _1795_ (
    .a(_0724_),
    .y(_0075_)
  );
  al_and3 _1796_ (
    .a(_0721_),
    .b(_0772_),
    .c(_0767_),
    .y(_0076_)
  );
  al_and3fft _1797_ (
    .a(_0725_),
    .b(_0076_),
    .c(_0075_),
    .y(_0077_)
  );
  al_inv _1798_ (
    .a(_0725_),
    .y(_0078_)
  );
  al_oai21ftf _1799_ (
    .a(_0078_),
    .b(_0076_),
    .c(_0075_),
    .y(_0079_)
  );
  al_nand2ft _1800_ (
    .a(_0077_),
    .b(_0079_),
    .y(N10907)
  );
  al_ao21ftf _1801_ (
    .a(_0725_),
    .b(_0721_),
    .c(_0071_),
    .y(_0080_)
  );
  al_ao21ftf _1802_ (
    .a(_0725_),
    .b(_0076_),
    .c(_0080_),
    .y(N10908)
  );
  al_oai21ftf _1803_ (
    .a(_0826_),
    .b(_0820_),
    .c(_0800_),
    .y(_0081_)
  );
  al_oa21 _1804_ (
    .a(_0797_),
    .b(_0798_),
    .c(_0713_),
    .y(_0082_)
  );
  al_and3ftt _1805_ (
    .a(_0082_),
    .b(_0820_),
    .c(_0801_),
    .y(_0083_)
  );
  al_ao21ftt _1806_ (
    .a(_0082_),
    .b(_0820_),
    .c(_0801_),
    .y(_0084_)
  );
  al_nor3fft _1807_ (
    .a(_0806_),
    .b(_0084_),
    .c(_0083_),
    .y(_0085_)
  );
  al_nand3ftt _1808_ (
    .a(_0368_),
    .b(N280),
    .c(_0712_),
    .y(_0086_)
  );
  al_aoi21ftf _1809_ (
    .a(_0712_),
    .b(_0797_),
    .c(_0086_),
    .y(_0087_)
  );
  al_oa21 _1810_ (
    .a(_0791_),
    .b(_0792_),
    .c(_0087_),
    .y(_0088_)
  );
  al_or3 _1811_ (
    .a(_0791_),
    .b(_0792_),
    .c(_0087_),
    .y(_0089_)
  );
  al_nand3ftt _1812_ (
    .a(_0088_),
    .b(_0089_),
    .c(_0085_),
    .y(_0090_)
  );
  al_ao21ftt _1813_ (
    .a(_0088_),
    .b(_0089_),
    .c(_0085_),
    .y(_0091_)
  );
  al_ao21 _1814_ (
    .a(_0090_),
    .b(_0091_),
    .c(_0081_),
    .y(_0092_)
  );
  al_nand3 _1815_ (
    .a(_0081_),
    .b(_0090_),
    .c(_0091_),
    .y(_0093_)
  );
  al_nand3 _1816_ (
    .a(_0092_),
    .b(_0093_),
    .c(_0825_),
    .y(_0094_)
  );
  al_mux2h _1817_ (
    .a(_0797_),
    .b(_0798_),
    .s(_0711_),
    .y(_0095_)
  );
  al_oai21 _1818_ (
    .a(_0792_),
    .b(_0791_),
    .c(_0095_),
    .y(_0096_)
  );
  al_or3 _1819_ (
    .a(_0792_),
    .b(_0791_),
    .c(_0095_),
    .y(_0097_)
  );
  al_or3fft _1820_ (
    .a(_0097_),
    .b(_0096_),
    .c(_0800_),
    .y(_0098_)
  );
  al_aoi21ttf _1821_ (
    .a(_0097_),
    .b(_0096_),
    .c(_0800_),
    .y(_0099_)
  );
  al_nand2ft _1822_ (
    .a(_0099_),
    .b(_0098_),
    .y(_0100_)
  );
  al_oai21ftf _1823_ (
    .a(_0084_),
    .b(_0083_),
    .c(_0100_),
    .y(_0101_)
  );
  al_nand3ftt _1824_ (
    .a(_0083_),
    .b(_0084_),
    .c(_0100_),
    .y(_0102_)
  );
  al_or3fft _1825_ (
    .a(_0101_),
    .b(_0102_),
    .c(_0825_),
    .y(_0103_)
  );
  al_ao21ftt _1826_ (
    .a(_0795_),
    .b(_0796_),
    .c(_0804_),
    .y(_0104_)
  );
  al_and2ft _1827_ (
    .a(_0805_),
    .b(_0104_),
    .y(_0105_)
  );
  al_ao21 _1828_ (
    .a(_0094_),
    .b(_0103_),
    .c(_0105_),
    .y(_0106_)
  );
  al_nand3 _1829_ (
    .a(_0105_),
    .b(_0094_),
    .c(_0103_),
    .y(_0107_)
  );
  al_mux2l _1830_ (
    .a(_0782_),
    .b(_0781_),
    .s(_0814_),
    .y(_0108_)
  );
  al_oai21ttf _1831_ (
    .a(_0786_),
    .b(_0055_),
    .c(_0788_),
    .y(_0109_)
  );
  al_oai21 _1832_ (
    .a(_0781_),
    .b(_0782_),
    .c(_0812_),
    .y(_0110_)
  );
  al_ao21ftf _1833_ (
    .a(_0811_),
    .b(_0810_),
    .c(_0783_),
    .y(_0111_)
  );
  al_nor3fft _1834_ (
    .a(_0111_),
    .b(_0110_),
    .c(_0109_),
    .y(_0112_)
  );
  al_ao21ttf _1835_ (
    .a(_0111_),
    .b(_0110_),
    .c(_0109_),
    .y(_0113_)
  );
  al_and3fft _1836_ (
    .a(_0108_),
    .b(_0112_),
    .c(_0113_),
    .y(_0114_)
  );
  al_oai21ftt _1837_ (
    .a(_0113_),
    .b(_0112_),
    .c(_0108_),
    .y(_0115_)
  );
  al_nand2ft _1838_ (
    .a(_0114_),
    .b(_0115_),
    .y(_0116_)
  );
  al_mux2h _1839_ (
    .a(_0787_),
    .b(_0785_),
    .s(_0786_),
    .y(_0117_)
  );
  al_oa21ttf _1840_ (
    .a(_0781_),
    .b(_0782_),
    .c(_0117_),
    .y(_0118_)
  );
  al_nand3fft _1841_ (
    .a(_0781_),
    .b(_0782_),
    .c(_0117_),
    .y(_0119_)
  );
  al_or2ft _1842_ (
    .a(_0119_),
    .b(_0118_),
    .y(_0120_)
  );
  al_ao21 _1843_ (
    .a(_0786_),
    .b(_0784_),
    .c(_0055_),
    .y(_0121_)
  );
  al_nand3 _1844_ (
    .a(_0812_),
    .b(_0789_),
    .c(_0121_),
    .y(_0122_)
  );
  al_ao21 _1845_ (
    .a(_0789_),
    .b(_0121_),
    .c(_0812_),
    .y(_0123_)
  );
  al_aoi21ttf _1846_ (
    .a(_0122_),
    .b(_0123_),
    .c(_0047_),
    .y(_0124_)
  );
  al_or3fft _1847_ (
    .a(_0122_),
    .b(_0123_),
    .c(_0047_),
    .y(_0125_)
  );
  al_nor3fft _1848_ (
    .a(_0120_),
    .b(_0125_),
    .c(_0124_),
    .y(_0126_)
  );
  al_oai21ftf _1849_ (
    .a(_0125_),
    .b(_0124_),
    .c(_0120_),
    .y(_0127_)
  );
  al_nand2ft _1850_ (
    .a(_0126_),
    .b(_0127_),
    .y(_0128_)
  );
  al_mux2l _1851_ (
    .a(_0116_),
    .b(_0128_),
    .s(_0048_),
    .y(_0129_)
  );
  al_aoi21 _1852_ (
    .a(_0107_),
    .b(_0106_),
    .c(_0129_),
    .y(_0130_)
  );
  al_nand3 _1853_ (
    .a(_0107_),
    .b(_0106_),
    .c(_0129_),
    .y(_0131_)
  );
  al_nand2ft _1854_ (
    .a(_0130_),
    .b(_0131_),
    .y(N11333)
  );
  al_nand3ftt _1855_ (
    .a(_0889_),
    .b(_0892_),
    .c(_0062_),
    .y(_0132_)
  );
  al_ao21ftf _1856_ (
    .a(_0835_),
    .b(_0836_),
    .c(_0844_),
    .y(_0133_)
  );
  al_aoi21ftf _1857_ (
    .a(_0837_),
    .b(_0838_),
    .c(_0854_),
    .y(_0134_)
  );
  al_nand2ft _1858_ (
    .a(_0134_),
    .b(_0133_),
    .y(_0135_)
  );
  al_and3 _1859_ (
    .a(N267),
    .b(N382),
    .c(_0135_),
    .y(_0136_)
  );
  al_ao21 _1860_ (
    .a(N267),
    .b(N382),
    .c(_0135_),
    .y(_0137_)
  );
  al_nand2ft _1861_ (
    .a(_0136_),
    .b(_0137_),
    .y(_0138_)
  );
  al_nand3 _1862_ (
    .a(_0777_),
    .b(_0778_),
    .c(_0845_),
    .y(_0139_)
  );
  al_aoi21 _1863_ (
    .a(_0777_),
    .b(_0778_),
    .c(_0845_),
    .y(_0140_)
  );
  al_nand3ftt _1864_ (
    .a(_0140_),
    .b(_0139_),
    .c(_0843_),
    .y(_0141_)
  );
  al_ao21ftt _1865_ (
    .a(_0140_),
    .b(_0139_),
    .c(_0843_),
    .y(_0142_)
  );
  al_or3fft _1866_ (
    .a(_0844_),
    .b(_0854_),
    .c(_0139_),
    .y(_0143_)
  );
  al_nand3 _1867_ (
    .a(_0143_),
    .b(_0141_),
    .c(_0142_),
    .y(_0144_)
  );
  al_nand3fft _1868_ (
    .a(_0573_),
    .b(_0387_),
    .c(_0778_),
    .y(_0145_)
  );
  al_aoi21ftf _1869_ (
    .a(_0778_),
    .b(_0839_),
    .c(_0145_),
    .y(_0146_)
  );
  al_or3 _1870_ (
    .a(_0849_),
    .b(_0850_),
    .c(_0146_),
    .y(_0147_)
  );
  al_and2ft _1871_ (
    .a(_0851_),
    .b(_0146_),
    .y(_0148_)
  );
  al_nand2ft _1872_ (
    .a(_0148_),
    .b(_0147_),
    .y(_0149_)
  );
  al_aoi21ftt _1873_ (
    .a(_0842_),
    .b(_0846_),
    .c(_0149_),
    .y(_0150_)
  );
  al_nand3ftt _1874_ (
    .a(_0842_),
    .b(_0846_),
    .c(_0149_),
    .y(_0151_)
  );
  al_or3ftt _1875_ (
    .a(_0151_),
    .b(_0150_),
    .c(_0144_),
    .y(_0152_)
  );
  al_aoi21ftf _1876_ (
    .a(_0150_),
    .b(_0151_),
    .c(_0144_),
    .y(_0153_)
  );
  al_nand2ft _1877_ (
    .a(_0153_),
    .b(_0152_),
    .y(_0154_)
  );
  al_ao21 _1878_ (
    .a(_0816_),
    .b(_0813_),
    .c(_0154_),
    .y(_0155_)
  );
  al_mux2l _1879_ (
    .a(_0839_),
    .b(_0840_),
    .s(_0777_),
    .y(_0156_)
  );
  al_nand3fft _1880_ (
    .a(_0849_),
    .b(_0850_),
    .c(_0156_),
    .y(_0157_)
  );
  al_oai21ttf _1881_ (
    .a(_0849_),
    .b(_0850_),
    .c(_0156_),
    .y(_0158_)
  );
  al_aoi21ttf _1882_ (
    .a(_0157_),
    .b(_0158_),
    .c(_0842_),
    .y(_0159_)
  );
  al_or3fft _1883_ (
    .a(_0157_),
    .b(_0158_),
    .c(_0842_),
    .y(_0160_)
  );
  al_nand2ft _1884_ (
    .a(_0159_),
    .b(_0160_),
    .y(_0161_)
  );
  al_or3fft _1885_ (
    .a(_0141_),
    .b(_0142_),
    .c(_0161_),
    .y(_0162_)
  );
  al_aoi21ttf _1886_ (
    .a(_0141_),
    .b(_0142_),
    .c(_0161_),
    .y(_0163_)
  );
  al_and2ft _1887_ (
    .a(_0163_),
    .b(_0162_),
    .y(_0164_)
  );
  al_nand3 _1888_ (
    .a(_0816_),
    .b(_0164_),
    .c(_0813_),
    .y(_0165_)
  );
  al_and3 _1889_ (
    .a(_0138_),
    .b(_0165_),
    .c(_0155_),
    .y(_0166_)
  );
  al_ao21 _1890_ (
    .a(_0165_),
    .b(_0155_),
    .c(_0138_),
    .y(_0167_)
  );
  al_nand2ft _1891_ (
    .a(_0166_),
    .b(_0167_),
    .y(_0168_)
  );
  al_ao21 _1892_ (
    .a(_0888_),
    .b(_0132_),
    .c(_0168_),
    .y(_0169_)
  );
  al_and3 _1893_ (
    .a(_0888_),
    .b(_0132_),
    .c(_0168_),
    .y(_0170_)
  );
  al_nand2ft _1894_ (
    .a(_0170_),
    .b(_0169_),
    .y(N11334)
  );
  al_ao21ftf _1895_ (
    .a(N358),
    .b(_0422_),
    .c(_0721_),
    .y(_0171_)
  );
  al_ao21 _1896_ (
    .a(_0719_),
    .b(_0725_),
    .c(_0171_),
    .y(_0172_)
  );
  al_aoi21ftf _1897_ (
    .a(_0721_),
    .b(_0720_),
    .c(_0172_),
    .y(_0173_)
  );
  al_and3 _1898_ (
    .a(_0715_),
    .b(_0714_),
    .c(_0070_),
    .y(_0174_)
  );
  al_nand3ftt _1899_ (
    .a(_0718_),
    .b(_0717_),
    .c(_0068_),
    .y(_0175_)
  );
  al_oai21ftt _1900_ (
    .a(_0175_),
    .b(_0174_),
    .c(_0173_),
    .y(_0176_)
  );
  al_or3ftt _1901_ (
    .a(_0175_),
    .b(_0174_),
    .c(_0173_),
    .y(_0177_)
  );
  al_and3 _1902_ (
    .a(_0727_),
    .b(_0176_),
    .c(_0177_),
    .y(_0178_)
  );
  al_ao21 _1903_ (
    .a(_0176_),
    .b(_0177_),
    .c(_0727_),
    .y(_0179_)
  );
  al_nand2ft _1904_ (
    .a(_0178_),
    .b(_0179_),
    .y(_0180_)
  );
  al_ao21 _1905_ (
    .a(_0717_),
    .b(_0722_),
    .c(_0718_),
    .y(_0181_)
  );
  al_and3fft _1906_ (
    .a(_0421_),
    .b(_0720_),
    .c(N355),
    .y(_0182_)
  );
  al_oai21ttf _1907_ (
    .a(_0725_),
    .b(_0722_),
    .c(_0182_),
    .y(_0183_)
  );
  al_aoi21ftf _1908_ (
    .a(_0720_),
    .b(_0719_),
    .c(_0068_),
    .y(_0184_)
  );
  al_nand3 _1909_ (
    .a(_0715_),
    .b(_0714_),
    .c(_0724_),
    .y(_0185_)
  );
  al_and3ftt _1910_ (
    .a(_0184_),
    .b(_0185_),
    .c(_0183_),
    .y(_0186_)
  );
  al_oai21ftf _1911_ (
    .a(_0185_),
    .b(_0184_),
    .c(_0183_),
    .y(_0187_)
  );
  al_oai21ftf _1912_ (
    .a(_0187_),
    .b(_0186_),
    .c(_0181_),
    .y(_0188_)
  );
  al_nor3fft _1913_ (
    .a(_0181_),
    .b(_0187_),
    .c(_0186_),
    .y(_0189_)
  );
  al_and2ft _1914_ (
    .a(_0189_),
    .b(_0188_),
    .y(_0190_)
  );
  al_mux2l _1915_ (
    .a(_0180_),
    .b(_0190_),
    .s(_0071_),
    .y(_0191_)
  );
  al_mux2h _1916_ (
    .a(_0741_),
    .b(_0875_),
    .s(_0871_),
    .y(_0192_)
  );
  al_and3 _1917_ (
    .a(_0548_),
    .b(_0413_),
    .c(_0733_),
    .y(_0193_)
  );
  al_aoi21 _1918_ (
    .a(_0734_),
    .b(_0732_),
    .c(_0193_),
    .y(_0194_)
  );
  al_ao21ttf _1919_ (
    .a(_0738_),
    .b(_0770_),
    .c(_0194_),
    .y(_0195_)
  );
  al_and3ftt _1920_ (
    .a(_0194_),
    .b(_0738_),
    .c(_0770_),
    .y(_0196_)
  );
  al_or3ftt _1921_ (
    .a(_0195_),
    .b(_0196_),
    .c(_0192_),
    .y(_0197_)
  );
  al_ao21ftf _1922_ (
    .a(_0196_),
    .b(_0195_),
    .c(_0192_),
    .y(_0198_)
  );
  al_ao21ttf _1923_ (
    .a(_0198_),
    .b(_0197_),
    .c(_0866_),
    .y(_0199_)
  );
  al_mux2l _1924_ (
    .a(_0736_),
    .b(_0735_),
    .s(_0769_),
    .y(_0200_)
  );
  al_ao21 _1925_ (
    .a(_0733_),
    .b(_0768_),
    .c(_0865_),
    .y(_0201_)
  );
  al_and3 _1926_ (
    .a(_0869_),
    .b(_0201_),
    .c(_0200_),
    .y(_0202_)
  );
  al_ao21 _1927_ (
    .a(_0869_),
    .b(_0201_),
    .c(_0200_),
    .y(_0203_)
  );
  al_or3ftt _1928_ (
    .a(_0203_),
    .b(_0202_),
    .c(_0875_),
    .y(_0204_)
  );
  al_ao21ftf _1929_ (
    .a(_0202_),
    .b(_0203_),
    .c(_0875_),
    .y(_0205_)
  );
  al_ao21 _1930_ (
    .a(_0205_),
    .b(_0204_),
    .c(_0866_),
    .y(_0206_)
  );
  al_oa21 _1931_ (
    .a(_0735_),
    .b(_0736_),
    .c(_0730_),
    .y(_0207_)
  );
  al_or2 _1932_ (
    .a(_0207_),
    .b(_0870_),
    .y(_0208_)
  );
  al_inv _1933_ (
    .a(_0208_),
    .y(_0209_)
  );
  al_ao21 _1934_ (
    .a(_0206_),
    .b(_0199_),
    .c(_0209_),
    .y(_0210_)
  );
  al_nand3 _1935_ (
    .a(_0206_),
    .b(_0209_),
    .c(_0199_),
    .y(_0211_)
  );
  al_aoi21ttf _1936_ (
    .a(_0211_),
    .b(_0210_),
    .c(_0191_),
    .y(_0212_)
  );
  al_and3ftt _1937_ (
    .a(_0191_),
    .b(_0211_),
    .c(_0210_),
    .y(_0213_)
  );
  al_or2 _1938_ (
    .a(_0213_),
    .b(_0212_),
    .y(N11340)
  );
  al_oai21 _1939_ (
    .a(_0745_),
    .b(_0746_),
    .c(_0760_),
    .y(_0214_)
  );
  al_ao21ftf _1940_ (
    .a(_0748_),
    .b(_0747_),
    .c(_0763_),
    .y(_0215_)
  );
  al_aoi21ttf _1941_ (
    .a(_0215_),
    .b(_0214_),
    .c(_0751_),
    .y(_0216_)
  );
  al_or3fft _1942_ (
    .a(_0215_),
    .b(_0214_),
    .c(_0751_),
    .y(_0217_)
  );
  al_nand2ft _1943_ (
    .a(_0216_),
    .b(_0217_),
    .y(_0218_)
  );
  al_inv _1944_ (
    .a(_0748_),
    .y(_0219_)
  );
  al_mux2h _1945_ (
    .a(_0219_),
    .b(_0750_),
    .s(_0761_),
    .y(_0220_)
  );
  al_nor2 _1946_ (
    .a(_0764_),
    .b(_0220_),
    .y(_0221_)
  );
  al_nand2 _1947_ (
    .a(_0764_),
    .b(_0220_),
    .y(_0222_)
  );
  al_ao21ftt _1948_ (
    .a(_0221_),
    .b(_0222_),
    .c(_0218_),
    .y(_0223_)
  );
  al_nand3ftt _1949_ (
    .a(_0221_),
    .b(_0222_),
    .c(_0218_),
    .y(_0224_)
  );
  al_ao21 _1950_ (
    .a(_0224_),
    .b(_0223_),
    .c(_0759_),
    .y(_0225_)
  );
  al_nand3fft _1951_ (
    .a(_0745_),
    .b(_0746_),
    .c(_0764_),
    .y(_0226_)
  );
  al_aoi21ftt _1952_ (
    .a(_0744_),
    .b(_0743_),
    .c(_0763_),
    .y(_0227_)
  );
  al_nor2ft _1953_ (
    .a(_0226_),
    .b(_0227_),
    .y(_0228_)
  );
  al_mux2h _1954_ (
    .a(_0747_),
    .b(_0219_),
    .s(_0749_),
    .y(_0229_)
  );
  al_mux2l _1955_ (
    .a(_0763_),
    .b(_0229_),
    .s(_0762_),
    .y(_0230_)
  );
  al_aoi21ftt _1956_ (
    .a(_0762_),
    .b(_0229_),
    .c(_0751_),
    .y(_0231_)
  );
  al_ao21 _1957_ (
    .a(_0751_),
    .b(_0230_),
    .c(_0231_),
    .y(_0232_)
  );
  al_or2 _1958_ (
    .a(_0228_),
    .b(_0232_),
    .y(_0233_)
  );
  al_and2 _1959_ (
    .a(_0228_),
    .b(_0232_),
    .y(_0234_)
  );
  al_nand2ft _1960_ (
    .a(_0234_),
    .b(_0233_),
    .y(_0235_)
  );
  al_ao21ttf _1961_ (
    .a(_0759_),
    .b(_0235_),
    .c(_0225_),
    .y(_0236_)
  );
  al_ao21 _1962_ (
    .a(_0224_),
    .b(_0223_),
    .c(_0755_),
    .y(_0237_)
  );
  al_inv _1963_ (
    .a(N367),
    .y(_0238_)
  );
  al_ao21ftf _1964_ (
    .a(_0282_),
    .b(_0754_),
    .c(_0238_),
    .y(_0239_)
  );
  al_ao21ftf _1965_ (
    .a(_0239_),
    .b(_0235_),
    .c(_0237_),
    .y(_0240_)
  );
  al_aoi21 _1966_ (
    .a(N367),
    .b(_0236_),
    .c(_0240_),
    .y(_0241_)
  );
  al_ao21ttf _1967_ (
    .a(_0287_),
    .b(_0300_),
    .c(_0753_),
    .y(_0242_)
  );
  al_ao21ttf _1968_ (
    .a(_0277_),
    .b(_0297_),
    .c(_0298_),
    .y(_0243_)
  );
  al_nand2ft _1969_ (
    .a(_0278_),
    .b(_0277_),
    .y(_0244_)
  );
  al_ao21ttf _1970_ (
    .a(_0297_),
    .b(_0292_),
    .c(_0244_),
    .y(_0245_)
  );
  al_or3fft _1971_ (
    .a(_0294_),
    .b(_0245_),
    .c(_0304_),
    .y(_0246_)
  );
  al_ao21ttf _1972_ (
    .a(_0294_),
    .b(_0245_),
    .c(_0304_),
    .y(_0247_)
  );
  al_ao21 _1973_ (
    .a(_0247_),
    .b(_0246_),
    .c(_0243_),
    .y(_0248_)
  );
  al_nand3 _1974_ (
    .a(_0243_),
    .b(_0247_),
    .c(_0246_),
    .y(_0249_)
  );
  al_ao21 _1975_ (
    .a(_0249_),
    .b(_0248_),
    .c(_0242_),
    .y(_0250_)
  );
  al_nand3 _1976_ (
    .a(_0242_),
    .b(_0249_),
    .c(_0248_),
    .y(_0251_)
  );
  al_nand3 _1977_ (
    .a(_0238_),
    .b(_0251_),
    .c(_0250_),
    .y(_0252_)
  );
  al_nand3 _1978_ (
    .a(_0278_),
    .b(_0297_),
    .c(_0298_),
    .y(_0253_)
  );
  al_ao21ftf _1979_ (
    .a(_0278_),
    .b(_0292_),
    .c(_0253_),
    .y(_0254_)
  );
  al_ao21ttf _1980_ (
    .a(_0295_),
    .b(_0300_),
    .c(_0254_),
    .y(_0255_)
  );
  al_and3ftt _1981_ (
    .a(_0254_),
    .b(_0295_),
    .c(_0300_),
    .y(_0256_)
  );
  al_nand2ft _1982_ (
    .a(_0256_),
    .b(_0255_),
    .y(_0257_)
  );
  al_or3fft _1983_ (
    .a(_0246_),
    .b(_0247_),
    .c(_0758_),
    .y(_0258_)
  );
  al_ao21ttf _1984_ (
    .a(_0246_),
    .b(_0247_),
    .c(_0758_),
    .y(_0259_)
  );
  al_ao21 _1985_ (
    .a(_0258_),
    .b(_0259_),
    .c(_0257_),
    .y(_0260_)
  );
  al_nand3 _1986_ (
    .a(_0259_),
    .b(_0258_),
    .c(_0257_),
    .y(_0261_)
  );
  al_nand3 _1987_ (
    .a(N367),
    .b(_0261_),
    .c(_0260_),
    .y(_0262_)
  );
  al_ao21ftt _1988_ (
    .a(_0286_),
    .b(_0306_),
    .c(_0756_),
    .y(_0263_)
  );
  al_and3ftt _1989_ (
    .a(_0286_),
    .b(_0306_),
    .c(_0756_),
    .y(_0264_)
  );
  al_nand2ft _1990_ (
    .a(_0264_),
    .b(_0263_),
    .y(_0265_)
  );
  al_ao21 _1991_ (
    .a(_0252_),
    .b(_0262_),
    .c(_0265_),
    .y(_0266_)
  );
  al_and3 _1992_ (
    .a(_0265_),
    .b(_0252_),
    .c(_0262_),
    .y(_0267_)
  );
  al_ao21ftt _1993_ (
    .a(_0267_),
    .b(_0266_),
    .c(_0241_),
    .y(_0268_)
  );
  al_and3ftt _1994_ (
    .a(_0267_),
    .b(_0266_),
    .c(_0241_),
    .y(_0269_)
  );
  al_nand2ft _1995_ (
    .a(_0269_),
    .b(_0268_),
    .y(N11342)
  );
  al_aoi21ttf _1996_ (
    .a(_0887_),
    .b(_0894_),
    .c(_0885_),
    .y(N10104)
  );
  al_aoi21 _1997_ (
    .a(_0032_),
    .b(_0027_),
    .c(_0896_),
    .y(N10628)
  );
  al_aoi21ttf _1998_ (
    .a(_0887_),
    .b(_0894_),
    .c(_0885_),
    .y(N10706)
  );
  al_aoi21ttf _1999_ (
    .a(_0887_),
    .b(_0894_),
    .c(_0885_),
    .y(N10759)
  );
  assign N10103 = N10102;
  assign N10778 = N10837;
  assign N10781 = N10839;
  assign N10838 = N10837;
  assign N10840 = N10839;
  assign N1112 = N1110;
  assign N1114 = N1111;
  assign N1116 = N1;
  assign N1125 = N18;
  assign N1136 = N18;
  assign N1147 = N18;
  assign N1160 = N18;
  assign N1175 = N18;
  assign N1182 = N18;
  assign N1233 = N18;
  assign N1244 = N18;
  assign N1249 = N18;
  assign N1256 = N18;
  assign N1270 = N18;
  assign N1277 = N18;
  assign N1287 = N38;
  assign N1299 = N38;
  assign N1308 = N38;
  assign N1311 = N38;
  assign N1428 = N38;
  assign N1431 = N38;
  assign N1489 = N1113;
  assign N1490 = N1;
  assign N1828 = N260;
  assign N1829 = N257;
  assign N1830 = N254;
  assign N1833 = N251;
  assign N1840 = N260;
  assign N1841 = N257;
  assign N1842 = N254;
  assign N1843 = N251;
  assign N1867 = N303;
  assign N1868 = N299;
  assign N1869 = N296;
  assign N1870 = N289;
  assign N1871 = N286;
  assign N1872 = N283;
  assign N1873 = N280;
  assign N1874 = N293;
  assign N1875 = N277;
  assign N1876 = N303;
  assign N1877 = N299;
  assign N1878 = N296;
  assign N1879 = N293;
  assign N1880 = N289;
  assign N1881 = N286;
  assign N1882 = N283;
  assign N1883 = N280;
  assign N1884 = N277;
  assign N1913 = N18;
  assign N1931 = N334;
  assign N1932 = N331;
  assign N1933 = N328;
  assign N1934 = N325;
  assign N1935 = N322;
  assign N1936 = N319;
  assign N1937 = N316;
  assign N1938 = N313;
  assign N1939 = N334;
  assign N1940 = N331;
  assign N1941 = N328;
  assign N1942 = N322;
  assign N1943 = N319;
  assign N1944 = N316;
  assign N1945 = N313;
  assign N1946 = N325;
  assign N1968 = N364;
  assign N1969 = N361;
  assign N1970 = N358;
  assign N1971 = N355;
  assign N1972 = N352;
  assign N1973 = N349;
  assign N1974 = N346;
  assign N1975 = N343;
  assign N1976 = N340;
  assign N1997 = N18;
  assign N2015 = N364;
  assign N2016 = N361;
  assign N2017 = N358;
  assign N2018 = N352;
  assign N2019 = N349;
  assign N2020 = N346;
  assign N2021 = N343;
  assign N2022 = N355;
  assign N2023 = N340;
  assign N2267 = N106;
  assign N2275 = N106;
  assign N2287 = N18;
  assign N2293 = N18;
  assign N2309 = N18;
  assign N2315 = N18;
  assign N2331 = N18;
  assign N2368 = N18;
  assign N2384 = N18;
  assign N2390 = N18;
  assign N2406 = N18;
  assign N2412 = N18;
  assign N241_O = N241_I;
  assign N387 = N1;
  assign N388 = N1;
  assign N478 = N248;
  assign N482 = N254;
  assign N484 = N257;
  assign N486 = N260;
  assign N489 = N263;
  assign N492 = N267;
  assign N501 = N274;
  assign N505 = N280;
  assign N507 = N283;
  assign N509 = N286;
  assign N511 = N289;
  assign N513 = N293;
  assign N515 = N296;
  assign N517 = N299;
  assign N519 = N303;
  assign N535 = N307;
  assign N537 = N310;
  assign N539 = N313;
  assign N541 = N316;
  assign N543 = N319;
  assign N545 = N322;
  assign N547 = N325;
  assign N549 = N328;
  assign N551 = N331;
  assign N553 = N334;
  assign N556 = N337;
  assign N559 = N343;
  assign N561 = N346;
  assign N563 = N349;
  assign N565 = N352;
  assign N567 = N355;
  assign N569 = N358;
  assign N571 = N361;
  assign N573 = N364;
  assign N582 = N1111;
  assign N590 = N1;
  assign N614 = N38;
  assign N625 = N15;
  assign N636 = N38;
  assign N643 = N251;
  assign N657 = N106;
  assign N676 = N18;
  assign N682 = N18;
  assign N689 = N18;
  assign N707 = N277;
  assign N750 = N367;
  assign N813 = N340;
  assign N871 = N367;
  assign N889 = N1;
  assign N945 = N106;
endmodule
