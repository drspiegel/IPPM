
module s838(GND, VDD, CK, C_0, C_1, C_10, C_11, C_12, C_13, C_14, C_15, C_16, C_17, C_18, C_19, C_2, C_20, C_21, C_22, C_23, C_24, C_25, C_26, C_27, C_28, C_29, C_3, C_30, C_31, C_32, C_4, C_5, C_6, C_7, C_8, C_9, P_0, Z);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  input CK;
  input C_0;
  input C_1;
  input C_10;
  input C_11;
  input C_12;
  input C_13;
  input C_14;
  input C_15;
  input C_16;
  input C_17;
  input C_18;
  input C_19;
  input C_2;
  input C_20;
  input C_21;
  input C_22;
  input C_23;
  input C_24;
  input C_25;
  input C_26;
  input C_27;
  input C_28;
  input C_29;
  input C_3;
  input C_30;
  input C_31;
  input C_32;
  input C_4;
  input C_5;
  input C_6;
  input C_7;
  input C_8;
  input C_9;
  wire \DFF_0.CK ;
  wire \DFF_0.D ;
  wire \DFF_0.Q ;
  wire \DFF_1.CK ;
  wire \DFF_1.D ;
  wire \DFF_1.Q ;
  wire \DFF_10.CK ;
  wire \DFF_10.D ;
  wire \DFF_10.Q ;
  wire \DFF_11.CK ;
  wire \DFF_11.D ;
  wire \DFF_11.Q ;
  wire \DFF_12.CK ;
  wire \DFF_12.D ;
  wire \DFF_12.Q ;
  wire \DFF_13.CK ;
  wire \DFF_13.D ;
  wire \DFF_13.Q ;
  wire \DFF_14.CK ;
  wire \DFF_14.D ;
  wire \DFF_14.Q ;
  wire \DFF_15.CK ;
  wire \DFF_15.D ;
  wire \DFF_15.Q ;
  wire \DFF_16.CK ;
  wire \DFF_16.D ;
  wire \DFF_16.Q ;
  wire \DFF_17.CK ;
  wire \DFF_17.D ;
  wire \DFF_17.Q ;
  wire \DFF_18.CK ;
  wire \DFF_18.D ;
  wire \DFF_18.Q ;
  wire \DFF_19.CK ;
  wire \DFF_19.D ;
  wire \DFF_19.Q ;
  wire \DFF_2.CK ;
  wire \DFF_2.D ;
  wire \DFF_2.Q ;
  wire \DFF_20.CK ;
  wire \DFF_20.D ;
  wire \DFF_20.Q ;
  wire \DFF_21.CK ;
  wire \DFF_21.D ;
  wire \DFF_21.Q ;
  wire \DFF_22.CK ;
  wire \DFF_22.D ;
  wire \DFF_22.Q ;
  wire \DFF_23.CK ;
  wire \DFF_23.D ;
  wire \DFF_23.Q ;
  wire \DFF_24.CK ;
  wire \DFF_24.D ;
  wire \DFF_24.Q ;
  wire \DFF_25.CK ;
  wire \DFF_25.D ;
  wire \DFF_25.Q ;
  wire \DFF_26.CK ;
  wire \DFF_26.D ;
  wire \DFF_26.Q ;
  wire \DFF_27.CK ;
  wire \DFF_27.D ;
  wire \DFF_27.Q ;
  wire \DFF_28.CK ;
  wire \DFF_28.D ;
  wire \DFF_28.Q ;
  wire \DFF_29.CK ;
  wire \DFF_29.D ;
  wire \DFF_29.Q ;
  wire \DFF_3.CK ;
  wire \DFF_3.D ;
  wire \DFF_3.Q ;
  wire \DFF_30.CK ;
  wire \DFF_30.D ;
  wire \DFF_30.Q ;
  wire \DFF_31.CK ;
  wire \DFF_31.D ;
  wire \DFF_31.Q ;
  wire \DFF_4.CK ;
  wire \DFF_4.D ;
  wire \DFF_4.Q ;
  wire \DFF_5.CK ;
  wire \DFF_5.D ;
  wire \DFF_5.Q ;
  wire \DFF_6.CK ;
  wire \DFF_6.D ;
  wire \DFF_6.Q ;
  wire \DFF_7.CK ;
  wire \DFF_7.D ;
  wire \DFF_7.Q ;
  wire \DFF_8.CK ;
  wire \DFF_8.D ;
  wire \DFF_8.Q ;
  wire \DFF_9.CK ;
  wire \DFF_9.D ;
  wire \DFF_9.Q ;
  input GND;
  wire I110;
  wire I111;
  wire I112;
  wire I113;
  wire I12;
  wire I13;
  wire I14;
  wire I15;
  wire I208;
  wire I209;
  wire I210;
  wire I211;
  wire I306;
  wire I307;
  wire I308;
  wire I309;
  wire I404;
  wire I405;
  wire I406;
  wire I407;
  wire I502;
  wire I503;
  wire I504;
  wire I505;
  wire I600;
  wire I601;
  wire I602;
  wire I603;
  wire I698;
  wire I699;
  wire I700;
  wire I701;
  input P_0;
  input VDD;
  wire X_1;
  wire X_10;
  wire X_11;
  wire X_12;
  wire X_13;
  wire X_14;
  wire X_15;
  wire X_16;
  wire X_17;
  wire X_18;
  wire X_19;
  wire X_2;
  wire X_20;
  wire X_21;
  wire X_22;
  wire X_23;
  wire X_24;
  wire X_25;
  wire X_26;
  wire X_27;
  wire X_28;
  wire X_29;
  wire X_3;
  wire X_30;
  wire X_31;
  wire X_32;
  wire X_4;
  wire X_5;
  wire X_6;
  wire X_7;
  wire X_8;
  wire X_9;
  output Z;
  al_aoi21 _137_ (
    .a(\DFF_3.Q ),
    .b(P_0),
    .c(\DFF_2.Q ),
    .y(_000_)
  );
  al_and3 _138_ (
    .a(\DFF_3.Q ),
    .b(\DFF_2.Q ),
    .c(P_0),
    .y(_001_)
  );
  al_nor2 _139_ (
    .a(_000_),
    .b(_001_),
    .y(\DFF_2.D )
  );
  al_and3 _140_ (
    .a(\DFF_1.Q ),
    .b(\DFF_0.Q ),
    .c(_001_),
    .y(_002_)
  );
  al_ao21 _141_ (
    .a(\DFF_7.Q ),
    .b(_002_),
    .c(\DFF_6.Q ),
    .y(_003_)
  );
  al_and3 _142_ (
    .a(\DFF_7.Q ),
    .b(\DFF_6.Q ),
    .c(_002_),
    .y(_004_)
  );
  al_and2ft _143_ (
    .a(_004_),
    .b(_003_),
    .y(\DFF_6.D )
  );
  al_and3 _144_ (
    .a(\DFF_5.Q ),
    .b(\DFF_4.Q ),
    .c(_004_),
    .y(_005_)
  );
  al_ao21 _145_ (
    .a(\DFF_11.Q ),
    .b(_005_),
    .c(\DFF_10.Q ),
    .y(_006_)
  );
  al_and3 _146_ (
    .a(\DFF_11.Q ),
    .b(\DFF_10.Q ),
    .c(_005_),
    .y(_007_)
  );
  al_and2ft _147_ (
    .a(_007_),
    .b(_006_),
    .y(\DFF_10.D )
  );
  al_and3 _148_ (
    .a(\DFF_9.Q ),
    .b(\DFF_8.Q ),
    .c(_007_),
    .y(_008_)
  );
  al_ao21 _149_ (
    .a(\DFF_15.Q ),
    .b(_008_),
    .c(\DFF_14.Q ),
    .y(_009_)
  );
  al_and3 _150_ (
    .a(\DFF_15.Q ),
    .b(\DFF_14.Q ),
    .c(_008_),
    .y(_010_)
  );
  al_and2ft _151_ (
    .a(_010_),
    .b(_009_),
    .y(\DFF_14.D )
  );
  al_and3 _152_ (
    .a(\DFF_13.Q ),
    .b(\DFF_12.Q ),
    .c(_010_),
    .y(_011_)
  );
  al_ao21 _153_ (
    .a(\DFF_19.Q ),
    .b(_011_),
    .c(\DFF_18.Q ),
    .y(_012_)
  );
  al_and3 _154_ (
    .a(\DFF_19.Q ),
    .b(\DFF_18.Q ),
    .c(_011_),
    .y(_013_)
  );
  al_and2ft _155_ (
    .a(_013_),
    .b(_012_),
    .y(\DFF_18.D )
  );
  al_and3 _156_ (
    .a(\DFF_17.Q ),
    .b(\DFF_16.Q ),
    .c(_013_),
    .y(_014_)
  );
  al_ao21 _157_ (
    .a(\DFF_23.Q ),
    .b(_014_),
    .c(\DFF_22.Q ),
    .y(_015_)
  );
  al_and3 _158_ (
    .a(\DFF_23.Q ),
    .b(\DFF_22.Q ),
    .c(_014_),
    .y(_016_)
  );
  al_and2ft _159_ (
    .a(_016_),
    .b(_015_),
    .y(\DFF_22.D )
  );
  al_and3 _160_ (
    .a(\DFF_21.Q ),
    .b(\DFF_20.Q ),
    .c(_016_),
    .y(_017_)
  );
  al_ao21 _161_ (
    .a(\DFF_27.Q ),
    .b(_017_),
    .c(\DFF_26.Q ),
    .y(_018_)
  );
  al_and3 _162_ (
    .a(\DFF_27.Q ),
    .b(\DFF_26.Q ),
    .c(_017_),
    .y(_019_)
  );
  al_and2ft _163_ (
    .a(_019_),
    .b(_018_),
    .y(\DFF_26.D )
  );
  al_and3 _164_ (
    .a(\DFF_25.Q ),
    .b(\DFF_24.Q ),
    .c(_019_),
    .y(_020_)
  );
  al_ao21 _165_ (
    .a(\DFF_31.Q ),
    .b(_020_),
    .c(\DFF_30.Q ),
    .y(_021_)
  );
  al_and3 _166_ (
    .a(\DFF_31.Q ),
    .b(\DFF_30.Q ),
    .c(_020_),
    .y(_022_)
  );
  al_and2ft _167_ (
    .a(_022_),
    .b(_021_),
    .y(\DFF_30.D )
  );
  al_ao21 _168_ (
    .a(\DFF_1.Q ),
    .b(_001_),
    .c(\DFF_0.Q ),
    .y(_023_)
  );
  al_and2ft _169_ (
    .a(_002_),
    .b(_023_),
    .y(\DFF_0.D )
  );
  al_ao21 _170_ (
    .a(\DFF_5.Q ),
    .b(_004_),
    .c(\DFF_4.Q ),
    .y(_024_)
  );
  al_and2ft _171_ (
    .a(_005_),
    .b(_024_),
    .y(\DFF_4.D )
  );
  al_ao21 _172_ (
    .a(\DFF_9.Q ),
    .b(_007_),
    .c(\DFF_8.Q ),
    .y(_025_)
  );
  al_and2ft _173_ (
    .a(_008_),
    .b(_025_),
    .y(\DFF_8.D )
  );
  al_ao21 _174_ (
    .a(\DFF_13.Q ),
    .b(_010_),
    .c(\DFF_12.Q ),
    .y(_026_)
  );
  al_and2ft _175_ (
    .a(_011_),
    .b(_026_),
    .y(\DFF_12.D )
  );
  al_ao21 _176_ (
    .a(\DFF_17.Q ),
    .b(_013_),
    .c(\DFF_16.Q ),
    .y(_027_)
  );
  al_and2ft _177_ (
    .a(_014_),
    .b(_027_),
    .y(\DFF_16.D )
  );
  al_ao21 _178_ (
    .a(\DFF_21.Q ),
    .b(_016_),
    .c(\DFF_20.Q ),
    .y(_028_)
  );
  al_and2ft _179_ (
    .a(_017_),
    .b(_028_),
    .y(\DFF_20.D )
  );
  al_ao21 _180_ (
    .a(\DFF_25.Q ),
    .b(_019_),
    .c(\DFF_24.Q ),
    .y(_029_)
  );
  al_and2ft _181_ (
    .a(_020_),
    .b(_029_),
    .y(\DFF_24.D )
  );
  al_inv _182_ (
    .a(\DFF_28.Q ),
    .y(_030_)
  );
  al_ao21 _183_ (
    .a(\DFF_29.Q ),
    .b(_022_),
    .c(_030_),
    .y(_031_)
  );
  al_and3 _184_ (
    .a(\DFF_29.Q ),
    .b(_030_),
    .c(_022_),
    .y(_032_)
  );
  al_nand2ft _185_ (
    .a(_032_),
    .b(_031_),
    .y(\DFF_28.D )
  );
  al_and2 _186_ (
    .a(\DFF_31.Q ),
    .b(_020_),
    .y(_033_)
  );
  al_nand3 _187_ (
    .a(\DFF_30.Q ),
    .b(\DFF_29.Q ),
    .c(_033_),
    .y(_034_)
  );
  al_nand3 _188_ (
    .a(\DFF_31.Q ),
    .b(\DFF_30.Q ),
    .c(_020_),
    .y(_035_)
  );
  al_and2ft _189_ (
    .a(\DFF_29.Q ),
    .b(_035_),
    .y(_036_)
  );
  al_and2ft _190_ (
    .a(_036_),
    .b(_034_),
    .y(\DFF_29.D )
  );
  al_and2 _191_ (
    .a(\DFF_1.Q ),
    .b(_001_),
    .y(_037_)
  );
  al_or2 _192_ (
    .a(\DFF_1.Q ),
    .b(_001_),
    .y(_038_)
  );
  al_and2ft _193_ (
    .a(_037_),
    .b(_038_),
    .y(\DFF_1.D )
  );
  al_and2ft _194_ (
    .a(P_0),
    .b(\DFF_3.Q ),
    .y(_039_)
  );
  al_nand2ft _195_ (
    .a(\DFF_3.Q ),
    .b(P_0),
    .y(_040_)
  );
  al_nand2ft _196_ (
    .a(_039_),
    .b(_040_),
    .y(\DFF_3.D )
  );
  al_and2 _197_ (
    .a(\DFF_5.Q ),
    .b(_004_),
    .y(_041_)
  );
  al_or2 _198_ (
    .a(\DFF_5.Q ),
    .b(_004_),
    .y(_042_)
  );
  al_and2ft _199_ (
    .a(_041_),
    .b(_042_),
    .y(\DFF_5.D )
  );
  al_and2 _200_ (
    .a(\DFF_7.Q ),
    .b(_002_),
    .y(_043_)
  );
  al_or2 _201_ (
    .a(\DFF_7.Q ),
    .b(_002_),
    .y(_044_)
  );
  al_and2ft _202_ (
    .a(_043_),
    .b(_044_),
    .y(\DFF_7.D )
  );
  al_and2 _203_ (
    .a(\DFF_9.Q ),
    .b(_007_),
    .y(_045_)
  );
  al_or2 _204_ (
    .a(\DFF_9.Q ),
    .b(_007_),
    .y(_046_)
  );
  al_and2ft _205_ (
    .a(_045_),
    .b(_046_),
    .y(\DFF_9.D )
  );
  al_and2 _206_ (
    .a(\DFF_11.Q ),
    .b(_005_),
    .y(_047_)
  );
  al_or2 _207_ (
    .a(\DFF_11.Q ),
    .b(_005_),
    .y(_048_)
  );
  al_and2ft _208_ (
    .a(_047_),
    .b(_048_),
    .y(\DFF_11.D )
  );
  al_and2 _209_ (
    .a(\DFF_13.Q ),
    .b(_010_),
    .y(_049_)
  );
  al_or2 _210_ (
    .a(\DFF_13.Q ),
    .b(_010_),
    .y(_050_)
  );
  al_and2ft _211_ (
    .a(_049_),
    .b(_050_),
    .y(\DFF_13.D )
  );
  al_and2 _212_ (
    .a(\DFF_15.Q ),
    .b(_008_),
    .y(_051_)
  );
  al_or2 _213_ (
    .a(\DFF_15.Q ),
    .b(_008_),
    .y(_052_)
  );
  al_and2ft _214_ (
    .a(_051_),
    .b(_052_),
    .y(\DFF_15.D )
  );
  al_and2 _215_ (
    .a(\DFF_17.Q ),
    .b(_013_),
    .y(_053_)
  );
  al_or2 _216_ (
    .a(\DFF_17.Q ),
    .b(_013_),
    .y(_054_)
  );
  al_and2ft _217_ (
    .a(_053_),
    .b(_054_),
    .y(\DFF_17.D )
  );
  al_and2 _218_ (
    .a(\DFF_19.Q ),
    .b(_011_),
    .y(_055_)
  );
  al_or2 _219_ (
    .a(\DFF_19.Q ),
    .b(_011_),
    .y(_056_)
  );
  al_and2ft _220_ (
    .a(_055_),
    .b(_056_),
    .y(\DFF_19.D )
  );
  al_and2 _221_ (
    .a(\DFF_21.Q ),
    .b(_016_),
    .y(_057_)
  );
  al_or2 _222_ (
    .a(\DFF_21.Q ),
    .b(_016_),
    .y(_058_)
  );
  al_and2ft _223_ (
    .a(_057_),
    .b(_058_),
    .y(\DFF_21.D )
  );
  al_and2 _224_ (
    .a(\DFF_23.Q ),
    .b(_014_),
    .y(_059_)
  );
  al_or2 _225_ (
    .a(\DFF_23.Q ),
    .b(_014_),
    .y(_060_)
  );
  al_and2ft _226_ (
    .a(_059_),
    .b(_060_),
    .y(\DFF_23.D )
  );
  al_and2 _227_ (
    .a(\DFF_25.Q ),
    .b(_019_),
    .y(_061_)
  );
  al_or2 _228_ (
    .a(\DFF_25.Q ),
    .b(_019_),
    .y(_062_)
  );
  al_and2ft _229_ (
    .a(_061_),
    .b(_062_),
    .y(\DFF_25.D )
  );
  al_and2 _230_ (
    .a(\DFF_27.Q ),
    .b(_017_),
    .y(_063_)
  );
  al_or2 _231_ (
    .a(\DFF_27.Q ),
    .b(_017_),
    .y(_064_)
  );
  al_and2ft _232_ (
    .a(_063_),
    .b(_064_),
    .y(\DFF_27.D )
  );
  al_or2 _233_ (
    .a(\DFF_31.Q ),
    .b(_020_),
    .y(_065_)
  );
  al_and2ft _234_ (
    .a(_033_),
    .b(_065_),
    .y(\DFF_31.D )
  );
  al_or3 _235_ (
    .a(\DFF_2.Q ),
    .b(\DFF_1.Q ),
    .c(\DFF_0.Q ),
    .y(_066_)
  );
  al_nor2 _236_ (
    .a(\DFF_3.Q ),
    .b(\DFF_7.Q ),
    .y(_067_)
  );
  al_or3 _237_ (
    .a(\DFF_6.Q ),
    .b(\DFF_5.Q ),
    .c(\DFF_4.Q ),
    .y(_068_)
  );
  al_and3fft _238_ (
    .a(_066_),
    .b(_068_),
    .c(_067_),
    .y(_069_)
  );
  al_and2ft _239_ (
    .a(\DFF_10.Q ),
    .b(_069_),
    .y(_070_)
  );
  al_nor2 _240_ (
    .a(\DFF_15.Q ),
    .b(\DFF_14.Q ),
    .y(_071_)
  );
  al_nor2 _241_ (
    .a(\DFF_11.Q ),
    .b(\DFF_9.Q ),
    .y(_072_)
  );
  al_or2 _242_ (
    .a(\DFF_8.Q ),
    .b(\DFF_13.Q ),
    .y(_073_)
  );
  al_and3ftt _243_ (
    .a(_073_),
    .b(_071_),
    .c(_072_),
    .y(_074_)
  );
  al_or2 _244_ (
    .a(\DFF_19.Q ),
    .b(\DFF_18.Q ),
    .y(_075_)
  );
  al_nor2 _245_ (
    .a(\DFF_12.Q ),
    .b(\DFF_17.Q ),
    .y(_076_)
  );
  al_and3fft _246_ (
    .a(\DFF_16.Q ),
    .b(_075_),
    .c(_076_),
    .y(_077_)
  );
  al_and3 _247_ (
    .a(_074_),
    .b(_077_),
    .c(_070_),
    .y(_078_)
  );
  al_nor2 _248_ (
    .a(\DFF_23.Q ),
    .b(\DFF_22.Q ),
    .y(_079_)
  );
  al_nand3fft _249_ (
    .a(\DFF_21.Q ),
    .b(\DFF_20.Q ),
    .c(_079_),
    .y(_080_)
  );
  al_aoi21 _250_ (
    .a(\DFF_28.Q ),
    .b(C_32),
    .c(\DFF_29.Q ),
    .y(_081_)
  );
  al_nand2ft _251_ (
    .a(C_31),
    .b(\DFF_29.Q ),
    .y(_082_)
  );
  al_and3fft _252_ (
    .a(\DFF_30.Q ),
    .b(_081_),
    .c(_082_),
    .y(_083_)
  );
  al_and2 _253_ (
    .a(\DFF_30.Q ),
    .b(C_30),
    .y(_084_)
  );
  al_mux2l _254_ (
    .a(_084_),
    .b(_083_),
    .s(\DFF_31.Q ),
    .y(_085_)
  );
  al_ao21 _255_ (
    .a(\DFF_31.Q ),
    .b(C_29),
    .c(\DFF_24.Q ),
    .y(_086_)
  );
  al_or3 _256_ (
    .a(\DFF_27.Q ),
    .b(\DFF_26.Q ),
    .c(\DFF_25.Q ),
    .y(_087_)
  );
  al_ao21ftt _257_ (
    .a(C_28),
    .b(\DFF_24.Q ),
    .c(_087_),
    .y(_088_)
  );
  al_mux2l _258_ (
    .a(_086_),
    .b(_085_),
    .s(_088_),
    .y(_089_)
  );
  al_nand3ftt _259_ (
    .a(\DFF_27.Q ),
    .b(\DFF_26.Q ),
    .c(C_26),
    .y(_090_)
  );
  al_ao21ttf _260_ (
    .a(\DFF_27.Q ),
    .b(C_25),
    .c(_090_),
    .y(_091_)
  );
  al_or2 _261_ (
    .a(_091_),
    .b(_089_),
    .y(_092_)
  );
  al_nand3ftt _262_ (
    .a(_080_),
    .b(_078_),
    .c(_092_),
    .y(_093_)
  );
  al_nand3ftt _263_ (
    .a(\DFF_23.Q ),
    .b(\DFF_22.Q ),
    .c(C_22),
    .y(_094_)
  );
  al_ao21ttf _264_ (
    .a(\DFF_23.Q ),
    .b(C_21),
    .c(_094_),
    .y(_095_)
  );
  al_ao21 _265_ (
    .a(\DFF_20.Q ),
    .b(C_24),
    .c(\DFF_21.Q ),
    .y(_096_)
  );
  al_aoi21ftf _266_ (
    .a(C_23),
    .b(\DFF_21.Q ),
    .c(_079_),
    .y(_097_)
  );
  al_ao21 _267_ (
    .a(_096_),
    .b(_097_),
    .c(_095_),
    .y(_098_)
  );
  al_aoi21 _268_ (
    .a(_098_),
    .b(_078_),
    .c(C_0),
    .y(_099_)
  );
  al_aoi21 _269_ (
    .a(\DFF_16.Q ),
    .b(C_20),
    .c(\DFF_17.Q ),
    .y(_100_)
  );
  al_nand2ft _270_ (
    .a(C_19),
    .b(\DFF_17.Q ),
    .y(_101_)
  );
  al_nand3fft _271_ (
    .a(_075_),
    .b(_100_),
    .c(_101_),
    .y(_102_)
  );
  al_ao21 _272_ (
    .a(\DFF_18.Q ),
    .b(C_18),
    .c(\DFF_19.Q ),
    .y(_103_)
  );
  al_ao21ftf _273_ (
    .a(C_17),
    .b(\DFF_19.Q ),
    .c(_103_),
    .y(_104_)
  );
  al_and3ftt _274_ (
    .a(\DFF_12.Q ),
    .b(_104_),
    .c(_102_),
    .y(_105_)
  );
  al_aoi21ftf _275_ (
    .a(C_16),
    .b(\DFF_12.Q ),
    .c(_074_),
    .y(_106_)
  );
  al_nand3ftt _276_ (
    .a(_105_),
    .b(_070_),
    .c(_106_),
    .y(_107_)
  );
  al_nand3 _277_ (
    .a(_099_),
    .b(_107_),
    .c(_093_),
    .y(_108_)
  );
  al_nand3 _278_ (
    .a(\DFF_13.Q ),
    .b(C_15),
    .c(_071_),
    .y(_109_)
  );
  al_nand3ftt _279_ (
    .a(\DFF_15.Q ),
    .b(\DFF_14.Q ),
    .c(C_14),
    .y(_110_)
  );
  al_aoi21 _280_ (
    .a(\DFF_15.Q ),
    .b(C_13),
    .c(\DFF_8.Q ),
    .y(_111_)
  );
  al_and3 _281_ (
    .a(_110_),
    .b(_111_),
    .c(_109_),
    .y(_112_)
  );
  al_ao21 _282_ (
    .a(\DFF_9.Q ),
    .b(C_11),
    .c(\DFF_10.Q ),
    .y(_113_)
  );
  al_oai21ftf _283_ (
    .a(\DFF_8.Q ),
    .b(C_12),
    .c(\DFF_9.Q ),
    .y(_114_)
  );
  al_mux2l _284_ (
    .a(_114_),
    .b(_112_),
    .s(_113_),
    .y(_115_)
  );
  al_and2ft _285_ (
    .a(C_10),
    .b(\DFF_10.Q ),
    .y(_116_)
  );
  al_mux2l _286_ (
    .a(_116_),
    .b(_115_),
    .s(\DFF_11.Q ),
    .y(_117_)
  );
  al_and2ft _287_ (
    .a(C_9),
    .b(\DFF_11.Q ),
    .y(_118_)
  );
  al_and3fft _288_ (
    .a(_118_),
    .b(_117_),
    .c(_069_),
    .y(_119_)
  );
  al_mux2h _289_ (
    .a(_119_),
    .b(_108_),
    .s(P_0),
    .y(_120_)
  );
  al_and3fft _290_ (
    .a(\DFF_27.Q ),
    .b(\DFF_26.Q ),
    .c(P_0),
    .y(_121_)
  );
  al_and3 _291_ (
    .a(\DFF_25.Q ),
    .b(C_27),
    .c(_121_),
    .y(_122_)
  );
  al_nand3ftt _292_ (
    .a(_080_),
    .b(_122_),
    .c(_078_),
    .y(_123_)
  );
  al_nand3 _293_ (
    .a(\DFF_3.Q ),
    .b(P_0),
    .c(C_1),
    .y(_124_)
  );
  al_ao21 _294_ (
    .a(\DFF_0.Q ),
    .b(C_4),
    .c(\DFF_1.Q ),
    .y(_125_)
  );
  al_ao21ftf _295_ (
    .a(C_3),
    .b(\DFF_1.Q ),
    .c(_125_),
    .y(_126_)
  );
  al_aoi21ftt _296_ (
    .a(C_2),
    .b(\DFF_2.Q ),
    .c(_040_),
    .y(_127_)
  );
  al_ao21ftf _297_ (
    .a(\DFF_2.Q ),
    .b(_126_),
    .c(_127_),
    .y(_128_)
  );
  al_ao21 _298_ (
    .a(\DFF_4.Q ),
    .b(C_8),
    .c(\DFF_5.Q ),
    .y(_129_)
  );
  al_nand2ft _299_ (
    .a(C_7),
    .b(\DFF_5.Q ),
    .y(_130_)
  );
  al_nand3ftt _300_ (
    .a(\DFF_6.Q ),
    .b(_130_),
    .c(_129_),
    .y(_131_)
  );
  al_ao21 _301_ (
    .a(\DFF_6.Q ),
    .b(C_6),
    .c(\DFF_7.Q ),
    .y(_132_)
  );
  al_nand2ft _302_ (
    .a(C_5),
    .b(\DFF_7.Q ),
    .y(_133_)
  );
  al_and3fft _303_ (
    .a(_040_),
    .b(_066_),
    .c(_133_),
    .y(_134_)
  );
  al_ao21ftf _304_ (
    .a(_132_),
    .b(_131_),
    .c(_134_),
    .y(_135_)
  );
  al_and3 _305_ (
    .a(_124_),
    .b(_128_),
    .c(_135_),
    .y(_136_)
  );
  al_or3fft _306_ (
    .a(_123_),
    .b(_136_),
    .c(_120_),
    .y(Z)
  );
  al_dffl _307_ (
    .clk(CK),
    .d(\DFF_0.D ),
    .q(\DFF_0.Q )
  );
  al_dffl _308_ (
    .clk(CK),
    .d(\DFF_1.D ),
    .q(\DFF_1.Q )
  );
  al_dffl _309_ (
    .clk(CK),
    .d(\DFF_2.D ),
    .q(\DFF_2.Q )
  );
  al_dffl _310_ (
    .clk(CK),
    .d(\DFF_3.D ),
    .q(\DFF_3.Q )
  );
  al_dffl _311_ (
    .clk(CK),
    .d(\DFF_4.D ),
    .q(\DFF_4.Q )
  );
  al_dffl _312_ (
    .clk(CK),
    .d(\DFF_5.D ),
    .q(\DFF_5.Q )
  );
  al_dffl _313_ (
    .clk(CK),
    .d(\DFF_6.D ),
    .q(\DFF_6.Q )
  );
  al_dffl _314_ (
    .clk(CK),
    .d(\DFF_7.D ),
    .q(\DFF_7.Q )
  );
  al_dffl _315_ (
    .clk(CK),
    .d(\DFF_8.D ),
    .q(\DFF_8.Q )
  );
  al_dffl _316_ (
    .clk(CK),
    .d(\DFF_9.D ),
    .q(\DFF_9.Q )
  );
  al_dffl _317_ (
    .clk(CK),
    .d(\DFF_10.D ),
    .q(\DFF_10.Q )
  );
  al_dffl _318_ (
    .clk(CK),
    .d(\DFF_11.D ),
    .q(\DFF_11.Q )
  );
  al_dffl _319_ (
    .clk(CK),
    .d(\DFF_12.D ),
    .q(\DFF_12.Q )
  );
  al_dffl _320_ (
    .clk(CK),
    .d(\DFF_13.D ),
    .q(\DFF_13.Q )
  );
  al_dffl _321_ (
    .clk(CK),
    .d(\DFF_14.D ),
    .q(\DFF_14.Q )
  );
  al_dffl _322_ (
    .clk(CK),
    .d(\DFF_15.D ),
    .q(\DFF_15.Q )
  );
  al_dffl _323_ (
    .clk(CK),
    .d(\DFF_16.D ),
    .q(\DFF_16.Q )
  );
  al_dffl _324_ (
    .clk(CK),
    .d(\DFF_17.D ),
    .q(\DFF_17.Q )
  );
  al_dffl _325_ (
    .clk(CK),
    .d(\DFF_18.D ),
    .q(\DFF_18.Q )
  );
  al_dffl _326_ (
    .clk(CK),
    .d(\DFF_19.D ),
    .q(\DFF_19.Q )
  );
  al_dffl _327_ (
    .clk(CK),
    .d(\DFF_20.D ),
    .q(\DFF_20.Q )
  );
  al_dffl _328_ (
    .clk(CK),
    .d(\DFF_21.D ),
    .q(\DFF_21.Q )
  );
  al_dffl _329_ (
    .clk(CK),
    .d(\DFF_22.D ),
    .q(\DFF_22.Q )
  );
  al_dffl _330_ (
    .clk(CK),
    .d(\DFF_23.D ),
    .q(\DFF_23.Q )
  );
  al_dffl _331_ (
    .clk(CK),
    .d(\DFF_24.D ),
    .q(\DFF_24.Q )
  );
  al_dffl _332_ (
    .clk(CK),
    .d(\DFF_25.D ),
    .q(\DFF_25.Q )
  );
  al_dffl _333_ (
    .clk(CK),
    .d(\DFF_26.D ),
    .q(\DFF_26.Q )
  );
  al_dffl _334_ (
    .clk(CK),
    .d(\DFF_27.D ),
    .q(\DFF_27.Q )
  );
  al_dffl _335_ (
    .clk(CK),
    .d(\DFF_28.D ),
    .q(\DFF_28.Q )
  );
  al_dffl _336_ (
    .clk(CK),
    .d(\DFF_29.D ),
    .q(\DFF_29.Q )
  );
  al_dffl _337_ (
    .clk(CK),
    .d(\DFF_30.D ),
    .q(\DFF_30.Q )
  );
  al_dffl _338_ (
    .clk(CK),
    .d(\DFF_31.D ),
    .q(\DFF_31.Q )
  );
  assign \DFF_0.CK  = CK;
  assign \DFF_1.CK  = CK;
  assign \DFF_10.CK  = CK;
  assign \DFF_11.CK  = CK;
  assign \DFF_12.CK  = CK;
  assign \DFF_13.CK  = CK;
  assign \DFF_14.CK  = CK;
  assign \DFF_15.CK  = CK;
  assign \DFF_16.CK  = CK;
  assign \DFF_17.CK  = CK;
  assign \DFF_18.CK  = CK;
  assign \DFF_19.CK  = CK;
  assign \DFF_2.CK  = CK;
  assign \DFF_20.CK  = CK;
  assign \DFF_21.CK  = CK;
  assign \DFF_22.CK  = CK;
  assign \DFF_23.CK  = CK;
  assign \DFF_24.CK  = CK;
  assign \DFF_25.CK  = CK;
  assign \DFF_26.CK  = CK;
  assign \DFF_27.CK  = CK;
  assign \DFF_28.CK  = CK;
  assign \DFF_29.CK  = CK;
  assign \DFF_3.CK  = CK;
  assign \DFF_30.CK  = CK;
  assign \DFF_31.CK  = CK;
  assign \DFF_4.CK  = CK;
  assign \DFF_5.CK  = CK;
  assign \DFF_6.CK  = CK;
  assign \DFF_7.CK  = CK;
  assign \DFF_8.CK  = CK;
  assign \DFF_9.CK  = CK;
  assign I110 = \DFF_4.D ;
  assign I111 = \DFF_5.D ;
  assign I112 = \DFF_6.D ;
  assign I113 = \DFF_7.D ;
  assign I12 = \DFF_0.D ;
  assign I13 = \DFF_1.D ;
  assign I14 = \DFF_2.D ;
  assign I15 = \DFF_3.D ;
  assign I208 = \DFF_8.D ;
  assign I209 = \DFF_9.D ;
  assign I210 = \DFF_10.D ;
  assign I211 = \DFF_11.D ;
  assign I306 = \DFF_12.D ;
  assign I307 = \DFF_13.D ;
  assign I308 = \DFF_14.D ;
  assign I309 = \DFF_15.D ;
  assign I404 = \DFF_16.D ;
  assign I405 = \DFF_17.D ;
  assign I406 = \DFF_18.D ;
  assign I407 = \DFF_19.D ;
  assign I502 = \DFF_20.D ;
  assign I503 = \DFF_21.D ;
  assign I504 = \DFF_22.D ;
  assign I505 = \DFF_23.D ;
  assign I600 = \DFF_24.D ;
  assign I601 = \DFF_25.D ;
  assign I602 = \DFF_26.D ;
  assign I603 = \DFF_27.D ;
  assign I698 = \DFF_28.D ;
  assign I699 = \DFF_29.D ;
  assign I700 = \DFF_30.D ;
  assign I701 = \DFF_31.D ;
  assign X_1 = \DFF_3.Q ;
  assign X_10 = \DFF_10.Q ;
  assign X_11 = \DFF_9.Q ;
  assign X_12 = \DFF_8.Q ;
  assign X_13 = \DFF_15.Q ;
  assign X_14 = \DFF_14.Q ;
  assign X_15 = \DFF_13.Q ;
  assign X_16 = \DFF_12.Q ;
  assign X_17 = \DFF_19.Q ;
  assign X_18 = \DFF_18.Q ;
  assign X_19 = \DFF_17.Q ;
  assign X_2 = \DFF_2.Q ;
  assign X_20 = \DFF_16.Q ;
  assign X_21 = \DFF_23.Q ;
  assign X_22 = \DFF_22.Q ;
  assign X_23 = \DFF_21.Q ;
  assign X_24 = \DFF_20.Q ;
  assign X_25 = \DFF_27.Q ;
  assign X_26 = \DFF_26.Q ;
  assign X_27 = \DFF_25.Q ;
  assign X_28 = \DFF_24.Q ;
  assign X_29 = \DFF_31.Q ;
  assign X_3 = \DFF_1.Q ;
  assign X_30 = \DFF_30.Q ;
  assign X_31 = \DFF_29.Q ;
  assign X_32 = \DFF_28.Q ;
  assign X_4 = \DFF_0.Q ;
  assign X_5 = \DFF_7.Q ;
  assign X_6 = \DFF_6.Q ;
  assign X_7 = \DFF_5.Q ;
  assign X_8 = \DFF_4.Q ;
  assign X_9 = \DFF_11.Q ;
endmodule
