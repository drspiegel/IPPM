
module s1488(GND, VDD, CK, CLR, v0, v1, v13_D_10, v13_D_11, v13_D_12, v13_D_13, v13_D_14, v13_D_15, v13_D_16, v13_D_17, v13_D_18, v13_D_19, v13_D_20, v13_D_21, v13_D_22, v13_D_23, v13_D_24, v13_D_6, v13_D_7, v13_D_8, v13_D_9, v2, v3, v4, v5, v6);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  wire _332_;
  wire _333_;
  wire _334_;
  wire _335_;
  wire _336_;
  wire _337_;
  wire _338_;
  wire _339_;
  wire _340_;
  wire _341_;
  wire Av13_D_10B;
  wire Av13_D_11B;
  wire Av13_D_12B;
  wire Av13_D_13B;
  wire Av13_D_14B;
  wire Av13_D_15B;
  wire Av13_D_16B;
  wire Av13_D_17B;
  wire Av13_D_18B;
  wire Av13_D_19B;
  wire Av13_D_20B;
  wire Av13_D_21B;
  wire Av13_D_22B;
  wire Av13_D_23B;
  wire Av13_D_24B;
  wire Av13_D_6B;
  wire Av13_D_7B;
  wire Av13_D_8B;
  wire Av13_D_9B;
  wire C193D;
  wire C79D;
  input CK;
  input CLR;
  wire \DFF_0.CK ;
  wire \DFF_0.D ;
  wire \DFF_0.Q ;
  wire \DFF_1.CK ;
  wire \DFF_1.D ;
  wire \DFF_1.Q ;
  wire \DFF_2.CK ;
  wire \DFF_2.D ;
  wire \DFF_2.Q ;
  wire \DFF_3.CK ;
  wire \DFF_3.D ;
  wire \DFF_3.Q ;
  wire \DFF_4.CK ;
  wire \DFF_4.D ;
  wire \DFF_4.Q ;
  wire \DFF_5.CK ;
  wire \DFF_5.D ;
  wire \DFF_5.Q ;
  input GND;
  wire II143;
  wire IIII518;
  input VDD;
  input v0;
  input v1;
  wire v10;
  wire v11;
  wire v12;
  wire v13_D_0C;
  output v13_D_10;
  output v13_D_11;
  output v13_D_12;
  output v13_D_13;
  output v13_D_14;
  output v13_D_15;
  output v13_D_16;
  output v13_D_17;
  output v13_D_18;
  output v13_D_19;
  wire v13_D_1C;
  output v13_D_20;
  output v13_D_21;
  output v13_D_22;
  output v13_D_23;
  output v13_D_24;
  wire v13_D_2C;
  wire v13_D_3C;
  wire v13_D_4C;
  wire v13_D_5C;
  output v13_D_6;
  output v13_D_7;
  output v13_D_8;
  output v13_D_9;
  input v2;
  input v3;
  input v4;
  input v5;
  input v6;
  wire v7;
  wire v8;
  wire v9;
  al_nand2ft _342_ (
    .a(v1),
    .b(v6),
    .y(_283_)
  );
  al_and3 _343_ (
    .a(\DFF_4.Q ),
    .b(\DFF_2.Q ),
    .c(_283_),
    .y(_290_)
  );
  al_and3 _344_ (
    .a(v3),
    .b(\DFF_0.Q ),
    .c(\DFF_3.Q ),
    .y(_291_)
  );
  al_nand2ft _345_ (
    .a(\DFF_5.Q ),
    .b(\DFF_1.Q ),
    .y(_292_)
  );
  al_and3ftt _346_ (
    .a(_292_),
    .b(_291_),
    .c(_290_),
    .y(v13_D_20)
  );
  al_inv _347_ (
    .a(\DFF_5.Q ),
    .y(_293_)
  );
  al_inv _348_ (
    .a(v2),
    .y(_294_)
  );
  al_and2 _349_ (
    .a(\DFF_4.Q ),
    .b(\DFF_3.Q ),
    .y(_295_)
  );
  al_nand2 _350_ (
    .a(v4),
    .b(v5),
    .y(_296_)
  );
  al_or2 _351_ (
    .a(\DFF_4.Q ),
    .b(\DFF_1.Q ),
    .y(_297_)
  );
  al_or3 _352_ (
    .a(\DFF_3.Q ),
    .b(_297_),
    .c(_296_),
    .y(_298_)
  );
  al_ao21ftf _353_ (
    .a(_294_),
    .b(_295_),
    .c(_298_),
    .y(_299_)
  );
  al_nor2 _354_ (
    .a(\DFF_0.Q ),
    .b(\DFF_2.Q ),
    .y(_300_)
  );
  al_and3 _355_ (
    .a(_293_),
    .b(_300_),
    .c(_299_),
    .y(v13_D_21)
  );
  al_nand3 _356_ (
    .a(\DFF_4.Q ),
    .b(v2),
    .c(\DFF_1.Q ),
    .y(_301_)
  );
  al_and2ft _357_ (
    .a(\DFF_3.Q ),
    .b(\DFF_0.Q ),
    .y(_302_)
  );
  al_and3 _358_ (
    .a(\DFF_5.Q ),
    .b(\DFF_2.Q ),
    .c(_302_),
    .y(_303_)
  );
  al_and3fft _359_ (
    .a(\DFF_5.Q ),
    .b(\DFF_1.Q ),
    .c(v3),
    .y(_304_)
  );
  al_nand3ftt _360_ (
    .a(\DFF_0.Q ),
    .b(v6),
    .c(\DFF_2.Q ),
    .y(_305_)
  );
  al_nand3ftt _361_ (
    .a(_305_),
    .b(_295_),
    .c(_304_),
    .y(_306_)
  );
  al_ao21ftf _362_ (
    .a(_301_),
    .b(_303_),
    .c(_306_),
    .y(v13_D_16)
  );
  al_nor2 _363_ (
    .a(\DFF_5.Q ),
    .b(\DFF_0.Q ),
    .y(_307_)
  );
  al_inv _364_ (
    .a(_307_),
    .y(_308_)
  );
  al_nor2 _365_ (
    .a(\DFF_3.Q ),
    .b(\DFF_2.Q ),
    .y(_309_)
  );
  al_nand3fft _366_ (
    .a(_297_),
    .b(_296_),
    .c(_309_),
    .y(_310_)
  );
  al_and2ft _367_ (
    .a(\DFF_3.Q ),
    .b(\DFF_2.Q ),
    .y(_311_)
  );
  al_nand3fft _368_ (
    .a(v0),
    .b(\DFF_4.Q ),
    .c(_311_),
    .y(_312_)
  );
  al_nand3ftt _369_ (
    .a(v2),
    .b(\DFF_4.Q ),
    .c(\DFF_3.Q ),
    .y(_313_)
  );
  al_oai21 _370_ (
    .a(v4),
    .b(v5),
    .c(\DFF_1.Q ),
    .y(_314_)
  );
  al_ao21 _371_ (
    .a(_313_),
    .b(_312_),
    .c(_314_),
    .y(_315_)
  );
  al_aoi21 _372_ (
    .a(_310_),
    .b(_315_),
    .c(_308_),
    .y(v13_D_18)
  );
  al_nor2 _373_ (
    .a(\DFF_5.Q ),
    .b(\DFF_4.Q ),
    .y(_316_)
  );
  al_inv _374_ (
    .a(_316_),
    .y(_317_)
  );
  al_and3fft _375_ (
    .a(\DFF_2.Q ),
    .b(\DFF_1.Q ),
    .c(v6),
    .y(_318_)
  );
  al_nand3ftt _376_ (
    .a(\DFF_3.Q ),
    .b(\DFF_0.Q ),
    .c(_318_),
    .y(_319_)
  );
  al_and2 _377_ (
    .a(\DFF_0.Q ),
    .b(\DFF_1.Q ),
    .y(_320_)
  );
  al_and2ft _378_ (
    .a(\DFF_0.Q ),
    .b(\DFF_1.Q ),
    .y(_321_)
  );
  al_nand3 _379_ (
    .a(v0),
    .b(_311_),
    .c(_321_),
    .y(_322_)
  );
  al_nand2 _380_ (
    .a(\DFF_3.Q ),
    .b(\DFF_2.Q ),
    .y(_323_)
  );
  al_aoi21ftf _381_ (
    .a(_323_),
    .b(_320_),
    .c(_322_),
    .y(_324_)
  );
  al_aoi21 _382_ (
    .a(_319_),
    .b(_324_),
    .c(_317_),
    .y(v13_D_23)
  );
  al_and2 _383_ (
    .a(\DFF_3.Q ),
    .b(\DFF_1.Q ),
    .y(_325_)
  );
  al_nand2ft _384_ (
    .a(v2),
    .b(\DFF_4.Q ),
    .y(_326_)
  );
  al_oai21ftt _385_ (
    .a(\DFF_2.Q ),
    .b(v0),
    .c(\DFF_1.Q ),
    .y(_327_)
  );
  al_nand3fft _386_ (
    .a(\DFF_4.Q ),
    .b(\DFF_3.Q ),
    .c(_327_),
    .y(_328_)
  );
  al_ao21ftf _387_ (
    .a(_326_),
    .b(_325_),
    .c(_328_),
    .y(_329_)
  );
  al_and2ft _388_ (
    .a(\DFF_1.Q ),
    .b(\DFF_2.Q ),
    .y(_330_)
  );
  al_inv _389_ (
    .a(_330_),
    .y(_331_)
  );
  al_and3ftt _390_ (
    .a(v5),
    .b(v4),
    .c(_307_),
    .y(_332_)
  );
  al_and3 _391_ (
    .a(_332_),
    .b(_331_),
    .c(_329_),
    .y(v13_D_15)
  );
  al_or2 _392_ (
    .a(\DFF_2.Q ),
    .b(\DFF_1.Q ),
    .y(_333_)
  );
  al_nand3 _393_ (
    .a(\DFF_5.Q ),
    .b(\DFF_4.Q ),
    .c(_333_),
    .y(_334_)
  );
  al_nand3ftt _394_ (
    .a(\DFF_4.Q ),
    .b(\DFF_2.Q ),
    .c(\DFF_1.Q ),
    .y(_335_)
  );
  al_ao21ttf _395_ (
    .a(_335_),
    .b(_334_),
    .c(\DFF_3.Q ),
    .y(_336_)
  );
  al_inv _396_ (
    .a(\DFF_2.Q ),
    .y(_337_)
  );
  al_and3ftt _397_ (
    .a(\DFF_4.Q ),
    .b(v0),
    .c(\DFF_1.Q ),
    .y(_338_)
  );
  al_oai21ttf _398_ (
    .a(\DFF_3.Q ),
    .b(_326_),
    .c(_338_),
    .y(_339_)
  );
  al_nand3fft _399_ (
    .a(\DFF_5.Q ),
    .b(_337_),
    .c(_339_),
    .y(_340_)
  );
  al_aoi21 _400_ (
    .a(_336_),
    .b(_340_),
    .c(\DFF_0.Q ),
    .y(v13_D_9)
  );
  al_inv _401_ (
    .a(CLR),
    .y(_341_)
  );
  al_and2ft _402_ (
    .a(\DFF_5.Q ),
    .b(\DFF_3.Q ),
    .y(_000_)
  );
  al_ao21ttf _403_ (
    .a(v3),
    .b(_283_),
    .c(_320_),
    .y(_001_)
  );
  al_aoi21 _404_ (
    .a(v1),
    .b(v3),
    .c(\DFF_1.Q ),
    .y(_002_)
  );
  al_nand3fft _405_ (
    .a(\DFF_4.Q ),
    .b(\DFF_0.Q ),
    .c(_002_),
    .y(_003_)
  );
  al_and3ftt _406_ (
    .a(\DFF_1.Q ),
    .b(\DFF_4.Q ),
    .c(\DFF_0.Q ),
    .y(_004_)
  );
  al_nand2ft _407_ (
    .a(\DFF_2.Q ),
    .b(\DFF_0.Q ),
    .y(_005_)
  );
  al_and3ftt _408_ (
    .a(_004_),
    .b(_005_),
    .c(_003_),
    .y(_006_)
  );
  al_ao21ttf _409_ (
    .a(_001_),
    .b(_006_),
    .c(_000_),
    .y(_007_)
  );
  al_nor2 _410_ (
    .a(\DFF_0.Q ),
    .b(\DFF_3.Q ),
    .y(_008_)
  );
  al_and3 _411_ (
    .a(v4),
    .b(v5),
    .c(_008_),
    .y(_009_)
  );
  al_nand2ft _412_ (
    .a(v0),
    .b(\DFF_1.Q ),
    .y(_010_)
  );
  al_nand3ftt _413_ (
    .a(_010_),
    .b(\DFF_2.Q ),
    .c(_009_),
    .y(_011_)
  );
  al_oai21ttf _414_ (
    .a(v6),
    .b(\DFF_0.Q ),
    .c(\DFF_1.Q ),
    .y(_012_)
  );
  al_oai21ftt _415_ (
    .a(\DFF_2.Q ),
    .b(\DFF_0.Q ),
    .c(\DFF_3.Q ),
    .y(_013_)
  );
  al_and2ft _416_ (
    .a(\DFF_0.Q ),
    .b(\DFF_2.Q ),
    .y(_014_)
  );
  al_nand3ftt _417_ (
    .a(\DFF_1.Q ),
    .b(\DFF_3.Q ),
    .c(_014_),
    .y(_015_)
  );
  al_aoi21ftf _418_ (
    .a(_013_),
    .b(_012_),
    .c(_015_),
    .y(_016_)
  );
  al_ao21 _419_ (
    .a(_011_),
    .b(_016_),
    .c(_317_),
    .y(_017_)
  );
  al_and2ft _420_ (
    .a(v2),
    .b(\DFF_3.Q ),
    .y(_018_)
  );
  al_and2 _421_ (
    .a(\DFF_4.Q ),
    .b(\DFF_1.Q ),
    .y(_019_)
  );
  al_and2 _422_ (
    .a(v4),
    .b(v5),
    .y(_020_)
  );
  al_ao21ttf _423_ (
    .a(_019_),
    .b(_020_),
    .c(_297_),
    .y(_021_)
  );
  al_nand3 _424_ (
    .a(_307_),
    .b(_018_),
    .c(_021_),
    .y(_022_)
  );
  al_and2 _425_ (
    .a(\DFF_5.Q ),
    .b(\DFF_4.Q ),
    .y(_023_)
  );
  al_and3ftt _426_ (
    .a(v2),
    .b(_302_),
    .c(_023_),
    .y(_024_)
  );
  al_nand2ft _427_ (
    .a(\DFF_1.Q ),
    .b(\DFF_3.Q ),
    .y(_025_)
  );
  al_ao21ftf _428_ (
    .a(\DFF_3.Q ),
    .b(\DFF_0.Q ),
    .c(_025_),
    .y(_026_)
  );
  al_nand2 _429_ (
    .a(\DFF_2.Q ),
    .b(\DFF_1.Q ),
    .y(_027_)
  );
  al_and3 _430_ (
    .a(_323_),
    .b(_027_),
    .c(_023_),
    .y(_028_)
  );
  al_aoi21 _431_ (
    .a(_026_),
    .b(_028_),
    .c(_024_),
    .y(_029_)
  );
  al_and3 _432_ (
    .a(_022_),
    .b(_029_),
    .c(_017_),
    .y(_030_)
  );
  al_aoi21 _433_ (
    .a(_007_),
    .b(_030_),
    .c(_341_),
    .y(\DFF_5.D )
  );
  al_nand3ftt _434_ (
    .a(v1),
    .b(v0),
    .c(v6),
    .y(_031_)
  );
  al_ao21ttf _435_ (
    .a(_031_),
    .b(_291_),
    .c(_025_),
    .y(_032_)
  );
  al_aoi21 _436_ (
    .a(\DFF_2.Q ),
    .b(\DFF_1.Q ),
    .c(\DFF_3.Q ),
    .y(_033_)
  );
  al_nand3ftt _437_ (
    .a(\DFF_0.Q ),
    .b(v2),
    .c(\DFF_2.Q ),
    .y(_034_)
  );
  al_nand3ftt _438_ (
    .a(\DFF_2.Q ),
    .b(\DFF_0.Q ),
    .c(\DFF_1.Q ),
    .y(_035_)
  );
  al_ao21ttf _439_ (
    .a(_034_),
    .b(_033_),
    .c(_035_),
    .y(_036_)
  );
  al_ao21 _440_ (
    .a(_012_),
    .b(_032_),
    .c(_036_),
    .y(_037_)
  );
  al_nand2 _441_ (
    .a(\DFF_4.Q ),
    .b(_037_),
    .y(_038_)
  );
  al_and2ft _442_ (
    .a(\DFF_4.Q ),
    .b(\DFF_0.Q ),
    .y(_039_)
  );
  al_ao21 _443_ (
    .a(\DFF_3.Q ),
    .b(\DFF_2.Q ),
    .c(_033_),
    .y(_040_)
  );
  al_ao21ftf _444_ (
    .a(_318_),
    .b(_040_),
    .c(_039_),
    .y(_041_)
  );
  al_nand2ft _445_ (
    .a(\DFF_0.Q ),
    .b(\DFF_4.Q ),
    .y(_042_)
  );
  al_or2 _446_ (
    .a(\DFF_0.Q ),
    .b(\DFF_3.Q ),
    .y(_043_)
  );
  al_nand3fft _447_ (
    .a(v3),
    .b(\DFF_1.Q ),
    .c(_043_),
    .y(_044_)
  );
  al_ao21 _448_ (
    .a(_005_),
    .b(_042_),
    .c(_044_),
    .y(_045_)
  );
  al_nand2ft _449_ (
    .a(\DFF_2.Q ),
    .b(\DFF_4.Q ),
    .y(_046_)
  );
  al_aoi21ftf _450_ (
    .a(_046_),
    .b(_296_),
    .c(_045_),
    .y(_047_)
  );
  al_aoi21 _451_ (
    .a(\DFF_3.Q ),
    .b(\DFF_2.Q ),
    .c(\DFF_4.Q ),
    .y(_048_)
  );
  al_nand2 _452_ (
    .a(\DFF_4.Q ),
    .b(\DFF_2.Q ),
    .y(_049_)
  );
  al_and3ftt _453_ (
    .a(\DFF_0.Q ),
    .b(v2),
    .c(_049_),
    .y(_050_)
  );
  al_nand3fft _454_ (
    .a(_333_),
    .b(_296_),
    .c(_008_),
    .y(_051_)
  );
  al_aoi21ftf _455_ (
    .a(_048_),
    .b(_050_),
    .c(_051_),
    .y(_052_)
  );
  al_and3 _456_ (
    .a(_041_),
    .b(_052_),
    .c(_047_),
    .y(_053_)
  );
  al_ao21 _457_ (
    .a(_038_),
    .b(_053_),
    .c(\DFF_5.Q ),
    .y(_054_)
  );
  al_nand3 _458_ (
    .a(\DFF_5.Q ),
    .b(\DFF_3.Q ),
    .c(_321_),
    .y(_055_)
  );
  al_and3fft _459_ (
    .a(\DFF_3.Q ),
    .b(\DFF_2.Q ),
    .c(\DFF_0.Q ),
    .y(_056_)
  );
  al_nand2ft _460_ (
    .a(\DFF_3.Q ),
    .b(\DFF_0.Q ),
    .y(_057_)
  );
  al_nand2ft _461_ (
    .a(\DFF_1.Q ),
    .b(\DFF_4.Q ),
    .y(_058_)
  );
  al_aoi21 _462_ (
    .a(\DFF_2.Q ),
    .b(_057_),
    .c(_058_),
    .y(_059_)
  );
  al_aoi21ftf _463_ (
    .a(_056_),
    .b(_059_),
    .c(_055_),
    .y(_060_)
  );
  al_aoi21 _464_ (
    .a(_060_),
    .b(_054_),
    .c(_341_),
    .y(\DFF_2.D )
  );
  al_inv _465_ (
    .a(\DFF_4.Q ),
    .y(_061_)
  );
  al_nor2 _466_ (
    .a(\DFF_2.Q ),
    .b(\DFF_1.Q ),
    .y(_062_)
  );
  al_oai21 _467_ (
    .a(v3),
    .b(v6),
    .c(_062_),
    .y(_063_)
  );
  al_nand3 _468_ (
    .a(\DFF_0.Q ),
    .b(_027_),
    .c(_063_),
    .y(_064_)
  );
  al_nand3ftt _469_ (
    .a(\DFF_0.Q ),
    .b(v4),
    .c(v5),
    .y(_065_)
  );
  al_and3fft _470_ (
    .a(_065_),
    .b(_330_),
    .c(_327_),
    .y(_066_)
  );
  al_ao21ftf _471_ (
    .a(_066_),
    .b(_064_),
    .c(_061_),
    .y(_067_)
  );
  al_nand3 _472_ (
    .a(\DFF_0.Q ),
    .b(\DFF_3.Q ),
    .c(\DFF_1.Q ),
    .y(_068_)
  );
  al_or3ftt _473_ (
    .a(\DFF_1.Q ),
    .b(v1),
    .c(_005_),
    .y(_069_)
  );
  al_and3ftt _474_ (
    .a(\DFF_4.Q ),
    .b(\DFF_0.Q ),
    .c(\DFF_2.Q ),
    .y(_070_)
  );
  al_nand2ft _475_ (
    .a(\DFF_4.Q ),
    .b(\DFF_3.Q ),
    .y(_071_)
  );
  al_aoi21ftf _476_ (
    .a(v3),
    .b(_070_),
    .c(_071_),
    .y(_072_)
  );
  al_ao21 _477_ (
    .a(_069_),
    .b(_072_),
    .c(_294_),
    .y(_073_)
  );
  al_or3ftt _478_ (
    .a(\DFF_2.Q ),
    .b(\DFF_0.Q ),
    .c(\DFF_1.Q ),
    .y(_074_)
  );
  al_nand3ftt _479_ (
    .a(\DFF_0.Q ),
    .b(\DFF_4.Q ),
    .c(_309_),
    .y(_075_)
  );
  al_aoi21ftf _480_ (
    .a(_071_),
    .b(_074_),
    .c(_075_),
    .y(_076_)
  );
  al_and3 _481_ (
    .a(_068_),
    .b(_076_),
    .c(_073_),
    .y(_077_)
  );
  al_ao21 _482_ (
    .a(_067_),
    .b(_077_),
    .c(\DFF_5.Q ),
    .y(_078_)
  );
  al_nand3ftt _483_ (
    .a(\DFF_2.Q ),
    .b(v1),
    .c(\DFF_0.Q ),
    .y(_079_)
  );
  al_or3fft _484_ (
    .a(v4),
    .b(v5),
    .c(_042_),
    .y(_080_)
  );
  al_ao21 _485_ (
    .a(_079_),
    .b(_080_),
    .c(_292_),
    .y(_081_)
  );
  al_nand2 _486_ (
    .a(\DFF_4.Q ),
    .b(\DFF_1.Q ),
    .y(_082_)
  );
  al_nand3 _487_ (
    .a(\DFF_5.Q ),
    .b(\DFF_4.Q ),
    .c(_302_),
    .y(_083_)
  );
  al_aoi21ftf _488_ (
    .a(_082_),
    .b(_014_),
    .c(_083_),
    .y(_084_)
  );
  al_ao21 _489_ (
    .a(_084_),
    .b(_081_),
    .c(v2),
    .y(_085_)
  );
  al_nand3 _490_ (
    .a(\DFF_3.Q ),
    .b(\DFF_1.Q ),
    .c(_014_),
    .y(_086_)
  );
  al_nand3fft _491_ (
    .a(\DFF_4.Q ),
    .b(\DFF_2.Q ),
    .c(_321_),
    .y(_087_)
  );
  al_aoi21ftf _492_ (
    .a(_082_),
    .b(_014_),
    .c(_087_),
    .y(_088_)
  );
  al_ao21 _493_ (
    .a(_086_),
    .b(_088_),
    .c(_293_),
    .y(_089_)
  );
  al_oai21ftt _494_ (
    .a(_333_),
    .b(_056_),
    .c(_023_),
    .y(_090_)
  );
  al_ao21ftf _495_ (
    .a(\DFF_0.Q ),
    .b(v3),
    .c(_057_),
    .y(_091_)
  );
  al_aoi21ttf _496_ (
    .a(_091_),
    .b(_059_),
    .c(_090_),
    .y(_092_)
  );
  al_and3 _497_ (
    .a(_092_),
    .b(_089_),
    .c(_085_),
    .y(_093_)
  );
  al_aoi21 _498_ (
    .a(_093_),
    .b(_078_),
    .c(_341_),
    .y(\DFF_4.D )
  );
  al_nand3 _499_ (
    .a(\DFF_2.Q ),
    .b(_018_),
    .c(_296_),
    .y(_094_)
  );
  al_oai21ftt _500_ (
    .a(\DFF_1.Q ),
    .b(\DFF_0.Q ),
    .c(\DFF_3.Q ),
    .y(_095_)
  );
  al_oai21 _501_ (
    .a(\DFF_3.Q ),
    .b(\DFF_2.Q ),
    .c(\DFF_4.Q ),
    .y(_096_)
  );
  al_nand3ftt _502_ (
    .a(_096_),
    .b(_095_),
    .c(_094_),
    .y(_097_)
  );
  al_nand3fft _503_ (
    .a(\DFF_4.Q ),
    .b(_057_),
    .c(_318_),
    .y(_098_)
  );
  al_and2ft _504_ (
    .a(\DFF_4.Q ),
    .b(\DFF_3.Q ),
    .y(_099_)
  );
  al_nand3fft _505_ (
    .a(\DFF_0.Q ),
    .b(\DFF_3.Q ),
    .c(_330_),
    .y(_100_)
  );
  al_aoi21ftf _506_ (
    .a(_027_),
    .b(_099_),
    .c(_100_),
    .y(_101_)
  );
  al_and3 _507_ (
    .a(_098_),
    .b(_101_),
    .c(_097_),
    .y(_102_)
  );
  al_nand2 _508_ (
    .a(v3),
    .b(\DFF_0.Q ),
    .y(_103_)
  );
  al_and2ft _509_ (
    .a(v0),
    .b(\DFF_2.Q ),
    .y(_104_)
  );
  al_nand3fft _510_ (
    .a(_283_),
    .b(_103_),
    .c(_019_),
    .y(_105_)
  );
  al_ao21ftf _511_ (
    .a(_009_),
    .b(_105_),
    .c(_104_),
    .y(_106_)
  );
  al_and2 _512_ (
    .a(v0),
    .b(\DFF_1.Q ),
    .y(_107_)
  );
  al_nand3fft _513_ (
    .a(\DFF_4.Q ),
    .b(\DFF_3.Q ),
    .c(_062_),
    .y(_108_)
  );
  al_ao21ttf _514_ (
    .a(_107_),
    .b(_290_),
    .c(_108_),
    .y(_109_)
  );
  al_aoi21ftf _515_ (
    .a(_103_),
    .b(_109_),
    .c(_106_),
    .y(_110_)
  );
  al_ao21 _516_ (
    .a(_102_),
    .b(_110_),
    .c(\DFF_5.Q ),
    .y(_111_)
  );
  al_nand3 _517_ (
    .a(\DFF_4.Q ),
    .b(\DFF_1.Q ),
    .c(_311_),
    .y(_112_)
  );
  al_and3 _518_ (
    .a(v1),
    .b(v6),
    .c(_300_),
    .y(_113_)
  );
  al_nand3ftt _519_ (
    .a(_297_),
    .b(_000_),
    .c(_113_),
    .y(_114_)
  );
  al_ao21 _520_ (
    .a(_112_),
    .b(_114_),
    .c(v2),
    .y(_115_)
  );
  al_nand3ftt _521_ (
    .a(\DFF_1.Q ),
    .b(\DFF_4.Q ),
    .c(_043_),
    .y(_116_)
  );
  al_nand3fft _522_ (
    .a(\DFF_4.Q ),
    .b(\DFF_0.Q ),
    .c(\DFF_1.Q ),
    .y(_117_)
  );
  al_nand2ft _523_ (
    .a(\DFF_2.Q ),
    .b(\DFF_5.Q ),
    .y(_118_)
  );
  al_ao21 _524_ (
    .a(_117_),
    .b(_116_),
    .c(_118_),
    .y(_119_)
  );
  al_and3fft _525_ (
    .a(\DFF_0.Q ),
    .b(\DFF_3.Q ),
    .c(\DFF_4.Q ),
    .y(_120_)
  );
  al_ao21ftf _526_ (
    .a(_120_),
    .b(_055_),
    .c(\DFF_2.Q ),
    .y(_121_)
  );
  al_and3 _527_ (
    .a(_119_),
    .b(_121_),
    .c(_115_),
    .y(_122_)
  );
  al_aoi21 _528_ (
    .a(_122_),
    .b(_111_),
    .c(_341_),
    .y(\DFF_0.D )
  );
  al_and3ftt _529_ (
    .a(_300_),
    .b(_333_),
    .c(_027_),
    .y(_123_)
  );
  al_nand2 _530_ (
    .a(\DFF_3.Q ),
    .b(_123_),
    .y(_124_)
  );
  al_nand2 _531_ (
    .a(\DFF_0.Q ),
    .b(\DFF_3.Q ),
    .y(_125_)
  );
  al_or3ftt _532_ (
    .a(\DFF_3.Q ),
    .b(\DFF_4.Q ),
    .c(\DFF_2.Q ),
    .y(_126_)
  );
  al_ao21ftf _533_ (
    .a(\DFF_1.Q ),
    .b(\DFF_0.Q ),
    .c(_126_),
    .y(_127_)
  );
  al_nand3ftt _534_ (
    .a(v6),
    .b(_125_),
    .c(_127_),
    .y(_128_)
  );
  al_oai21 _535_ (
    .a(\DFF_0.Q ),
    .b(\DFF_3.Q ),
    .c(_065_),
    .y(_129_)
  );
  al_nand3fft _536_ (
    .a(_309_),
    .b(_326_),
    .c(_129_),
    .y(_130_)
  );
  al_and3 _537_ (
    .a(_130_),
    .b(_128_),
    .c(_124_),
    .y(_131_)
  );
  al_and3ftt _538_ (
    .a(\DFF_1.Q ),
    .b(\DFF_0.Q ),
    .c(\DFF_2.Q ),
    .y(_132_)
  );
  al_nand2 _539_ (
    .a(v1),
    .b(\DFF_3.Q ),
    .y(_133_)
  );
  al_nand3fft _540_ (
    .a(\DFF_4.Q ),
    .b(\DFF_0.Q ),
    .c(_133_),
    .y(_134_)
  );
  al_oa21ttf _541_ (
    .a(_134_),
    .b(_040_),
    .c(_132_),
    .y(_135_)
  );
  al_nand2ft _542_ (
    .a(\DFF_0.Q ),
    .b(\DFF_1.Q ),
    .y(_136_)
  );
  al_or3 _543_ (
    .a(v3),
    .b(\DFF_3.Q ),
    .c(\DFF_2.Q ),
    .y(_137_)
  );
  al_aoi21ftf _544_ (
    .a(\DFF_2.Q ),
    .b(_136_),
    .c(_137_),
    .y(_138_)
  );
  al_ao21ttf _545_ (
    .a(_291_),
    .b(_031_),
    .c(_138_),
    .y(_139_)
  );
  al_aoi21ftf _546_ (
    .a(_061_),
    .b(_139_),
    .c(_135_),
    .y(_140_)
  );
  al_ao21 _547_ (
    .a(_131_),
    .b(_140_),
    .c(\DFF_5.Q ),
    .y(_141_)
  );
  al_and2ft _548_ (
    .a(_301_),
    .b(_303_),
    .y(_142_)
  );
  al_oai21ftf _549_ (
    .a(\DFF_3.Q ),
    .b(_117_),
    .c(_004_),
    .y(_143_)
  );
  al_and3 _550_ (
    .a(v2),
    .b(_000_),
    .c(_300_),
    .y(_144_)
  );
  al_aoi21 _551_ (
    .a(_337_),
    .b(_143_),
    .c(_144_),
    .y(_145_)
  );
  al_nand2ft _552_ (
    .a(\DFF_0.Q ),
    .b(\DFF_5.Q ),
    .y(_146_)
  );
  al_nand3fft _553_ (
    .a(\DFF_4.Q ),
    .b(\DFF_2.Q ),
    .c(\DFF_1.Q ),
    .y(_147_)
  );
  al_nand3ftt _554_ (
    .a(\DFF_3.Q ),
    .b(\DFF_4.Q ),
    .c(_330_),
    .y(_148_)
  );
  al_ao21 _555_ (
    .a(_147_),
    .b(_148_),
    .c(_146_),
    .y(_149_)
  );
  al_and3ftt _556_ (
    .a(_142_),
    .b(_149_),
    .c(_145_),
    .y(_150_)
  );
  al_aoi21 _557_ (
    .a(_150_),
    .b(_141_),
    .c(_341_),
    .y(\DFF_1.D )
  );
  al_nand3fft _558_ (
    .a(\DFF_0.Q ),
    .b(\DFF_1.Q ),
    .c(_099_),
    .y(_151_)
  );
  al_or2 _559_ (
    .a(v1),
    .b(\DFF_3.Q ),
    .y(_152_)
  );
  al_nand3fft _560_ (
    .a(_008_),
    .b(_082_),
    .c(_152_),
    .y(_153_)
  );
  al_ao21 _561_ (
    .a(_151_),
    .b(_153_),
    .c(\DFF_2.Q ),
    .y(_154_)
  );
  al_ao21 _562_ (
    .a(_100_),
    .b(_154_),
    .c(_294_),
    .y(_155_)
  );
  al_nand2ft _563_ (
    .a(\DFF_0.Q ),
    .b(\DFF_2.Q ),
    .y(_156_)
  );
  al_or2 _564_ (
    .a(\DFF_4.Q ),
    .b(\DFF_3.Q ),
    .y(_157_)
  );
  al_ao21 _565_ (
    .a(_035_),
    .b(_156_),
    .c(_157_),
    .y(_158_)
  );
  al_nand3ftt _566_ (
    .a(_046_),
    .b(_296_),
    .c(_325_),
    .y(_159_)
  );
  al_and3ftt _567_ (
    .a(_010_),
    .b(_020_),
    .c(_005_),
    .y(_160_)
  );
  al_ao21 _568_ (
    .a(_159_),
    .b(_158_),
    .c(_160_),
    .y(_161_)
  );
  al_and2 _569_ (
    .a(\DFF_3.Q ),
    .b(_132_),
    .y(_162_)
  );
  al_or3 _570_ (
    .a(v1),
    .b(_035_),
    .c(_326_),
    .y(_163_)
  );
  al_nor2 _571_ (
    .a(v6),
    .b(\DFF_0.Q ),
    .y(_164_)
  );
  al_nand3ftt _572_ (
    .a(_071_),
    .b(_062_),
    .c(_164_),
    .y(_165_)
  );
  al_and3ftt _573_ (
    .a(_162_),
    .b(_163_),
    .c(_165_),
    .y(_166_)
  );
  al_nand3 _574_ (
    .a(\DFF_0.Q ),
    .b(\DFF_3.Q ),
    .c(_027_),
    .y(_167_)
  );
  al_and2ft _575_ (
    .a(\DFF_0.Q ),
    .b(v3),
    .y(_168_)
  );
  al_nand3fft _576_ (
    .a(\DFF_2.Q ),
    .b(\DFF_1.Q ),
    .c(_168_),
    .y(_169_)
  );
  al_ao21 _577_ (
    .a(_169_),
    .b(_167_),
    .c(_061_),
    .y(_170_)
  );
  al_or3ftt _578_ (
    .a(_337_),
    .b(v1),
    .c(_151_),
    .y(_171_)
  );
  al_and3 _579_ (
    .a(_051_),
    .b(_171_),
    .c(_170_),
    .y(_172_)
  );
  al_and3 _580_ (
    .a(_161_),
    .b(_166_),
    .c(_172_),
    .y(_173_)
  );
  al_ao21 _581_ (
    .a(_155_),
    .b(_173_),
    .c(\DFF_5.Q ),
    .y(_174_)
  );
  al_oai21ttf _582_ (
    .a(\DFF_2.Q ),
    .b(\DFF_1.Q ),
    .c(\DFF_0.Q ),
    .y(_175_)
  );
  al_nand3 _583_ (
    .a(v2),
    .b(\DFF_2.Q ),
    .c(\DFF_1.Q ),
    .y(_176_)
  );
  al_nand3ftt _584_ (
    .a(\DFF_3.Q ),
    .b(_333_),
    .c(_176_),
    .y(_177_)
  );
  al_ao21ttf _585_ (
    .a(_175_),
    .b(_177_),
    .c(_023_),
    .y(_178_)
  );
  al_nand3fft _586_ (
    .a(v6),
    .b(\DFF_4.Q ),
    .c(\DFF_0.Q ),
    .y(_179_)
  );
  al_or3 _587_ (
    .a(\DFF_5.Q ),
    .b(_179_),
    .c(_137_),
    .y(_180_)
  );
  al_or3fft _588_ (
    .a(\DFF_5.Q ),
    .b(_321_),
    .c(_311_),
    .y(_181_)
  );
  al_inv _589_ (
    .a(\DFF_1.Q ),
    .y(_182_)
  );
  al_ao21ftt _590_ (
    .a(_182_),
    .b(v3),
    .c(_075_),
    .y(_183_)
  );
  al_and3 _591_ (
    .a(_180_),
    .b(_181_),
    .c(_183_),
    .y(_184_)
  );
  al_and2 _592_ (
    .a(_178_),
    .b(_184_),
    .y(_185_)
  );
  al_aoi21 _593_ (
    .a(_185_),
    .b(_174_),
    .c(_341_),
    .y(\DFF_3.D )
  );
  al_and3ftt _594_ (
    .a(_025_),
    .b(_014_),
    .c(_023_),
    .y(_186_)
  );
  al_or2 _595_ (
    .a(\DFF_0.Q ),
    .b(v2),
    .y(_187_)
  );
  al_and3ftt _596_ (
    .a(\DFF_4.Q ),
    .b(\DFF_0.Q ),
    .c(\DFF_3.Q ),
    .y(_188_)
  );
  al_oai21ttf _597_ (
    .a(_058_),
    .b(_187_),
    .c(_188_),
    .y(_189_)
  );
  al_nor2 _598_ (
    .a(\DFF_5.Q ),
    .b(\DFF_2.Q ),
    .y(_190_)
  );
  al_ao21 _599_ (
    .a(_190_),
    .b(_189_),
    .c(_186_),
    .y(v13_D_22)
  );
  al_nand3ftt _600_ (
    .a(_179_),
    .b(_304_),
    .c(_309_),
    .y(_191_)
  );
  al_or3fft _601_ (
    .a(_191_),
    .b(_306_),
    .c(_142_),
    .y(v13_D_19)
  );
  al_and3fft _602_ (
    .a(\DFF_4.Q ),
    .b(_062_),
    .c(_010_),
    .y(_192_)
  );
  al_nand2 _603_ (
    .a(v3),
    .b(v6),
    .y(_193_)
  );
  al_mux2h _604_ (
    .a(_193_),
    .b(_020_),
    .s(_058_),
    .y(_194_)
  );
  al_nand3ftt _605_ (
    .a(\DFF_0.Q ),
    .b(_071_),
    .c(_301_),
    .y(_195_)
  );
  al_or3 _606_ (
    .a(_195_),
    .b(_192_),
    .c(_194_),
    .y(_196_)
  );
  al_aoi21ttf _607_ (
    .a(\DFF_3.Q ),
    .b(\DFF_2.Q ),
    .c(\DFF_4.Q ),
    .y(_197_)
  );
  al_ao21ftf _608_ (
    .a(_325_),
    .b(_197_),
    .c(_087_),
    .y(_198_)
  );
  al_ao21 _609_ (
    .a(_293_),
    .b(_196_),
    .c(_198_),
    .y(v13_D_11)
  );
  al_nand3ftt _610_ (
    .a(v2),
    .b(\DFF_3.Q ),
    .c(\DFF_1.Q ),
    .y(_199_)
  );
  al_and3ftt _611_ (
    .a(\DFF_1.Q ),
    .b(v2),
    .c(\DFF_2.Q ),
    .y(_200_)
  );
  al_nor3fft _612_ (
    .a(\DFF_4.Q ),
    .b(_199_),
    .c(_200_),
    .y(_201_)
  );
  al_ao21 _613_ (
    .a(\DFF_0.Q ),
    .b(\DFF_2.Q ),
    .c(\DFF_3.Q ),
    .y(_202_)
  );
  al_ao21ftf _614_ (
    .a(\DFF_0.Q ),
    .b(\DFF_1.Q ),
    .c(_202_),
    .y(_203_)
  );
  al_and2ft _615_ (
    .a(v4),
    .b(v5),
    .y(_204_)
  );
  al_aoi21ftf _616_ (
    .a(_204_),
    .b(_062_),
    .c(_203_),
    .y(_205_)
  );
  al_nand3fft _617_ (
    .a(_127_),
    .b(_201_),
    .c(_205_),
    .y(_206_)
  );
  al_nand3ftt _618_ (
    .a(\DFF_2.Q ),
    .b(\DFF_5.Q ),
    .c(_008_),
    .y(_207_)
  );
  al_mux2l _619_ (
    .a(_057_),
    .b(_125_),
    .s(_333_),
    .y(_208_)
  );
  al_aoi21 _620_ (
    .a(_207_),
    .b(_208_),
    .c(_061_),
    .y(_209_)
  );
  al_ao21 _621_ (
    .a(_293_),
    .b(_206_),
    .c(_209_),
    .y(v13_D_6)
  );
  al_ao21 _622_ (
    .a(\DFF_3.Q ),
    .b(\DFF_1.Q ),
    .c(_316_),
    .y(_210_)
  );
  al_and3 _623_ (
    .a(_020_),
    .b(_071_),
    .c(_210_),
    .y(_211_)
  );
  al_or2 _624_ (
    .a(_200_),
    .b(_192_),
    .y(_212_)
  );
  al_nor2 _625_ (
    .a(\DFF_5.Q ),
    .b(\DFF_3.Q ),
    .y(_213_)
  );
  al_ao21 _626_ (
    .a(_213_),
    .b(_212_),
    .c(_211_),
    .y(_214_)
  );
  al_aoi21ttf _627_ (
    .a(\DFF_0.Q ),
    .b(\DFF_3.Q ),
    .c(\DFF_1.Q ),
    .y(_215_)
  );
  al_or3fft _628_ (
    .a(_187_),
    .b(_215_),
    .c(_096_),
    .y(_216_)
  );
  al_oai21ftf _629_ (
    .a(_323_),
    .b(_309_),
    .c(_117_),
    .y(_217_)
  );
  al_oai21 _630_ (
    .a(\DFF_0.Q ),
    .b(\DFF_2.Q ),
    .c(_202_),
    .y(_218_)
  );
  al_and3ftt _631_ (
    .a(\DFF_1.Q ),
    .b(\DFF_5.Q ),
    .c(\DFF_4.Q ),
    .y(_219_)
  );
  al_or3fft _632_ (
    .a(\DFF_5.Q ),
    .b(_321_),
    .c(_096_),
    .y(_220_)
  );
  al_aoi21ttf _633_ (
    .a(_219_),
    .b(_218_),
    .c(_220_),
    .y(_221_)
  );
  al_and3 _634_ (
    .a(_216_),
    .b(_217_),
    .c(_221_),
    .y(_222_)
  );
  al_ao21ftf _635_ (
    .a(\DFF_0.Q ),
    .b(_214_),
    .c(_222_),
    .y(v13_D_10)
  );
  al_oai21ftt _636_ (
    .a(_156_),
    .b(_058_),
    .c(_005_),
    .y(_223_)
  );
  al_ao21ttf _637_ (
    .a(\DFF_1.Q ),
    .b(_309_),
    .c(_095_),
    .y(_224_)
  );
  al_nand2ft _638_ (
    .a(\DFF_4.Q ),
    .b(\DFF_1.Q ),
    .y(_225_)
  );
  al_oai21ftf _639_ (
    .a(_225_),
    .b(_018_),
    .c(_204_),
    .y(_226_)
  );
  al_aoi21ftf _640_ (
    .a(\DFF_0.Q ),
    .b(_200_),
    .c(_226_),
    .y(_227_)
  );
  al_nand3fft _641_ (
    .a(_223_),
    .b(_224_),
    .c(_227_),
    .y(_228_)
  );
  al_ao21 _642_ (
    .a(\DFF_0.Q ),
    .b(\DFF_1.Q ),
    .c(\DFF_3.Q ),
    .y(_229_)
  );
  al_oai21 _643_ (
    .a(\DFF_0.Q ),
    .b(\DFF_1.Q ),
    .c(_229_),
    .y(_230_)
  );
  al_nand3fft _644_ (
    .a(_293_),
    .b(_049_),
    .c(_230_),
    .y(_231_)
  );
  al_and3fft _645_ (
    .a(\DFF_0.Q ),
    .b(_147_),
    .c(\DFF_5.Q ),
    .y(_232_)
  );
  al_aoi21ftt _646_ (
    .a(_046_),
    .b(_026_),
    .c(_232_),
    .y(_233_)
  );
  al_aoi21ttf _647_ (
    .a(v0),
    .b(\DFF_1.Q ),
    .c(_074_),
    .y(_234_)
  );
  al_ao21ftf _648_ (
    .a(_229_),
    .b(_234_),
    .c(_316_),
    .y(_235_)
  );
  al_and3 _649_ (
    .a(_231_),
    .b(_233_),
    .c(_235_),
    .y(_236_)
  );
  al_ao21ttf _650_ (
    .a(_293_),
    .b(_228_),
    .c(_236_),
    .y(v13_D_8)
  );
  al_nand3fft _651_ (
    .a(v5),
    .b(\DFF_0.Q ),
    .c(\DFF_3.Q ),
    .y(_237_)
  );
  al_ao21ftt _652_ (
    .a(_237_),
    .b(_118_),
    .c(_303_),
    .y(_238_)
  );
  al_oa21ftf _653_ (
    .a(\DFF_2.Q ),
    .b(_295_),
    .c(_146_),
    .y(_239_)
  );
  al_ao21ftf _654_ (
    .a(\DFF_2.Q ),
    .b(_295_),
    .c(_239_),
    .y(_240_)
  );
  al_ao21ftf _655_ (
    .a(_326_),
    .b(_238_),
    .c(_240_),
    .y(_241_)
  );
  al_and3fft _656_ (
    .a(v5),
    .b(_027_),
    .c(_316_),
    .y(_242_)
  );
  al_oai21ttf _657_ (
    .a(_326_),
    .b(_118_),
    .c(_242_),
    .y(_243_)
  );
  al_nand3fft _658_ (
    .a(v0),
    .b(_043_),
    .c(_243_),
    .y(_244_)
  );
  al_nor2 _659_ (
    .a(v5),
    .b(\DFF_0.Q ),
    .y(_245_)
  );
  al_ao21 _660_ (
    .a(_333_),
    .b(_027_),
    .c(_245_),
    .y(_246_)
  );
  al_or3 _661_ (
    .a(\DFF_5.Q ),
    .b(\DFF_4.Q ),
    .c(\DFF_3.Q ),
    .y(_247_)
  );
  al_nand3ftt _662_ (
    .a(_247_),
    .b(_175_),
    .c(_246_),
    .y(_248_)
  );
  al_and3 _663_ (
    .a(_306_),
    .b(_248_),
    .c(_244_),
    .y(_249_)
  );
  al_ao21ftf _664_ (
    .a(_182_),
    .b(_241_),
    .c(_249_),
    .y(v13_D_24)
  );
  al_aoi21 _665_ (
    .a(\DFF_4.Q ),
    .b(v2),
    .c(\DFF_0.Q ),
    .y(_250_)
  );
  al_or2 _666_ (
    .a(v4),
    .b(v5),
    .y(_251_)
  );
  al_and3ftt _667_ (
    .a(_330_),
    .b(_296_),
    .c(_251_),
    .y(_252_)
  );
  al_ao21 _668_ (
    .a(_250_),
    .b(_252_),
    .c(\DFF_5.Q ),
    .y(_253_)
  );
  al_ao21ftf _669_ (
    .a(\DFF_3.Q ),
    .b(_327_),
    .c(_316_),
    .y(_254_)
  );
  al_nand3fft _670_ (
    .a(\DFF_4.Q ),
    .b(\DFF_3.Q ),
    .c(\DFF_2.Q ),
    .y(_255_)
  );
  al_nand3ftt _671_ (
    .a(_146_),
    .b(_297_),
    .c(_255_),
    .y(_256_)
  );
  al_aoi21ftf _672_ (
    .a(_325_),
    .b(_197_),
    .c(_256_),
    .y(_257_)
  );
  al_nand3 _673_ (
    .a(_254_),
    .b(_257_),
    .c(_253_),
    .y(v13_D_14)
  );
  al_ao21ftf _674_ (
    .a(_326_),
    .b(_325_),
    .c(_312_),
    .y(_258_)
  );
  al_nand3fft _675_ (
    .a(_204_),
    .b(_308_),
    .c(_258_),
    .y(_259_)
  );
  al_ao21 _676_ (
    .a(_035_),
    .b(_074_),
    .c(_157_),
    .y(_260_)
  );
  al_aoi21ftf _677_ (
    .a(_043_),
    .b(_200_),
    .c(_260_),
    .y(_261_)
  );
  al_or2 _678_ (
    .a(\DFF_5.Q ),
    .b(_261_),
    .y(_262_)
  );
  al_oa21ttf _679_ (
    .a(\DFF_3.Q ),
    .b(\DFF_2.Q ),
    .c(\DFF_0.Q ),
    .y(_263_)
  );
  al_oa21 _680_ (
    .a(_056_),
    .b(_263_),
    .c(_219_),
    .y(_264_)
  );
  al_aoi21ftt _681_ (
    .a(_055_),
    .b(_046_),
    .c(_264_),
    .y(_265_)
  );
  al_nand3 _682_ (
    .a(_259_),
    .b(_265_),
    .c(_262_),
    .y(v13_D_7)
  );
  al_nand3fft _683_ (
    .a(_156_),
    .b(_107_),
    .c(_213_),
    .y(_266_)
  );
  al_ao21 _684_ (
    .a(_323_),
    .b(_096_),
    .c(_136_),
    .y(_267_)
  );
  al_ao21 _685_ (
    .a(_266_),
    .b(_267_),
    .c(_294_),
    .y(_268_)
  );
  al_nand3 _686_ (
    .a(_316_),
    .b(_062_),
    .c(_009_),
    .y(_269_)
  );
  al_nand3fft _687_ (
    .a(\DFF_0.Q ),
    .b(\DFF_2.Q ),
    .c(\DFF_1.Q ),
    .y(_270_)
  );
  al_nand3 _688_ (
    .a(_042_),
    .b(_270_),
    .c(_112_),
    .y(_271_)
  );
  al_nand3fft _689_ (
    .a(_293_),
    .b(_294_),
    .c(_271_),
    .y(_272_)
  );
  al_nand3 _690_ (
    .a(_269_),
    .b(_268_),
    .c(_272_),
    .y(v13_D_17)
  );
  al_nand3 _691_ (
    .a(v4),
    .b(v5),
    .c(_300_),
    .y(_273_)
  );
  al_aoi21 _692_ (
    .a(v0),
    .b(_321_),
    .c(_132_),
    .y(_274_)
  );
  al_ao21 _693_ (
    .a(_273_),
    .b(_274_),
    .c(\DFF_3.Q ),
    .y(_275_)
  );
  al_ao21 _694_ (
    .a(_086_),
    .b(_275_),
    .c(_317_),
    .y(_276_)
  );
  al_or3 _695_ (
    .a(\DFF_3.Q ),
    .b(\DFF_2.Q ),
    .c(_117_),
    .y(_277_)
  );
  al_aoi21ftf _696_ (
    .a(_146_),
    .b(\DFF_4.Q ),
    .c(_216_),
    .y(_278_)
  );
  al_nand3 _697_ (
    .a(_277_),
    .b(_278_),
    .c(_276_),
    .y(v13_D_12)
  );
  al_nand2ft _698_ (
    .a(_065_),
    .b(_329_),
    .y(_279_)
  );
  al_aoi21ftf _699_ (
    .a(_301_),
    .b(_263_),
    .c(_100_),
    .y(_280_)
  );
  al_aoi21ftf _700_ (
    .a(_157_),
    .b(_123_),
    .c(_280_),
    .y(_281_)
  );
  al_ao21 _701_ (
    .a(_279_),
    .b(_281_),
    .c(\DFF_5.Q ),
    .y(_282_)
  );
  al_nand3 _702_ (
    .a(v1),
    .b(\DFF_3.Q ),
    .c(_321_),
    .y(_284_)
  );
  al_oai21ftf _703_ (
    .a(v1),
    .b(\DFF_0.Q ),
    .c(\DFF_3.Q ),
    .y(_285_)
  );
  al_oai21ftf _704_ (
    .a(_082_),
    .b(_307_),
    .c(_285_),
    .y(_286_)
  );
  al_ao21 _705_ (
    .a(_284_),
    .b(_286_),
    .c(_337_),
    .y(_287_)
  );
  al_nand3ftt _706_ (
    .a(_320_),
    .b(_309_),
    .c(_023_),
    .y(_288_)
  );
  al_and3fft _707_ (
    .a(_232_),
    .b(_186_),
    .c(_288_),
    .y(_289_)
  );
  al_nand3 _708_ (
    .a(_287_),
    .b(_289_),
    .c(_282_),
    .y(v13_D_13)
  );
  al_dffl _709_ (
    .clk(CK),
    .d(\DFF_0.D ),
    .q(\DFF_0.Q )
  );
  al_dffl _710_ (
    .clk(CK),
    .d(\DFF_1.D ),
    .q(\DFF_1.Q )
  );
  al_dffl _711_ (
    .clk(CK),
    .d(\DFF_2.D ),
    .q(\DFF_2.Q )
  );
  al_dffl _712_ (
    .clk(CK),
    .d(\DFF_3.D ),
    .q(\DFF_3.Q )
  );
  al_dffl _713_ (
    .clk(CK),
    .d(\DFF_4.D ),
    .q(\DFF_4.Q )
  );
  al_dffl _714_ (
    .clk(CK),
    .d(\DFF_5.D ),
    .q(\DFF_5.Q )
  );
  assign Av13_D_10B = v13_D_10;
  assign Av13_D_11B = v13_D_11;
  assign Av13_D_12B = v13_D_12;
  assign Av13_D_13B = v13_D_13;
  assign Av13_D_14B = v13_D_14;
  assign Av13_D_15B = v13_D_15;
  assign Av13_D_16B = v13_D_16;
  assign Av13_D_17B = v13_D_17;
  assign Av13_D_18B = v13_D_18;
  assign Av13_D_19B = v13_D_19;
  assign Av13_D_20B = v13_D_20;
  assign Av13_D_21B = v13_D_21;
  assign Av13_D_22B = v13_D_22;
  assign Av13_D_23B = v13_D_23;
  assign Av13_D_24B = v13_D_24;
  assign Av13_D_6B = v13_D_6;
  assign Av13_D_7B = v13_D_7;
  assign Av13_D_8B = v13_D_8;
  assign Av13_D_9B = v13_D_9;
  assign C193D = v2;
  assign C79D = \DFF_1.Q ;
  assign \DFF_0.CK  = CK;
  assign \DFF_1.CK  = CK;
  assign \DFF_2.CK  = CK;
  assign \DFF_3.CK  = CK;
  assign \DFF_4.CK  = CK;
  assign \DFF_5.CK  = CK;
  assign II143 = \DFF_2.Q ;
  assign IIII518 = \DFF_3.Q ;
  assign v10 = \DFF_2.Q ;
  assign v11 = \DFF_1.Q ;
  assign v12 = \DFF_0.Q ;
  assign v13_D_0C = \DFF_5.D ;
  assign v13_D_1C = \DFF_4.D ;
  assign v13_D_2C = \DFF_3.D ;
  assign v13_D_3C = \DFF_2.D ;
  assign v13_D_4C = \DFF_1.D ;
  assign v13_D_5C = \DFF_0.D ;
  assign v7 = \DFF_5.Q ;
  assign v8 = \DFF_4.Q ;
  assign v9 = \DFF_3.Q ;
endmodule
