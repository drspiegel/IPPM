
module s713(GND, VDD, CK, G1, G10, G100BF, G101BF, G103BF, G104BF, G105BF, G106BF, G107, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G4, G5, G6, G8, G83, G84, G85, G86BF, G87BF, G88BF, G89BF, G9, G90, G91, G92, G94, G95BF, G96BF, G97BF, G98BF, G99BF);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  input CK;
  wire \DFF_0.CK ;
  wire \DFF_0.D ;
  wire \DFF_0.Q ;
  wire \DFF_1.CK ;
  wire \DFF_1.D ;
  wire \DFF_1.Q ;
  wire \DFF_10.CK ;
  wire \DFF_10.D ;
  wire \DFF_10.Q ;
  wire \DFF_11.CK ;
  wire \DFF_11.D ;
  wire \DFF_11.Q ;
  wire \DFF_12.CK ;
  wire \DFF_12.D ;
  wire \DFF_12.Q ;
  wire \DFF_13.CK ;
  wire \DFF_13.D ;
  wire \DFF_13.Q ;
  wire \DFF_14.CK ;
  wire \DFF_14.D ;
  wire \DFF_14.Q ;
  wire \DFF_15.CK ;
  wire \DFF_15.D ;
  wire \DFF_15.Q ;
  wire \DFF_16.CK ;
  wire \DFF_16.D ;
  wire \DFF_16.Q ;
  wire \DFF_17.CK ;
  wire \DFF_17.D ;
  wire \DFF_17.Q ;
  wire \DFF_18.CK ;
  wire \DFF_18.D ;
  wire \DFF_18.Q ;
  wire \DFF_2.CK ;
  wire \DFF_2.D ;
  wire \DFF_2.Q ;
  wire \DFF_3.CK ;
  wire \DFF_3.D ;
  wire \DFF_3.Q ;
  wire \DFF_4.CK ;
  wire \DFF_4.D ;
  wire \DFF_4.Q ;
  wire \DFF_5.CK ;
  wire \DFF_5.D ;
  wire \DFF_5.Q ;
  wire \DFF_6.CK ;
  wire \DFF_6.D ;
  wire \DFF_6.Q ;
  wire \DFF_7.CK ;
  wire \DFF_7.D ;
  wire \DFF_7.Q ;
  wire \DFF_8.CK ;
  wire \DFF_8.D ;
  wire \DFF_8.Q ;
  wire \DFF_9.CK ;
  wire \DFF_9.D ;
  wire \DFF_9.Q ;
  input G1;
  input G10;
  output G100BF;
  output G101BF;
  output G103BF;
  output G104BF;
  output G105BF;
  output G106BF;
  output G107;
  wire G109;
  input G11;
  wire G111;
  wire G113;
  wire G115;
  wire G117;
  wire G119;
  input G12;
  wire G121;
  wire G122;
  wire G125;
  wire G126;
  wire G127;
  wire G128;
  wire G129;
  input G13;
  wire G130;
  wire G131;
  wire G132;
  wire G133;
  wire G138;
  wire G139;
  input G14;
  wire G140;
  wire G141;
  wire G142;
  input G15;
  wire G150;
  wire G158;
  input G16;
  input G17;
  input G18;
  input G19;
  input G2;
  input G20;
  wire G209;
  input G21;
  wire G211;
  wire G213;
  wire G215;
  wire G217;
  wire G219;
  input G22;
  wire G221;
  wire G223;
  wire G229;
  input G23;
  input G24;
  input G25;
  wire G250;
  input G26;
  wire G262;
  input G27;
  wire G271;
  wire G272;
  wire G273;
  wire G274;
  wire G275;
  wire G276;
  wire G277;
  wire G278;
  input G28;
  input G29;
  input G3;
  input G30;
  wire G300;
  wire G301;
  wire G306;
  wire G307;
  input G31;
  input G32;
  input G33;
  input G34;
  input G35;
  wire G352;
  wire G354;
  wire G356;
  wire G358;
  wire G359;
  input G36;
  wire G360;
  wire G361;
  wire G362;
  wire G363;
  wire G364;
  wire G367;
  wire G380;
  wire G386;
  wire G388;
  wire G389;
  wire G394;
  input G4;
  input G5;
  input G6;
  wire G64;
  wire G65;
  wire G66;
  wire G67;
  wire G68;
  wire G69;
  wire G70;
  wire G71;
  wire G72;
  wire G73;
  wire G74;
  wire G75;
  wire G76;
  wire G77;
  wire G78;
  wire G79;
  input G8;
  wire G80;
  wire G81;
  wire G82;
  output G83;
  output G84;
  output G85;
  output G86BF;
  output G87BF;
  output G88BF;
  output G89BF;
  input G9;
  output G90;
  output G91;
  output G92;
  output G94;
  output G95BF;
  output G96BF;
  output G97BF;
  output G98BF;
  output G99BF;
  input GND;
  wire II335;
  wire II338;
  wire II341;
  wire II449;
  wire II452;
  wire II524;
  wire II527;
  wire IIII398;
  wire IIII406;
  wire IIII414;
  wire IIII422;
  input VDD;
  al_nand3ftt _057_ (
    .a(G4),
    .b(\DFF_5.Q ),
    .c(G35),
    .y(G100BF)
  );
  al_nand3ftt _058_ (
    .a(G4),
    .b(\DFF_7.Q ),
    .c(G33),
    .y(G98BF)
  );
  al_nand3ftt _059_ (
    .a(G4),
    .b(\DFF_9.Q ),
    .c(G31),
    .y(G96BF)
  );
  al_and2ft _060_ (
    .a(G13),
    .b(G10),
    .y(_051_)
  );
  al_nand3ftt _061_ (
    .a(G3),
    .b(G9),
    .c(_051_),
    .y(_052_)
  );
  al_or2 _062_ (
    .a(G3),
    .b(G11),
    .y(_053_)
  );
  al_and3ftt _063_ (
    .a(\DFF_18.Q ),
    .b(G25),
    .c(_053_),
    .y(_054_)
  );
  al_nand2 _064_ (
    .a(_052_),
    .b(_054_),
    .y(G89BF)
  );
  al_nand3fft _065_ (
    .a(G3),
    .b(G9),
    .c(_051_),
    .y(_055_)
  );
  al_and2ft _066_ (
    .a(\DFF_16.Q ),
    .b(G23),
    .y(_056_)
  );
  al_nand3 _067_ (
    .a(_053_),
    .b(_056_),
    .c(_055_),
    .y(G87BF)
  );
  al_and3 _068_ (
    .a(\DFF_4.Q ),
    .b(_052_),
    .c(_054_),
    .y(\DFF_4.D )
  );
  al_nand2 _069_ (
    .a(G36),
    .b(\DFF_4.D ),
    .y(G101BF)
  );
  al_ao21 _070_ (
    .a(_052_),
    .b(_054_),
    .c(G3),
    .y(_000_)
  );
  al_nand3 _071_ (
    .a(\DFF_14.Q ),
    .b(G17),
    .c(_000_),
    .y(G106BF)
  );
  al_or3fft _072_ (
    .a(\DFF_8.Q ),
    .b(G32),
    .c(G87BF),
    .y(G97BF)
  );
  al_inv _073_ (
    .a(G3),
    .y(_001_)
  );
  al_inv _074_ (
    .a(\DFF_12.Q ),
    .y(_002_)
  );
  al_aoi21 _075_ (
    .a(_001_),
    .b(G87BF),
    .c(_002_),
    .y(_003_)
  );
  al_nand2 _076_ (
    .a(G15),
    .b(_003_),
    .y(G104BF)
  );
  al_and2ft _077_ (
    .a(G2),
    .b(\DFF_2.Q ),
    .y(_004_)
  );
  al_ao21ttf _078_ (
    .a(\DFF_14.Q ),
    .b(_000_),
    .c(_004_),
    .y(_005_)
  );
  al_and3fft _079_ (
    .a(G10),
    .b(G13),
    .c(G9),
    .y(_006_)
  );
  al_oa21 _080_ (
    .a(G3),
    .b(G11),
    .c(G24),
    .y(_007_)
  );
  al_aoi21ftf _081_ (
    .a(G3),
    .b(_006_),
    .c(_007_),
    .y(_008_)
  );
  al_nand2 _082_ (
    .a(_008_),
    .b(_005_),
    .y(G88BF)
  );
  al_or3fft _083_ (
    .a(\DFF_6.Q ),
    .b(G34),
    .c(G88BF),
    .y(G99BF)
  );
  al_aoi21ttf _084_ (
    .a(_001_),
    .b(G88BF),
    .c(\DFF_13.Q ),
    .y(\DFF_2.D )
  );
  al_ao21 _085_ (
    .a(_008_),
    .b(_005_),
    .c(G3),
    .y(_009_)
  );
  al_nand3 _086_ (
    .a(\DFF_13.Q ),
    .b(G16),
    .c(_009_),
    .y(G105BF)
  );
  al_inv _087_ (
    .a(_003_),
    .y(_010_)
  );
  al_and2 _088_ (
    .a(\DFF_14.Q ),
    .b(_000_),
    .y(_011_)
  );
  al_aoi21 _089_ (
    .a(\DFF_13.Q ),
    .b(_009_),
    .c(_011_),
    .y(_012_)
  );
  al_and2ft _090_ (
    .a(G2),
    .b(\DFF_0.Q ),
    .y(_013_)
  );
  al_nand3 _091_ (
    .a(_010_),
    .b(_013_),
    .c(_012_),
    .y(_014_)
  );
  al_nor2 _092_ (
    .a(G10),
    .b(G13),
    .y(_015_)
  );
  al_nand3fft _093_ (
    .a(G3),
    .b(G9),
    .c(_015_),
    .y(_016_)
  );
  al_and3 _094_ (
    .a(G22),
    .b(_053_),
    .c(_016_),
    .y(_017_)
  );
  al_nand2 _095_ (
    .a(_017_),
    .b(_014_),
    .y(G86BF)
  );
  al_and3 _096_ (
    .a(\DFF_10.Q ),
    .b(_017_),
    .c(_014_),
    .y(_018_)
  );
  al_nand2 _097_ (
    .a(G30),
    .b(_018_),
    .y(G95BF)
  );
  al_inv _098_ (
    .a(\DFF_11.Q ),
    .y(_019_)
  );
  al_aoi21 _099_ (
    .a(_001_),
    .b(G86BF),
    .c(_019_),
    .y(\DFF_0.D )
  );
  al_ao21 _100_ (
    .a(_017_),
    .b(_014_),
    .c(G3),
    .y(_020_)
  );
  al_nand3 _101_ (
    .a(\DFF_11.Q ),
    .b(G14),
    .c(_020_),
    .y(G103BF)
  );
  al_and2ft _102_ (
    .a(G4),
    .b(\DFF_7.Q ),
    .y(_021_)
  );
  al_oai21ftt _103_ (
    .a(\DFF_8.Q ),
    .b(G87BF),
    .c(_021_),
    .y(\DFF_8.D )
  );
  al_mux2l _104_ (
    .a(_021_),
    .b(\DFF_8.Q ),
    .s(G87BF),
    .y(\DFF_7.D )
  );
  al_and2ft _105_ (
    .a(G4),
    .b(\DFF_5.Q ),
    .y(_022_)
  );
  al_nand3 _106_ (
    .a(\DFF_6.Q ),
    .b(_008_),
    .c(_005_),
    .y(_023_)
  );
  al_nand2 _107_ (
    .a(_022_),
    .b(_023_),
    .y(\DFF_6.D )
  );
  al_ao21ttf _108_ (
    .a(_022_),
    .b(G88BF),
    .c(_023_),
    .y(\DFF_5.D )
  );
  al_or3ftt _109_ (
    .a(\DFF_9.Q ),
    .b(G4),
    .c(_018_),
    .y(\DFF_10.D )
  );
  al_and2ft _110_ (
    .a(G4),
    .b(\DFF_9.Q ),
    .y(_024_)
  );
  al_ao21 _111_ (
    .a(_024_),
    .b(G86BF),
    .c(_018_),
    .y(\DFF_9.D )
  );
  al_and3ftt _112_ (
    .a(G4),
    .b(\DFF_15.Q ),
    .c(G18),
    .y(G107)
  );
  al_and3ftt _113_ (
    .a(G4),
    .b(\DFF_16.Q ),
    .c(G19),
    .y(G83)
  );
  al_and3ftt _114_ (
    .a(G4),
    .b(\DFF_17.Q ),
    .c(G20),
    .y(G84)
  );
  al_and3ftt _115_ (
    .a(G4),
    .b(\DFF_18.Q ),
    .c(G21),
    .y(G85)
  );
  al_and2 _116_ (
    .a(G11),
    .b(G12),
    .y(_025_)
  );
  al_and3 _117_ (
    .a(G13),
    .b(G28),
    .c(_025_),
    .y(G92)
  );
  al_inv _118_ (
    .a(G2),
    .y(_026_)
  );
  al_and3 _119_ (
    .a(_026_),
    .b(\DFF_14.Q ),
    .c(_000_),
    .y(\DFF_18.D )
  );
  al_inv _120_ (
    .a(_011_),
    .y(_027_)
  );
  al_and3 _121_ (
    .a(_026_),
    .b(_027_),
    .c(\DFF_2.D ),
    .y(\DFF_17.D )
  );
  al_and3 _122_ (
    .a(_026_),
    .b(_003_),
    .c(_012_),
    .y(\DFF_16.D )
  );
  al_and3fft _123_ (
    .a(_003_),
    .b(\DFF_2.D ),
    .c(_027_),
    .y(_028_)
  );
  al_and3 _124_ (
    .a(_026_),
    .b(_028_),
    .c(\DFF_0.D ),
    .y(\DFF_15.D )
  );
  al_nor3fft _125_ (
    .a(\DFF_6.Q ),
    .b(_022_),
    .c(G88BF),
    .y(_029_)
  );
  al_inv _126_ (
    .a(_006_),
    .y(_030_)
  );
  al_nor3fft _127_ (
    .a(\DFF_8.Q ),
    .b(_021_),
    .c(G87BF),
    .y(_031_)
  );
  al_and3ftt _128_ (
    .a(G11),
    .b(\DFF_4.D ),
    .c(_031_),
    .y(_032_)
  );
  al_nand3 _129_ (
    .a(_024_),
    .b(_032_),
    .c(_018_),
    .y(_033_)
  );
  al_nand2 _130_ (
    .a(_030_),
    .b(_033_),
    .y(_034_)
  );
  al_and2ft _131_ (
    .a(G9),
    .b(_015_),
    .y(_035_)
  );
  al_nand3 _132_ (
    .a(_024_),
    .b(_035_),
    .c(_018_),
    .y(_036_)
  );
  al_oa21ftt _133_ (
    .a(G9),
    .b(\DFF_4.D ),
    .c(_051_),
    .y(_037_)
  );
  al_oai21 _134_ (
    .a(G9),
    .b(_031_),
    .c(_037_),
    .y(_038_)
  );
  al_and3 _135_ (
    .a(G12),
    .b(G26),
    .c(_038_),
    .y(_039_)
  );
  al_nand2 _136_ (
    .a(_039_),
    .b(_036_),
    .y(_040_)
  );
  al_aoi21 _137_ (
    .a(_029_),
    .b(_034_),
    .c(_040_),
    .y(G90)
  );
  al_nand3 _138_ (
    .a(_024_),
    .b(_028_),
    .c(_018_),
    .y(_041_)
  );
  al_nand3fft _139_ (
    .a(G2),
    .b(_019_),
    .c(_020_),
    .y(_042_)
  );
  al_nand2ft _140_ (
    .a(G8),
    .b(_042_),
    .y(_043_)
  );
  al_aoi21ftf _141_ (
    .a(\DFF_0.D ),
    .b(_041_),
    .c(_043_),
    .y(\DFF_11.D )
  );
  al_aoi21ftf _142_ (
    .a(G5),
    .b(G2),
    .c(_003_),
    .y(_044_)
  );
  al_and3 _143_ (
    .a(G5),
    .b(_031_),
    .c(_012_),
    .y(_045_)
  );
  al_oai21ftf _144_ (
    .a(_045_),
    .b(\DFF_0.D ),
    .c(_044_),
    .y(\DFF_12.D )
  );
  al_aoi21 _145_ (
    .a(\DFF_11.Q ),
    .b(_020_),
    .c(_003_),
    .y(_046_)
  );
  al_and3 _146_ (
    .a(G6),
    .b(_027_),
    .c(_029_),
    .y(_047_)
  );
  al_aoi21ftf _147_ (
    .a(G6),
    .b(G2),
    .c(\DFF_2.D ),
    .y(_048_)
  );
  al_ao21 _148_ (
    .a(_047_),
    .b(_046_),
    .c(_048_),
    .y(\DFF_13.D )
  );
  al_nor3fft _149_ (
    .a(G1),
    .b(\DFF_4.D ),
    .c(\DFF_2.D ),
    .y(_049_)
  );
  al_aoi21ftf _150_ (
    .a(G1),
    .b(G2),
    .c(_011_),
    .y(_050_)
  );
  al_ao21 _151_ (
    .a(_049_),
    .b(_046_),
    .c(_050_),
    .y(\DFF_14.D )
  );
  al_dffl _152_ (
    .clk(CK),
    .d(\DFF_0.D ),
    .q(\DFF_0.Q )
  );
  al_dffl _153_ (
    .clk(CK),
    .d(\DFF_2.D ),
    .q(\DFF_2.Q )
  );
  al_dffl _154_ (
    .clk(CK),
    .d(\DFF_4.D ),
    .q(\DFF_4.Q )
  );
  al_dffl _155_ (
    .clk(CK),
    .d(\DFF_5.D ),
    .q(\DFF_5.Q )
  );
  al_dffl _156_ (
    .clk(CK),
    .d(\DFF_6.D ),
    .q(\DFF_6.Q )
  );
  al_dffl _157_ (
    .clk(CK),
    .d(\DFF_7.D ),
    .q(\DFF_7.Q )
  );
  al_dffl _158_ (
    .clk(CK),
    .d(\DFF_8.D ),
    .q(\DFF_8.Q )
  );
  al_dffl _159_ (
    .clk(CK),
    .d(\DFF_9.D ),
    .q(\DFF_9.Q )
  );
  al_dffl _160_ (
    .clk(CK),
    .d(\DFF_10.D ),
    .q(\DFF_10.Q )
  );
  al_dffl _161_ (
    .clk(CK),
    .d(\DFF_11.D ),
    .q(\DFF_11.Q )
  );
  al_dffl _162_ (
    .clk(CK),
    .d(\DFF_12.D ),
    .q(\DFF_12.Q )
  );
  al_dffl _163_ (
    .clk(CK),
    .d(\DFF_13.D ),
    .q(\DFF_13.Q )
  );
  al_dffl _164_ (
    .clk(CK),
    .d(\DFF_14.D ),
    .q(\DFF_14.Q )
  );
  al_dffl _165_ (
    .clk(CK),
    .d(\DFF_15.D ),
    .q(\DFF_15.Q )
  );
  al_dffl _166_ (
    .clk(CK),
    .d(\DFF_16.D ),
    .q(\DFF_16.Q )
  );
  al_dffl _167_ (
    .clk(CK),
    .d(\DFF_17.D ),
    .q(\DFF_17.Q )
  );
  al_dffl _168_ (
    .clk(CK),
    .d(\DFF_18.D ),
    .q(\DFF_18.Q )
  );
  assign \DFF_0.CK  = CK;
  assign \DFF_1.CK  = CK;
  assign \DFF_1.D  = \DFF_16.D ;
  assign \DFF_1.Q  = \DFF_16.Q ;
  assign \DFF_10.CK  = CK;
  assign \DFF_11.CK  = CK;
  assign \DFF_12.CK  = CK;
  assign \DFF_13.CK  = CK;
  assign \DFF_14.CK  = CK;
  assign \DFF_15.CK  = CK;
  assign \DFF_16.CK  = CK;
  assign \DFF_17.CK  = CK;
  assign \DFF_18.CK  = CK;
  assign \DFF_2.CK  = CK;
  assign \DFF_3.CK  = CK;
  assign \DFF_3.D  = \DFF_18.D ;
  assign \DFF_3.Q  = \DFF_18.Q ;
  assign \DFF_4.CK  = CK;
  assign \DFF_5.CK  = CK;
  assign \DFF_6.CK  = CK;
  assign \DFF_7.CK  = CK;
  assign \DFF_8.CK  = CK;
  assign \DFF_9.CK  = CK;
  assign G109 = \DFF_4.Q ;
  assign G111 = \DFF_5.Q ;
  assign G113 = \DFF_6.Q ;
  assign G115 = \DFF_7.Q ;
  assign G117 = \DFF_8.Q ;
  assign G119 = \DFF_9.Q ;
  assign G121 = \DFF_10.Q ;
  assign G122 = \DFF_4.D ;
  assign G125 = \DFF_11.D ;
  assign G126 = \DFF_12.D ;
  assign G127 = \DFF_13.D ;
  assign G128 = \DFF_14.D ;
  assign G129 = \DFF_15.D ;
  assign G130 = \DFF_16.D ;
  assign G131 = \DFF_17.D ;
  assign G132 = \DFF_18.D ;
  assign G133 = \DFF_5.D ;
  assign G138 = \DFF_6.D ;
  assign G139 = \DFF_7.D ;
  assign G140 = \DFF_8.D ;
  assign G141 = \DFF_9.D ;
  assign G142 = \DFF_10.D ;
  assign G150 = \DFF_0.D ;
  assign G158 = \DFF_2.D ;
  assign G209 = \DFF_11.Q ;
  assign G211 = \DFF_12.Q ;
  assign G213 = \DFF_13.Q ;
  assign G215 = \DFF_14.Q ;
  assign G217 = \DFF_15.Q ;
  assign G219 = \DFF_16.Q ;
  assign G221 = \DFF_17.Q ;
  assign G223 = \DFF_18.Q ;
  assign G229 = \DFF_18.D ;
  assign G250 = \DFF_18.D ;
  assign G262 = \DFF_16.D ;
  assign G271 = \DFF_11.D ;
  assign G272 = \DFF_12.D ;
  assign G273 = \DFF_13.D ;
  assign G274 = \DFF_14.D ;
  assign G275 = \DFF_15.D ;
  assign G276 = \DFF_16.D ;
  assign G277 = \DFF_17.D ;
  assign G278 = \DFF_18.D ;
  assign G300 = \DFF_0.D ;
  assign G301 = \DFF_0.D ;
  assign G306 = \DFF_2.D ;
  assign G307 = \DFF_2.D ;
  assign G352 = G1;
  assign G354 = G86BF;
  assign G356 = G87BF;
  assign G358 = G88BF;
  assign G359 = G89BF;
  assign G360 = G4;
  assign G361 = G5;
  assign G362 = G6;
  assign G363 = G8;
  assign G364 = G9;
  assign G367 = G10;
  assign G380 = \DFF_0.D ;
  assign G386 = G11;
  assign G388 = G12;
  assign G389 = G13;
  assign G394 = \DFF_2.D ;
  assign G64 = \DFF_0.Q ;
  assign G65 = \DFF_16.Q ;
  assign G66 = \DFF_2.Q ;
  assign G67 = \DFF_18.Q ;
  assign G68 = \DFF_4.Q ;
  assign G69 = \DFF_5.Q ;
  assign G70 = \DFF_6.Q ;
  assign G71 = \DFF_7.Q ;
  assign G72 = \DFF_8.Q ;
  assign G73 = \DFF_9.Q ;
  assign G74 = \DFF_10.Q ;
  assign G75 = \DFF_11.Q ;
  assign G76 = \DFF_12.Q ;
  assign G77 = \DFF_13.Q ;
  assign G78 = \DFF_14.Q ;
  assign G79 = \DFF_15.Q ;
  assign G80 = \DFF_16.Q ;
  assign G81 = \DFF_17.Q ;
  assign G82 = \DFF_18.Q ;
  assign G91 = G27;
  assign G94 = G29;
  assign II335 = G87BF;
  assign II338 = G89BF;
  assign II341 = G87BF;
  assign II449 = G88BF;
  assign II452 = G88BF;
  assign II524 = G86BF;
  assign II527 = G86BF;
  assign IIII398 = G86BF;
  assign IIII406 = G87BF;
  assign IIII414 = G88BF;
  assign IIII422 = G89BF;
endmodule
