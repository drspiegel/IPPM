
module c432(N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  input N1;
  input N102;
  input N105;
  input N108;
  input N11;
  input N112;
  input N115;
  input N14;
  input N17;
  wire N203;
  input N21;
  wire N213;
  output N223;
  input N24;
  input N27;
  input N30;
  wire N309;
  wire N319;
  output N329;
  input N34;
  wire N360;
  input N37;
  output N370;
  input N4;
  input N40;
  output N421;
  input N43;
  output N430;
  output N431;
  output N432;
  input N47;
  input N50;
  input N53;
  input N56;
  input N60;
  input N63;
  input N66;
  input N69;
  input N73;
  input N76;
  input N79;
  input N8;
  input N82;
  input N86;
  input N89;
  input N92;
  input N95;
  input N99;
  al_nand2ft _097_ (
    .a(N24),
    .b(N30),
    .y(_043_)
  );
  al_ao21ftf _098_ (
    .a(N102),
    .b(N108),
    .c(_043_),
    .y(_044_)
  );
  al_and2ft _099_ (
    .a(N76),
    .b(N82),
    .y(_045_)
  );
  al_and2ft _100_ (
    .a(N1),
    .b(N4),
    .y(_046_)
  );
  al_nand2ft _101_ (
    .a(N89),
    .b(N95),
    .y(_047_)
  );
  al_nand3fft _102_ (
    .a(_045_),
    .b(_046_),
    .c(_047_),
    .y(_048_)
  );
  al_nand2ft _103_ (
    .a(N63),
    .b(N69),
    .y(_049_)
  );
  al_nand2ft _104_ (
    .a(N37),
    .b(N43),
    .y(_050_)
  );
  al_nand2ft _105_ (
    .a(N50),
    .b(N56),
    .y(_051_)
  );
  al_aoi21ftf _106_ (
    .a(N11),
    .b(N17),
    .c(_051_),
    .y(_052_)
  );
  al_and3 _107_ (
    .a(_049_),
    .b(_050_),
    .c(_052_),
    .y(_053_)
  );
  al_nand3fft _108_ (
    .a(_044_),
    .b(_048_),
    .c(_053_),
    .y(N223)
  );
  al_inv _109_ (
    .a(N69),
    .y(_054_)
  );
  al_and3ftt _110_ (
    .a(_045_),
    .b(_049_),
    .c(_050_),
    .y(_055_)
  );
  al_aoi21ftf _111_ (
    .a(N1),
    .b(N4),
    .c(_047_),
    .y(_056_)
  );
  al_and3ftt _112_ (
    .a(_044_),
    .b(_056_),
    .c(_052_),
    .y(_057_)
  );
  al_ao21ttf _113_ (
    .a(_055_),
    .b(_057_),
    .c(N63),
    .y(_058_)
  );
  al_nand3fft _114_ (
    .a(_054_),
    .b(N73),
    .c(_058_),
    .y(_059_)
  );
  al_ao21ttf _115_ (
    .a(N76),
    .b(N223),
    .c(N82),
    .y(_060_)
  );
  al_or2 _116_ (
    .a(N86),
    .b(_060_),
    .y(_061_)
  );
  al_aoi21ttf _117_ (
    .a(N24),
    .b(N223),
    .c(N30),
    .y(_062_)
  );
  al_inv _118_ (
    .a(N108),
    .y(_063_)
  );
  al_ao21ttf _119_ (
    .a(_055_),
    .b(_057_),
    .c(N102),
    .y(_064_)
  );
  al_nand3fft _120_ (
    .a(_063_),
    .b(N112),
    .c(_064_),
    .y(_065_)
  );
  al_aoi21ftf _121_ (
    .a(N34),
    .b(_062_),
    .c(_065_),
    .y(_066_)
  );
  al_nand3 _122_ (
    .a(_059_),
    .b(_061_),
    .c(_066_),
    .y(_067_)
  );
  al_inv _123_ (
    .a(N95),
    .y(_068_)
  );
  al_ao21ttf _124_ (
    .a(_055_),
    .b(_057_),
    .c(N89),
    .y(_069_)
  );
  al_nand3fft _125_ (
    .a(_068_),
    .b(N99),
    .c(_069_),
    .y(_070_)
  );
  al_inv _126_ (
    .a(N17),
    .y(_071_)
  );
  al_aoi21 _127_ (
    .a(N11),
    .b(N223),
    .c(_071_),
    .y(_072_)
  );
  al_nand2ft _128_ (
    .a(N21),
    .b(_072_),
    .y(_073_)
  );
  al_ao21ttf _129_ (
    .a(N1),
    .b(N223),
    .c(N4),
    .y(_074_)
  );
  al_or2 _130_ (
    .a(N8),
    .b(_074_),
    .y(_075_)
  );
  al_nand3 _131_ (
    .a(_070_),
    .b(_073_),
    .c(_075_),
    .y(_076_)
  );
  al_ao21ttf _132_ (
    .a(N37),
    .b(N223),
    .c(N43),
    .y(_077_)
  );
  al_inv _133_ (
    .a(N56),
    .y(_078_)
  );
  al_ao21ttf _134_ (
    .a(_055_),
    .b(_057_),
    .c(N50),
    .y(_079_)
  );
  al_nand3fft _135_ (
    .a(_078_),
    .b(N60),
    .c(_079_),
    .y(_080_)
  );
  al_oai21 _136_ (
    .a(N47),
    .b(_077_),
    .c(_080_),
    .y(_081_)
  );
  al_or3 _137_ (
    .a(_081_),
    .b(_076_),
    .c(_067_),
    .y(N329)
  );
  al_nand2ft _138_ (
    .a(N40),
    .b(_062_),
    .y(_082_)
  );
  al_aoi21 _139_ (
    .a(N34),
    .b(N329),
    .c(_082_),
    .y(_083_)
  );
  al_ao21ftf _140_ (
    .a(N21),
    .b(_072_),
    .c(_070_),
    .y(_084_)
  );
  al_nor3ftt _141_ (
    .a(_075_),
    .b(_084_),
    .c(_081_),
    .y(_085_)
  );
  al_nand3fft _142_ (
    .a(_060_),
    .b(_067_),
    .c(_085_),
    .y(_086_)
  );
  al_aoi21 _143_ (
    .a(_061_),
    .b(_086_),
    .c(N92),
    .y(_087_)
  );
  al_ao21 _144_ (
    .a(N63),
    .b(N223),
    .c(_054_),
    .y(_088_)
  );
  al_and3 _145_ (
    .a(_059_),
    .b(_061_),
    .c(_066_),
    .y(_089_)
  );
  al_ao21ttf _146_ (
    .a(_089_),
    .b(_085_),
    .c(N73),
    .y(_090_)
  );
  al_nand3fft _147_ (
    .a(N79),
    .b(_088_),
    .c(_090_),
    .y(_091_)
  );
  al_nand3fft _148_ (
    .a(_083_),
    .b(_087_),
    .c(_091_),
    .y(_092_)
  );
  al_inv _149_ (
    .a(N105),
    .y(_093_)
  );
  al_ao21ttf _150_ (
    .a(_089_),
    .b(_085_),
    .c(N8),
    .y(_094_)
  );
  al_nand3fft _151_ (
    .a(N14),
    .b(_074_),
    .c(_094_),
    .y(_095_)
  );
  al_ao21 _152_ (
    .a(N89),
    .b(N223),
    .c(_068_),
    .y(_096_)
  );
  al_aoi21 _153_ (
    .a(N99),
    .b(N329),
    .c(_096_),
    .y(_000_)
  );
  al_ao21ttf _154_ (
    .a(_093_),
    .b(_000_),
    .c(_095_),
    .y(_001_)
  );
  al_inv _155_ (
    .a(_072_),
    .y(_002_)
  );
  al_nand3fft _156_ (
    .a(_002_),
    .b(_067_),
    .c(_085_),
    .y(_003_)
  );
  al_nand2 _157_ (
    .a(_073_),
    .b(_003_),
    .y(_004_)
  );
  al_ao21 _158_ (
    .a(N102),
    .b(N223),
    .c(_063_),
    .y(_005_)
  );
  al_ao21ttf _159_ (
    .a(_089_),
    .b(_085_),
    .c(N112),
    .y(_006_)
  );
  al_nand3fft _160_ (
    .a(N115),
    .b(_005_),
    .c(_006_),
    .y(_007_)
  );
  al_aoi21ftf _161_ (
    .a(N27),
    .b(_004_),
    .c(_007_),
    .y(_008_)
  );
  al_ao21ttf _162_ (
    .a(_089_),
    .b(_085_),
    .c(N47),
    .y(_009_)
  );
  al_nand3fft _163_ (
    .a(N53),
    .b(_077_),
    .c(_009_),
    .y(_010_)
  );
  al_ao21 _164_ (
    .a(N50),
    .b(N223),
    .c(_078_),
    .y(_011_)
  );
  al_nand3fft _165_ (
    .a(_011_),
    .b(_067_),
    .c(_085_),
    .y(_012_)
  );
  al_ao21 _166_ (
    .a(_080_),
    .b(_012_),
    .c(N66),
    .y(_013_)
  );
  al_and3 _167_ (
    .a(_010_),
    .b(_013_),
    .c(_008_),
    .y(_014_)
  );
  al_nand3fft _168_ (
    .a(_092_),
    .b(_001_),
    .c(_014_),
    .y(N370)
  );
  al_ao21ttf _169_ (
    .a(N34),
    .b(N329),
    .c(_062_),
    .y(_015_)
  );
  al_ao21 _170_ (
    .a(N40),
    .b(N370),
    .c(_015_),
    .y(_016_)
  );
  al_ao21ttf _171_ (
    .a(N27),
    .b(N370),
    .c(_004_),
    .y(_017_)
  );
  al_ao21 _172_ (
    .a(N47),
    .b(N329),
    .c(_077_),
    .y(_018_)
  );
  al_ao21 _173_ (
    .a(N53),
    .b(N370),
    .c(_018_),
    .y(_019_)
  );
  al_and2 _174_ (
    .a(_080_),
    .b(_012_),
    .y(_020_)
  );
  al_and2 _175_ (
    .a(_061_),
    .b(_086_),
    .y(_021_)
  );
  al_oa21 _176_ (
    .a(N92),
    .b(_021_),
    .c(_010_),
    .y(_022_)
  );
  al_nand3ftt _177_ (
    .a(_083_),
    .b(_013_),
    .c(_022_),
    .y(_023_)
  );
  al_ao21ttf _178_ (
    .a(_093_),
    .b(_000_),
    .c(_091_),
    .y(_024_)
  );
  al_nor3fft _179_ (
    .a(_095_),
    .b(_008_),
    .c(_024_),
    .y(_025_)
  );
  al_nand3fft _180_ (
    .a(_020_),
    .b(_023_),
    .c(_025_),
    .y(_026_)
  );
  al_and3 _181_ (
    .a(_013_),
    .b(_026_),
    .c(_019_),
    .y(_027_)
  );
  al_and3 _182_ (
    .a(_016_),
    .b(_017_),
    .c(_027_),
    .y(_028_)
  );
  al_ao21 _183_ (
    .a(N73),
    .b(N329),
    .c(_088_),
    .y(_029_)
  );
  al_aoi21 _184_ (
    .a(N79),
    .b(N370),
    .c(_029_),
    .y(_030_)
  );
  al_and3fft _185_ (
    .a(_021_),
    .b(_023_),
    .c(_025_),
    .y(_031_)
  );
  al_or3 _186_ (
    .a(_087_),
    .b(_031_),
    .c(_030_),
    .y(_032_)
  );
  al_aoi21ttf _187_ (
    .a(N105),
    .b(N370),
    .c(_000_),
    .y(_033_)
  );
  al_ao21 _188_ (
    .a(N112),
    .b(N329),
    .c(_005_),
    .y(_034_)
  );
  al_ao21 _189_ (
    .a(N115),
    .b(N370),
    .c(_034_),
    .y(_035_)
  );
  al_and3fft _190_ (
    .a(_033_),
    .b(_032_),
    .c(_035_),
    .y(_036_)
  );
  al_ao21 _191_ (
    .a(N8),
    .b(N329),
    .c(_074_),
    .y(_037_)
  );
  al_aoi21 _192_ (
    .a(N14),
    .b(N370),
    .c(_037_),
    .y(_038_)
  );
  al_aoi21 _193_ (
    .a(_028_),
    .b(_036_),
    .c(_038_),
    .y(N421)
  );
  al_inv _194_ (
    .a(_028_),
    .y(N430)
  );
  al_and2 _195_ (
    .a(_016_),
    .b(_017_),
    .y(_039_)
  );
  al_ao21ttf _196_ (
    .a(_027_),
    .b(_032_),
    .c(_039_),
    .y(N431)
  );
  al_nand3fft _197_ (
    .a(_087_),
    .b(_031_),
    .c(_033_),
    .y(_040_)
  );
  al_nand3 _198_ (
    .a(_013_),
    .b(_026_),
    .c(_030_),
    .y(_041_)
  );
  al_nand3 _199_ (
    .a(_019_),
    .b(_040_),
    .c(_041_),
    .y(_042_)
  );
  al_ao21ttf _200_ (
    .a(_016_),
    .b(_042_),
    .c(_017_),
    .y(N432)
  );
  assign N203 = N223;
  assign N213 = N223;
  assign N309 = N329;
  assign N319 = N329;
  assign N360 = N370;
endmodule
