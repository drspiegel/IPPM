
module s526(GND, VDD, CK, G0, G1, G147, G148, G198, G199, G2, G213, G214);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  input CK;
  wire \DFF_0.CK ;
  wire \DFF_0.D ;
  wire \DFF_0.Q ;
  wire \DFF_1.CK ;
  wire \DFF_1.D ;
  wire \DFF_1.Q ;
  wire \DFF_10.CK ;
  wire \DFF_10.D ;
  wire \DFF_10.Q ;
  wire \DFF_11.CK ;
  wire \DFF_11.D ;
  wire \DFF_11.Q ;
  wire \DFF_12.CK ;
  wire \DFF_12.D ;
  wire \DFF_12.Q ;
  wire \DFF_13.CK ;
  wire \DFF_13.D ;
  wire \DFF_13.Q ;
  wire \DFF_14.CK ;
  wire \DFF_14.D ;
  wire \DFF_14.Q ;
  wire \DFF_15.CK ;
  wire \DFF_15.D ;
  wire \DFF_15.Q ;
  wire \DFF_16.CK ;
  wire \DFF_16.D ;
  wire \DFF_16.Q ;
  wire \DFF_17.CK ;
  wire \DFF_17.D ;
  wire \DFF_17.Q ;
  wire \DFF_18.CK ;
  wire \DFF_18.D ;
  wire \DFF_18.Q ;
  wire \DFF_19.CK ;
  wire \DFF_19.D ;
  wire \DFF_19.Q ;
  wire \DFF_2.CK ;
  wire \DFF_2.D ;
  wire \DFF_2.Q ;
  wire \DFF_20.CK ;
  wire \DFF_20.D ;
  wire \DFF_20.Q ;
  wire \DFF_3.CK ;
  wire \DFF_3.D ;
  wire \DFF_3.Q ;
  wire \DFF_4.CK ;
  wire \DFF_4.D ;
  wire \DFF_4.Q ;
  wire \DFF_5.CK ;
  wire \DFF_5.D ;
  wire \DFF_5.Q ;
  wire \DFF_6.CK ;
  wire \DFF_6.D ;
  wire \DFF_6.Q ;
  wire \DFF_7.CK ;
  wire \DFF_7.D ;
  wire \DFF_7.Q ;
  wire \DFF_8.CK ;
  wire \DFF_8.D ;
  wire \DFF_8.Q ;
  wire \DFF_9.CK ;
  wire \DFF_9.D ;
  wire \DFF_9.Q ;
  input G0;
  input G1;
  wire G10;
  wire G101;
  wire G106;
  wire G11;
  wire G115;
  wire G12;
  wire G126;
  wire G127;
  wire G13;
  wire G137;
  wire G14;
  output G147;
  output G148;
  wire G15;
  wire G16;
  wire G167;
  wire G17;
  wire G173;
  wire G179;
  wire G18;
  wire G183;
  wire G188;
  wire G19;
  wire G194;
  output G198;
  output G199;
  input G2;
  wire G20;
  wire G200;
  wire G205;
  wire G206;
  wire G21;
  wire G211;
  wire G212;
  output G213;
  output G214;
  wire G22;
  wire G23;
  wire G24;
  wire G25;
  wire G26;
  wire G27;
  wire G28;
  wire G29;
  wire G30;
  wire G60;
  wire G61;
  wire G62;
  wire G69;
  wire G79;
  wire G84;
  wire G89;
  wire G96;
  input GND;
  input VDD;
  al_inv _061_ (
    .a(G0),
    .y(_019_)
  );
  al_and2ft _062_ (
    .a(\DFF_1.Q ),
    .b(\DFF_0.Q ),
    .y(_020_)
  );
  al_and2ft _063_ (
    .a(\DFF_4.Q ),
    .b(\DFF_5.Q ),
    .y(_021_)
  );
  al_ao21 _064_ (
    .a(_020_),
    .b(_021_),
    .c(\DFF_20.Q ),
    .y(_022_)
  );
  al_and3fft _065_ (
    .a(\DFF_7.Q ),
    .b(\DFF_8.Q ),
    .c(\DFF_9.Q ),
    .y(_023_)
  );
  al_and3 _066_ (
    .a(\DFF_6.Q ),
    .b(_023_),
    .c(_022_),
    .y(_024_)
  );
  al_and2 _067_ (
    .a(\DFF_11.Q ),
    .b(\DFF_2.Q ),
    .y(_025_)
  );
  al_nand3 _068_ (
    .a(\DFF_10.Q ),
    .b(_025_),
    .c(_024_),
    .y(_026_)
  );
  al_inv _069_ (
    .a(\DFF_2.Q ),
    .y(_027_)
  );
  al_nand3 _070_ (
    .a(\DFF_10.Q ),
    .b(\DFF_11.Q ),
    .c(_024_),
    .y(_028_)
  );
  al_nand2 _071_ (
    .a(_027_),
    .b(_028_),
    .y(_029_)
  );
  al_and3 _072_ (
    .a(_019_),
    .b(_026_),
    .c(_029_),
    .y(\DFF_2.D )
  );
  al_inv _073_ (
    .a(\DFF_3.Q ),
    .y(_030_)
  );
  al_nand2 _074_ (
    .a(_030_),
    .b(_026_),
    .y(_031_)
  );
  al_or2 _075_ (
    .a(\DFF_11.Q ),
    .b(\DFF_2.Q ),
    .y(_032_)
  );
  al_oa21ftf _076_ (
    .a(_032_),
    .b(_025_),
    .c(_030_),
    .y(_033_)
  );
  al_nand3 _077_ (
    .a(\DFF_10.Q ),
    .b(_033_),
    .c(_024_),
    .y(_034_)
  );
  al_and3 _078_ (
    .a(_019_),
    .b(_034_),
    .c(_031_),
    .y(\DFF_3.D )
  );
  al_inv _079_ (
    .a(\DFF_11.Q ),
    .y(_035_)
  );
  al_nand2ft _080_ (
    .a(\DFF_2.Q ),
    .b(\DFF_3.Q ),
    .y(_036_)
  );
  al_nand3 _081_ (
    .a(\DFF_10.Q ),
    .b(_036_),
    .c(_024_),
    .y(_037_)
  );
  al_nand2 _082_ (
    .a(_035_),
    .b(_037_),
    .y(_038_)
  );
  al_and3 _083_ (
    .a(_019_),
    .b(_028_),
    .c(_038_),
    .y(\DFF_11.D )
  );
  al_nor2 _084_ (
    .a(\DFF_0.Q ),
    .b(G0),
    .y(\DFF_0.D )
  );
  al_and3fft _085_ (
    .a(\DFF_0.Q ),
    .b(G0),
    .c(\DFF_1.Q ),
    .y(_039_)
  );
  al_and3fft _086_ (
    .a(\DFF_1.Q ),
    .b(G0),
    .c(\DFF_0.Q ),
    .y(_040_)
  );
  al_oai21ftf _087_ (
    .a(_040_),
    .b(_021_),
    .c(_039_),
    .y(\DFF_1.D )
  );
  al_and3 _088_ (
    .a(\DFF_0.Q ),
    .b(\DFF_4.Q ),
    .c(\DFF_1.Q ),
    .y(_041_)
  );
  al_ao21 _089_ (
    .a(\DFF_0.Q ),
    .b(\DFF_1.Q ),
    .c(\DFF_4.Q ),
    .y(_042_)
  );
  al_and3fft _090_ (
    .a(G0),
    .b(_041_),
    .c(_042_),
    .y(\DFF_4.D )
  );
  al_or2ft _091_ (
    .a(\DFF_5.Q ),
    .b(_041_),
    .y(_043_)
  );
  al_nand2ft _092_ (
    .a(\DFF_5.Q ),
    .b(_041_),
    .y(_044_)
  );
  al_ao21ftf _093_ (
    .a(\DFF_4.Q ),
    .b(_020_),
    .c(_019_),
    .y(_045_)
  );
  al_aoi21 _094_ (
    .a(_044_),
    .b(_043_),
    .c(_045_),
    .y(\DFF_5.D )
  );
  al_and2 _095_ (
    .a(\DFF_6.Q ),
    .b(_022_),
    .y(_046_)
  );
  al_or2 _096_ (
    .a(\DFF_6.Q ),
    .b(_022_),
    .y(_047_)
  );
  al_nor3fft _097_ (
    .a(_019_),
    .b(_047_),
    .c(_046_),
    .y(\DFF_6.D )
  );
  al_aoi21 _098_ (
    .a(\DFF_6.Q ),
    .b(_022_),
    .c(\DFF_7.Q ),
    .y(_048_)
  );
  al_and3 _099_ (
    .a(\DFF_6.Q ),
    .b(\DFF_7.Q ),
    .c(_022_),
    .y(_049_)
  );
  al_nor2 _100_ (
    .a(G0),
    .b(_023_),
    .y(_050_)
  );
  al_nor3ftt _101_ (
    .a(_050_),
    .b(_049_),
    .c(_048_),
    .y(\DFF_7.D )
  );
  al_inv _102_ (
    .a(\DFF_8.Q ),
    .y(_051_)
  );
  al_oa21ftf _103_ (
    .a(_051_),
    .b(_049_),
    .c(G0),
    .y(_052_)
  );
  al_aoi21ftf _104_ (
    .a(_051_),
    .b(_049_),
    .c(_052_),
    .y(\DFF_8.D )
  );
  al_and3 _105_ (
    .a(\DFF_9.Q ),
    .b(\DFF_8.Q ),
    .c(_049_),
    .y(_053_)
  );
  al_nor2 _106_ (
    .a(\DFF_7.Q ),
    .b(\DFF_8.Q ),
    .y(_054_)
  );
  al_aoi21 _107_ (
    .a(_054_),
    .b(_046_),
    .c(G0),
    .y(_055_)
  );
  al_ao21 _108_ (
    .a(\DFF_8.Q ),
    .b(_049_),
    .c(\DFF_9.Q ),
    .y(_056_)
  );
  al_and3ftt _109_ (
    .a(_053_),
    .b(_056_),
    .c(_055_),
    .y(\DFF_9.D )
  );
  al_aoi21 _110_ (
    .a(\DFF_10.Q ),
    .b(_024_),
    .c(G0),
    .y(_057_)
  );
  al_oa21 _111_ (
    .a(\DFF_10.Q ),
    .b(_024_),
    .c(_057_),
    .y(\DFF_10.D )
  );
  al_and2ft _112_ (
    .a(\DFF_3.Q ),
    .b(\DFF_2.Q ),
    .y(_058_)
  );
  al_and2ft _113_ (
    .a(\DFF_11.Q ),
    .b(\DFF_10.Q ),
    .y(_059_)
  );
  al_ao21ttf _114_ (
    .a(_058_),
    .b(_059_),
    .c(\DFF_12.Q ),
    .y(_060_)
  );
  al_nor2 _115_ (
    .a(\DFF_10.Q ),
    .b(\DFF_11.Q ),
    .y(_000_)
  );
  al_ao21 _116_ (
    .a(_058_),
    .b(_000_),
    .c(\DFF_12.Q ),
    .y(_001_)
  );
  al_ao21ttf _117_ (
    .a(\DFF_19.Q ),
    .b(_001_),
    .c(_060_),
    .y(_002_)
  );
  al_and2 _118_ (
    .a(_019_),
    .b(_002_),
    .y(\DFF_12.D )
  );
  al_aoi21ttf _119_ (
    .a(\DFF_19.Q ),
    .b(_001_),
    .c(_060_),
    .y(_003_)
  );
  al_ao21 _120_ (
    .a(\DFF_11.Q ),
    .b(\DFF_3.Q ),
    .c(\DFF_2.Q ),
    .y(_004_)
  );
  al_aoi21ftf _121_ (
    .a(\DFF_13.Q ),
    .b(\DFF_3.Q ),
    .c(_004_),
    .y(_005_)
  );
  al_and2 _122_ (
    .a(_005_),
    .b(_003_),
    .y(\DFF_13.D )
  );
  al_nand3ftt _123_ (
    .a(\DFF_3.Q ),
    .b(\DFF_10.Q ),
    .c(\DFF_11.Q ),
    .y(_006_)
  );
  al_aoi21ftf _124_ (
    .a(\DFF_14.Q ),
    .b(_004_),
    .c(_006_),
    .y(_007_)
  );
  al_aoi21ftt _125_ (
    .a(_036_),
    .b(_000_),
    .c(_058_),
    .y(_008_)
  );
  al_and3 _126_ (
    .a(_007_),
    .b(_008_),
    .c(_003_),
    .y(\DFF_14.D )
  );
  al_nand2ft _127_ (
    .a(\DFF_15.Q ),
    .b(_004_),
    .y(_009_)
  );
  al_and3 _128_ (
    .a(_008_),
    .b(_009_),
    .c(_003_),
    .y(\DFF_15.D )
  );
  al_nand2 _129_ (
    .a(\DFF_16.Q ),
    .b(_004_),
    .y(_010_)
  );
  al_nand3 _130_ (
    .a(_008_),
    .b(_010_),
    .c(_003_),
    .y(_011_)
  );
  al_aoi21ftf _131_ (
    .a(_051_),
    .b(_002_),
    .c(_011_),
    .y(\DFF_16.D )
  );
  al_oai21ttf _132_ (
    .a(\DFF_11.Q ),
    .b(\DFF_2.Q ),
    .c(\DFF_17.Q ),
    .y(_012_)
  );
  al_and3fft _133_ (
    .a(\DFF_11.Q ),
    .b(\DFF_2.Q ),
    .c(\DFF_10.Q ),
    .y(_013_)
  );
  al_nor3fft _134_ (
    .a(\DFF_3.Q ),
    .b(_012_),
    .c(_013_),
    .y(_014_)
  );
  al_mux2l _135_ (
    .a(_051_),
    .b(_014_),
    .s(_002_),
    .y(\DFF_17.D )
  );
  al_mux2l _136_ (
    .a(\DFF_18.Q ),
    .b(\DFF_10.Q ),
    .s(\DFF_3.Q ),
    .y(_015_)
  );
  al_and3ftt _137_ (
    .a(_058_),
    .b(_032_),
    .c(_015_),
    .y(_016_)
  );
  al_and2 _138_ (
    .a(_016_),
    .b(_003_),
    .y(\DFF_18.D )
  );
  al_oa21ttf _139_ (
    .a(\DFF_19.Q ),
    .b(G2),
    .c(G0),
    .y(_017_)
  );
  al_aoi21ttf _140_ (
    .a(\DFF_19.Q ),
    .b(G2),
    .c(_017_),
    .y(\DFF_19.D )
  );
  al_oa21ttf _141_ (
    .a(\DFF_20.Q ),
    .b(G1),
    .c(G0),
    .y(_018_)
  );
  al_aoi21ttf _142_ (
    .a(\DFF_20.Q ),
    .b(G1),
    .c(_018_),
    .y(\DFF_20.D )
  );
  al_dffl _143_ (
    .clk(CK),
    .d(\DFF_0.D ),
    .q(\DFF_0.Q )
  );
  al_dffl _144_ (
    .clk(CK),
    .d(\DFF_1.D ),
    .q(\DFF_1.Q )
  );
  al_dffl _145_ (
    .clk(CK),
    .d(\DFF_2.D ),
    .q(\DFF_2.Q )
  );
  al_dffl _146_ (
    .clk(CK),
    .d(\DFF_3.D ),
    .q(\DFF_3.Q )
  );
  al_dffl _147_ (
    .clk(CK),
    .d(\DFF_4.D ),
    .q(\DFF_4.Q )
  );
  al_dffl _148_ (
    .clk(CK),
    .d(\DFF_5.D ),
    .q(\DFF_5.Q )
  );
  al_dffl _149_ (
    .clk(CK),
    .d(\DFF_6.D ),
    .q(\DFF_6.Q )
  );
  al_dffl _150_ (
    .clk(CK),
    .d(\DFF_7.D ),
    .q(\DFF_7.Q )
  );
  al_dffl _151_ (
    .clk(CK),
    .d(\DFF_8.D ),
    .q(\DFF_8.Q )
  );
  al_dffl _152_ (
    .clk(CK),
    .d(\DFF_9.D ),
    .q(\DFF_9.Q )
  );
  al_dffl _153_ (
    .clk(CK),
    .d(\DFF_10.D ),
    .q(\DFF_10.Q )
  );
  al_dffl _154_ (
    .clk(CK),
    .d(\DFF_11.D ),
    .q(\DFF_11.Q )
  );
  al_dffl _155_ (
    .clk(CK),
    .d(\DFF_12.D ),
    .q(\DFF_12.Q )
  );
  al_dffl _156_ (
    .clk(CK),
    .d(\DFF_13.D ),
    .q(\DFF_13.Q )
  );
  al_dffl _157_ (
    .clk(CK),
    .d(\DFF_14.D ),
    .q(\DFF_14.Q )
  );
  al_dffl _158_ (
    .clk(CK),
    .d(\DFF_15.D ),
    .q(\DFF_15.Q )
  );
  al_dffl _159_ (
    .clk(CK),
    .d(\DFF_16.D ),
    .q(\DFF_16.Q )
  );
  al_dffl _160_ (
    .clk(CK),
    .d(\DFF_17.D ),
    .q(\DFF_17.Q )
  );
  al_dffl _161_ (
    .clk(CK),
    .d(\DFF_18.D ),
    .q(\DFF_18.Q )
  );
  al_dffl _162_ (
    .clk(CK),
    .d(\DFF_19.D ),
    .q(\DFF_19.Q )
  );
  al_dffl _163_ (
    .clk(CK),
    .d(\DFF_20.D ),
    .q(\DFF_20.Q )
  );
  assign \DFF_0.CK  = CK;
  assign \DFF_1.CK  = CK;
  assign \DFF_10.CK  = CK;
  assign \DFF_11.CK  = CK;
  assign \DFF_12.CK  = CK;
  assign \DFF_13.CK  = CK;
  assign \DFF_14.CK  = CK;
  assign \DFF_15.CK  = CK;
  assign \DFF_16.CK  = CK;
  assign \DFF_17.CK  = CK;
  assign \DFF_18.CK  = CK;
  assign \DFF_19.CK  = CK;
  assign \DFF_2.CK  = CK;
  assign \DFF_20.CK  = CK;
  assign \DFF_3.CK  = CK;
  assign \DFF_4.CK  = CK;
  assign \DFF_5.CK  = CK;
  assign \DFF_6.CK  = CK;
  assign \DFF_7.CK  = CK;
  assign \DFF_8.CK  = CK;
  assign \DFF_9.CK  = CK;
  assign G10 = \DFF_0.Q ;
  assign G101 = \DFF_8.D ;
  assign G106 = \DFF_9.D ;
  assign G11 = \DFF_1.Q ;
  assign G115 = \DFF_10.D ;
  assign G12 = \DFF_2.Q ;
  assign G126 = G0;
  assign G127 = \DFF_11.D ;
  assign G13 = \DFF_3.Q ;
  assign G137 = \DFF_12.D ;
  assign G14 = \DFF_4.Q ;
  assign G147 = \DFF_13.Q ;
  assign G148 = \DFF_14.Q ;
  assign G15 = \DFF_5.Q ;
  assign G16 = \DFF_6.Q ;
  assign G167 = \DFF_13.D ;
  assign G17 = \DFF_7.Q ;
  assign G173 = \DFF_14.D ;
  assign G179 = \DFF_15.D ;
  assign G18 = \DFF_8.Q ;
  assign G183 = \DFF_16.D ;
  assign G188 = \DFF_17.D ;
  assign G19 = \DFF_9.Q ;
  assign G194 = \DFF_18.D ;
  assign G198 = \DFF_15.Q ;
  assign G199 = \DFF_16.Q ;
  assign G20 = \DFF_10.Q ;
  assign G200 = \DFF_19.D ;
  assign G205 = G2;
  assign G206 = \DFF_20.D ;
  assign G21 = \DFF_11.Q ;
  assign G211 = G0;
  assign G212 = G1;
  assign G213 = \DFF_17.Q ;
  assign G214 = \DFF_18.Q ;
  assign G22 = \DFF_12.Q ;
  assign G23 = \DFF_13.Q ;
  assign G24 = \DFF_14.Q ;
  assign G25 = \DFF_15.Q ;
  assign G26 = \DFF_16.Q ;
  assign G27 = \DFF_17.Q ;
  assign G28 = \DFF_18.Q ;
  assign G29 = \DFF_19.Q ;
  assign G30 = \DFF_20.Q ;
  assign G60 = \DFF_0.D ;
  assign G61 = \DFF_1.D ;
  assign G62 = \DFF_2.D ;
  assign G69 = \DFF_3.D ;
  assign G79 = \DFF_4.D ;
  assign G84 = \DFF_5.D ;
  assign G89 = \DFF_6.D ;
  assign G96 = \DFF_7.D ;
endmodule
