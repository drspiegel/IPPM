
module s641(GND, VDD, CK, G1, G10, G100BF, G101BF, G103BF, G104BF, G105BF, G106BF, G107, G11, G12, G13, G138, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G4, G5, G6, G8, G83, G84, G85, G86BF, G87BF, G88BF, G89BF, G9, G90, G91, G92, G94, G95BF, G96BF, G97BF, G98BF, G99BF);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  input CK;
  wire \DFF_0.CK ;
  wire \DFF_0.D ;
  wire \DFF_0.Q ;
  wire \DFF_1.CK ;
  wire \DFF_1.D ;
  wire \DFF_1.Q ;
  wire \DFF_10.CK ;
  wire \DFF_10.D ;
  wire \DFF_10.Q ;
  wire \DFF_11.CK ;
  wire \DFF_11.D ;
  wire \DFF_11.Q ;
  wire \DFF_12.CK ;
  wire \DFF_12.D ;
  wire \DFF_12.Q ;
  wire \DFF_13.CK ;
  wire \DFF_13.D ;
  wire \DFF_13.Q ;
  wire \DFF_14.CK ;
  wire \DFF_14.D ;
  wire \DFF_14.Q ;
  wire \DFF_15.CK ;
  wire \DFF_15.D ;
  wire \DFF_15.Q ;
  wire \DFF_16.CK ;
  wire \DFF_16.D ;
  wire \DFF_16.Q ;
  wire \DFF_17.CK ;
  wire \DFF_17.D ;
  wire \DFF_17.Q ;
  wire \DFF_18.CK ;
  wire \DFF_18.D ;
  wire \DFF_18.Q ;
  wire \DFF_2.CK ;
  wire \DFF_2.D ;
  wire \DFF_2.Q ;
  wire \DFF_3.CK ;
  wire \DFF_3.D ;
  wire \DFF_3.Q ;
  wire \DFF_4.CK ;
  wire \DFF_4.D ;
  wire \DFF_4.Q ;
  wire \DFF_5.CK ;
  wire \DFF_5.D ;
  wire \DFF_5.Q ;
  wire \DFF_6.CK ;
  wire \DFF_6.D ;
  wire \DFF_6.Q ;
  wire \DFF_7.CK ;
  wire \DFF_7.D ;
  wire \DFF_7.Q ;
  wire \DFF_8.CK ;
  wire \DFF_8.D ;
  wire \DFF_8.Q ;
  wire \DFF_9.CK ;
  wire \DFF_9.D ;
  wire \DFF_9.Q ;
  input G1;
  input G10;
  output G100BF;
  output G101BF;
  output G103BF;
  output G104BF;
  output G105BF;
  output G106BF;
  output G107;
  wire G109;
  input G11;
  wire G111;
  wire G113;
  wire G115;
  wire G117;
  wire G119;
  input G12;
  wire G121;
  wire G122;
  wire G125;
  wire G126;
  wire G127;
  wire G128;
  wire G129;
  input G13;
  wire G130;
  wire G131;
  wire G132;
  wire G133;
  output G138;
  wire G139;
  input G14;
  wire G140;
  wire G141;
  wire G142;
  wire G146;
  input G15;
  wire G150;
  wire G158;
  input G16;
  input G17;
  input G18;
  input G19;
  input G2;
  input G20;
  wire G209;
  input G21;
  wire G211;
  wire G213;
  wire G215;
  wire G217;
  wire G219;
  input G22;
  wire G221;
  wire G223;
  wire G229;
  input G23;
  input G24;
  input G25;
  wire G250;
  input G26;
  wire G262;
  input G27;
  wire G271;
  wire G272;
  wire G273;
  wire G274;
  wire G275;
  wire G276;
  wire G277;
  wire G278;
  input G28;
  input G29;
  wire G293;
  wire G294;
  input G3;
  input G30;
  wire G300;
  wire G301;
  wire G306;
  wire G307;
  input G31;
  input G32;
  input G33;
  input G34;
  input G35;
  wire G352;
  wire G354;
  wire G356;
  wire G358;
  wire G359;
  input G36;
  wire G360;
  wire G361;
  wire G362;
  wire G363;
  wire G364;
  wire G367;
  wire G380;
  wire G383;
  wire G386;
  wire G388;
  wire G389;
  wire G394;
  input G4;
  input G5;
  input G6;
  wire G64;
  wire G65;
  wire G66;
  wire G67;
  wire G68;
  wire G69;
  wire G70;
  wire G71;
  wire G72;
  wire G73;
  wire G74;
  wire G75;
  wire G76;
  wire G77;
  wire G78;
  wire G79;
  input G8;
  wire G80;
  wire G81;
  wire G82;
  output G83;
  output G84;
  output G85;
  output G86BF;
  output G87BF;
  output G88BF;
  output G89BF;
  input G9;
  output G90;
  output G91;
  output G92;
  output G94;
  output G95BF;
  output G96BF;
  output G97BF;
  output G98BF;
  output G99BF;
  input GND;
  wire II335;
  wire II338;
  wire II341;
  wire II373;
  wire II440;
  wire II449;
  wire II452;
  wire II511;
  wire II524;
  wire II527;
  wire IIII208;
  wire IIII285;
  wire IIII320;
  wire IIII327;
  wire IIII334;
  wire IIII341;
  wire IIII348;
  wire IIII398;
  wire IIII406;
  wire IIII414;
  wire IIII422;
  wire IIII476;
  input VDD;
  al_nand3ftt _056_ (
    .a(G4),
    .b(\DFF_5.Q ),
    .c(G35),
    .y(G100BF)
  );
  al_nand3ftt _057_ (
    .a(G4),
    .b(\DFF_7.Q ),
    .c(G33),
    .y(G98BF)
  );
  al_nand3ftt _058_ (
    .a(G4),
    .b(\DFF_9.Q ),
    .c(G31),
    .y(G96BF)
  );
  al_and2ft _059_ (
    .a(G13),
    .b(G10),
    .y(_050_)
  );
  al_nand3ftt _060_ (
    .a(G3),
    .b(G9),
    .c(_050_),
    .y(_051_)
  );
  al_or2 _061_ (
    .a(G3),
    .b(G11),
    .y(_052_)
  );
  al_and3ftt _062_ (
    .a(\DFF_18.Q ),
    .b(G25),
    .c(_052_),
    .y(_053_)
  );
  al_nand2 _063_ (
    .a(_051_),
    .b(_053_),
    .y(G89BF)
  );
  al_nand3fft _064_ (
    .a(G3),
    .b(G9),
    .c(_050_),
    .y(_054_)
  );
  al_and2ft _065_ (
    .a(\DFF_16.Q ),
    .b(G23),
    .y(_055_)
  );
  al_nand3 _066_ (
    .a(_052_),
    .b(_055_),
    .c(_054_),
    .y(G87BF)
  );
  al_and3 _067_ (
    .a(\DFF_4.Q ),
    .b(_051_),
    .c(_053_),
    .y(\DFF_4.D )
  );
  al_nand2 _068_ (
    .a(G36),
    .b(\DFF_4.D ),
    .y(G101BF)
  );
  al_ao21 _069_ (
    .a(_051_),
    .b(_053_),
    .c(G3),
    .y(_000_)
  );
  al_nand3 _070_ (
    .a(\DFF_14.Q ),
    .b(G17),
    .c(_000_),
    .y(G106BF)
  );
  al_or3fft _071_ (
    .a(\DFF_8.Q ),
    .b(G32),
    .c(G87BF),
    .y(G97BF)
  );
  al_inv _072_ (
    .a(G3),
    .y(_001_)
  );
  al_inv _073_ (
    .a(\DFF_12.Q ),
    .y(_002_)
  );
  al_aoi21 _074_ (
    .a(_001_),
    .b(G87BF),
    .c(_002_),
    .y(_003_)
  );
  al_nand2 _075_ (
    .a(G15),
    .b(_003_),
    .y(G104BF)
  );
  al_and2ft _076_ (
    .a(G4),
    .b(\DFF_7.Q ),
    .y(_004_)
  );
  al_oai21ftt _077_ (
    .a(\DFF_8.Q ),
    .b(G87BF),
    .c(_004_),
    .y(\DFF_8.D )
  );
  al_mux2l _078_ (
    .a(_004_),
    .b(\DFF_8.Q ),
    .s(G87BF),
    .y(\DFF_7.D )
  );
  al_and2ft _079_ (
    .a(G2),
    .b(\DFF_2.Q ),
    .y(_005_)
  );
  al_ao21ttf _080_ (
    .a(\DFF_14.Q ),
    .b(_000_),
    .c(_005_),
    .y(_006_)
  );
  al_nor2 _081_ (
    .a(G10),
    .b(G13),
    .y(_007_)
  );
  al_nand3ftt _082_ (
    .a(G3),
    .b(G9),
    .c(_007_),
    .y(_008_)
  );
  al_and3 _083_ (
    .a(G24),
    .b(_052_),
    .c(_008_),
    .y(_009_)
  );
  al_nand2 _084_ (
    .a(_009_),
    .b(_006_),
    .y(G88BF)
  );
  al_aoi21ttf _085_ (
    .a(_001_),
    .b(G88BF),
    .c(\DFF_13.Q ),
    .y(\DFF_2.D )
  );
  al_or3fft _086_ (
    .a(\DFF_6.Q ),
    .b(G34),
    .c(G88BF),
    .y(G99BF)
  );
  al_ao21 _087_ (
    .a(_009_),
    .b(_006_),
    .c(G3),
    .y(_010_)
  );
  al_nand3 _088_ (
    .a(\DFF_13.Q ),
    .b(G16),
    .c(_010_),
    .y(G105BF)
  );
  al_and2ft _089_ (
    .a(G4),
    .b(\DFF_5.Q ),
    .y(_011_)
  );
  al_nand3 _090_ (
    .a(\DFF_6.Q ),
    .b(_009_),
    .c(_006_),
    .y(_012_)
  );
  al_nand2 _091_ (
    .a(_011_),
    .b(_012_),
    .y(\DFF_6.D )
  );
  al_ao21ttf _092_ (
    .a(_011_),
    .b(G88BF),
    .c(_012_),
    .y(\DFF_5.D )
  );
  al_inv _093_ (
    .a(_003_),
    .y(_013_)
  );
  al_and2 _094_ (
    .a(\DFF_14.Q ),
    .b(_000_),
    .y(_014_)
  );
  al_aoi21 _095_ (
    .a(\DFF_13.Q ),
    .b(_010_),
    .c(_014_),
    .y(_015_)
  );
  al_and2ft _096_ (
    .a(G2),
    .b(\DFF_0.Q ),
    .y(_016_)
  );
  al_nand3 _097_ (
    .a(_013_),
    .b(_016_),
    .c(_015_),
    .y(_017_)
  );
  al_nand3fft _098_ (
    .a(G3),
    .b(G9),
    .c(_007_),
    .y(_018_)
  );
  al_and3 _099_ (
    .a(G22),
    .b(_052_),
    .c(_018_),
    .y(_019_)
  );
  al_nand2 _100_ (
    .a(_019_),
    .b(_017_),
    .y(G86BF)
  );
  al_inv _101_ (
    .a(\DFF_11.Q ),
    .y(_020_)
  );
  al_aoi21 _102_ (
    .a(_001_),
    .b(G86BF),
    .c(_020_),
    .y(\DFF_0.D )
  );
  al_and3 _103_ (
    .a(\DFF_10.Q ),
    .b(_019_),
    .c(_017_),
    .y(_021_)
  );
  al_nand2 _104_ (
    .a(G30),
    .b(_021_),
    .y(G95BF)
  );
  al_ao21 _105_ (
    .a(_019_),
    .b(_017_),
    .c(G3),
    .y(_022_)
  );
  al_nand3 _106_ (
    .a(\DFF_11.Q ),
    .b(G14),
    .c(_022_),
    .y(G103BF)
  );
  al_or3ftt _107_ (
    .a(\DFF_9.Q ),
    .b(G4),
    .c(_021_),
    .y(\DFF_10.D )
  );
  al_and2ft _108_ (
    .a(G4),
    .b(\DFF_9.Q ),
    .y(_023_)
  );
  al_ao21 _109_ (
    .a(_023_),
    .b(G86BF),
    .c(_021_),
    .y(\DFF_9.D )
  );
  al_and3ftt _110_ (
    .a(G4),
    .b(\DFF_15.Q ),
    .c(G18),
    .y(G107)
  );
  al_and3ftt _111_ (
    .a(G4),
    .b(\DFF_16.Q ),
    .c(G19),
    .y(G83)
  );
  al_and3ftt _112_ (
    .a(G4),
    .b(\DFF_17.Q ),
    .c(G20),
    .y(G84)
  );
  al_and3ftt _113_ (
    .a(G4),
    .b(\DFF_18.Q ),
    .c(G21),
    .y(G85)
  );
  al_and2 _114_ (
    .a(G11),
    .b(G12),
    .y(_024_)
  );
  al_and3 _115_ (
    .a(G13),
    .b(G28),
    .c(_024_),
    .y(G92)
  );
  al_inv _116_ (
    .a(G2),
    .y(_025_)
  );
  al_and3 _117_ (
    .a(_025_),
    .b(\DFF_14.Q ),
    .c(_000_),
    .y(\DFF_18.D )
  );
  al_inv _118_ (
    .a(_014_),
    .y(_026_)
  );
  al_and3 _119_ (
    .a(_025_),
    .b(_026_),
    .c(\DFF_2.D ),
    .y(\DFF_17.D )
  );
  al_and3 _120_ (
    .a(_025_),
    .b(_003_),
    .c(_015_),
    .y(\DFF_16.D )
  );
  al_and3fft _121_ (
    .a(_003_),
    .b(\DFF_2.D ),
    .c(_026_),
    .y(_027_)
  );
  al_and3 _122_ (
    .a(_025_),
    .b(_027_),
    .c(\DFF_0.D ),
    .y(\DFF_15.D )
  );
  al_nor3fft _123_ (
    .a(\DFF_6.Q ),
    .b(_011_),
    .c(G88BF),
    .y(_028_)
  );
  al_nand2 _124_ (
    .a(G9),
    .b(_007_),
    .y(_029_)
  );
  al_nor3fft _125_ (
    .a(\DFF_8.Q ),
    .b(_004_),
    .c(G87BF),
    .y(_030_)
  );
  al_and3ftt _126_ (
    .a(G11),
    .b(\DFF_4.D ),
    .c(_030_),
    .y(_031_)
  );
  al_nand3 _127_ (
    .a(_023_),
    .b(_031_),
    .c(_021_),
    .y(_032_)
  );
  al_nand2 _128_ (
    .a(_029_),
    .b(_032_),
    .y(_033_)
  );
  al_and2ft _129_ (
    .a(G9),
    .b(_007_),
    .y(_034_)
  );
  al_nand3 _130_ (
    .a(_023_),
    .b(_034_),
    .c(_021_),
    .y(_035_)
  );
  al_oa21ftt _131_ (
    .a(G9),
    .b(\DFF_4.D ),
    .c(_050_),
    .y(_036_)
  );
  al_oai21 _132_ (
    .a(G9),
    .b(_030_),
    .c(_036_),
    .y(_037_)
  );
  al_and3 _133_ (
    .a(G12),
    .b(G26),
    .c(_037_),
    .y(_038_)
  );
  al_nand2 _134_ (
    .a(_038_),
    .b(_035_),
    .y(_039_)
  );
  al_aoi21 _135_ (
    .a(_028_),
    .b(_033_),
    .c(_039_),
    .y(G90)
  );
  al_nand3 _136_ (
    .a(_023_),
    .b(_027_),
    .c(_021_),
    .y(_040_)
  );
  al_nand3fft _137_ (
    .a(G2),
    .b(_020_),
    .c(_022_),
    .y(_041_)
  );
  al_nand2ft _138_ (
    .a(G8),
    .b(_041_),
    .y(_042_)
  );
  al_aoi21ftf _139_ (
    .a(\DFF_0.D ),
    .b(_040_),
    .c(_042_),
    .y(\DFF_11.D )
  );
  al_and3 _140_ (
    .a(G5),
    .b(_030_),
    .c(_015_),
    .y(_043_)
  );
  al_aoi21ftf _141_ (
    .a(G5),
    .b(G2),
    .c(_003_),
    .y(_044_)
  );
  al_oai21ftf _142_ (
    .a(_043_),
    .b(\DFF_0.D ),
    .c(_044_),
    .y(\DFF_12.D )
  );
  al_aoi21 _143_ (
    .a(\DFF_11.Q ),
    .b(_022_),
    .c(_003_),
    .y(_045_)
  );
  al_and3 _144_ (
    .a(G6),
    .b(_026_),
    .c(_028_),
    .y(_046_)
  );
  al_aoi21ftf _145_ (
    .a(G6),
    .b(G2),
    .c(\DFF_2.D ),
    .y(_047_)
  );
  al_ao21 _146_ (
    .a(_046_),
    .b(_045_),
    .c(_047_),
    .y(\DFF_13.D )
  );
  al_nor3fft _147_ (
    .a(G1),
    .b(\DFF_4.D ),
    .c(\DFF_2.D ),
    .y(_048_)
  );
  al_aoi21ftf _148_ (
    .a(G1),
    .b(G2),
    .c(_014_),
    .y(_049_)
  );
  al_ao21 _149_ (
    .a(_048_),
    .b(_045_),
    .c(_049_),
    .y(\DFF_14.D )
  );
  al_dffl _150_ (
    .clk(CK),
    .d(\DFF_0.D ),
    .q(\DFF_0.Q )
  );
  al_dffl _151_ (
    .clk(CK),
    .d(\DFF_2.D ),
    .q(\DFF_2.Q )
  );
  al_dffl _152_ (
    .clk(CK),
    .d(\DFF_4.D ),
    .q(\DFF_4.Q )
  );
  al_dffl _153_ (
    .clk(CK),
    .d(\DFF_5.D ),
    .q(\DFF_5.Q )
  );
  al_dffl _154_ (
    .clk(CK),
    .d(\DFF_6.D ),
    .q(\DFF_6.Q )
  );
  al_dffl _155_ (
    .clk(CK),
    .d(\DFF_7.D ),
    .q(\DFF_7.Q )
  );
  al_dffl _156_ (
    .clk(CK),
    .d(\DFF_8.D ),
    .q(\DFF_8.Q )
  );
  al_dffl _157_ (
    .clk(CK),
    .d(\DFF_9.D ),
    .q(\DFF_9.Q )
  );
  al_dffl _158_ (
    .clk(CK),
    .d(\DFF_10.D ),
    .q(\DFF_10.Q )
  );
  al_dffl _159_ (
    .clk(CK),
    .d(\DFF_11.D ),
    .q(\DFF_11.Q )
  );
  al_dffl _160_ (
    .clk(CK),
    .d(\DFF_12.D ),
    .q(\DFF_12.Q )
  );
  al_dffl _161_ (
    .clk(CK),
    .d(\DFF_13.D ),
    .q(\DFF_13.Q )
  );
  al_dffl _162_ (
    .clk(CK),
    .d(\DFF_14.D ),
    .q(\DFF_14.Q )
  );
  al_dffl _163_ (
    .clk(CK),
    .d(\DFF_15.D ),
    .q(\DFF_15.Q )
  );
  al_dffl _164_ (
    .clk(CK),
    .d(\DFF_16.D ),
    .q(\DFF_16.Q )
  );
  al_dffl _165_ (
    .clk(CK),
    .d(\DFF_17.D ),
    .q(\DFF_17.Q )
  );
  al_dffl _166_ (
    .clk(CK),
    .d(\DFF_18.D ),
    .q(\DFF_18.Q )
  );
  assign \DFF_0.CK  = CK;
  assign \DFF_1.CK  = CK;
  assign \DFF_1.D  = \DFF_16.D ;
  assign \DFF_1.Q  = \DFF_16.Q ;
  assign \DFF_10.CK  = CK;
  assign \DFF_11.CK  = CK;
  assign \DFF_12.CK  = CK;
  assign \DFF_13.CK  = CK;
  assign \DFF_14.CK  = CK;
  assign \DFF_15.CK  = CK;
  assign \DFF_16.CK  = CK;
  assign \DFF_17.CK  = CK;
  assign \DFF_18.CK  = CK;
  assign \DFF_2.CK  = CK;
  assign \DFF_3.CK  = CK;
  assign \DFF_3.D  = \DFF_18.D ;
  assign \DFF_3.Q  = \DFF_18.Q ;
  assign \DFF_4.CK  = CK;
  assign \DFF_5.CK  = CK;
  assign \DFF_6.CK  = CK;
  assign \DFF_7.CK  = CK;
  assign \DFF_8.CK  = CK;
  assign \DFF_9.CK  = CK;
  assign G109 = \DFF_4.Q ;
  assign G111 = \DFF_5.Q ;
  assign G113 = \DFF_6.Q ;
  assign G115 = \DFF_7.Q ;
  assign G117 = \DFF_8.Q ;
  assign G119 = \DFF_9.Q ;
  assign G121 = \DFF_10.Q ;
  assign G122 = \DFF_4.D ;
  assign G125 = \DFF_11.D ;
  assign G126 = \DFF_12.D ;
  assign G127 = \DFF_13.D ;
  assign G128 = \DFF_14.D ;
  assign G129 = \DFF_15.D ;
  assign G130 = \DFF_16.D ;
  assign G131 = \DFF_17.D ;
  assign G132 = \DFF_18.D ;
  assign G133 = \DFF_5.D ;
  assign G138 = \DFF_6.D ;
  assign G139 = \DFF_7.D ;
  assign G140 = \DFF_8.D ;
  assign G141 = \DFF_9.D ;
  assign G142 = \DFF_10.D ;
  assign G146 = \DFF_4.D ;
  assign G150 = \DFF_0.D ;
  assign G158 = \DFF_2.D ;
  assign G209 = \DFF_11.Q ;
  assign G211 = \DFF_12.Q ;
  assign G213 = \DFF_13.Q ;
  assign G215 = \DFF_14.Q ;
  assign G217 = \DFF_15.Q ;
  assign G219 = \DFF_16.Q ;
  assign G221 = \DFF_17.Q ;
  assign G223 = \DFF_18.Q ;
  assign G229 = \DFF_18.D ;
  assign G250 = \DFF_18.D ;
  assign G262 = \DFF_16.D ;
  assign G271 = \DFF_11.D ;
  assign G272 = \DFF_12.D ;
  assign G273 = \DFF_13.D ;
  assign G274 = \DFF_14.D ;
  assign G275 = \DFF_15.D ;
  assign G276 = \DFF_16.D ;
  assign G277 = \DFF_17.D ;
  assign G278 = \DFF_18.D ;
  assign G293 = \DFF_4.D ;
  assign G294 = \DFF_4.D ;
  assign G300 = \DFF_0.D ;
  assign G301 = \DFF_0.D ;
  assign G306 = \DFF_2.D ;
  assign G307 = \DFF_2.D ;
  assign G352 = G1;
  assign G354 = G86BF;
  assign G356 = G87BF;
  assign G358 = G88BF;
  assign G359 = G89BF;
  assign G360 = G4;
  assign G361 = G5;
  assign G362 = G6;
  assign G363 = G8;
  assign G364 = G9;
  assign G367 = G10;
  assign G380 = \DFF_0.D ;
  assign G383 = \DFF_4.D ;
  assign G386 = G11;
  assign G388 = G12;
  assign G389 = G13;
  assign G394 = \DFF_2.D ;
  assign G64 = \DFF_0.Q ;
  assign G65 = \DFF_16.Q ;
  assign G66 = \DFF_2.Q ;
  assign G67 = \DFF_18.Q ;
  assign G68 = \DFF_4.Q ;
  assign G69 = \DFF_5.Q ;
  assign G70 = \DFF_6.Q ;
  assign G71 = \DFF_7.Q ;
  assign G72 = \DFF_8.Q ;
  assign G73 = \DFF_9.Q ;
  assign G74 = \DFF_10.Q ;
  assign G75 = \DFF_11.Q ;
  assign G76 = \DFF_12.Q ;
  assign G77 = \DFF_13.Q ;
  assign G78 = \DFF_14.Q ;
  assign G79 = \DFF_15.Q ;
  assign G80 = \DFF_16.Q ;
  assign G81 = \DFF_17.Q ;
  assign G82 = \DFF_18.Q ;
  assign G91 = G27;
  assign G94 = G29;
  assign II335 = G87BF;
  assign II338 = G89BF;
  assign II341 = G87BF;
  assign II373 = \DFF_8.D ;
  assign II440 = \DFF_6.D ;
  assign II449 = G88BF;
  assign II452 = G88BF;
  assign II511 = \DFF_10.D ;
  assign II524 = G86BF;
  assign II527 = G86BF;
  assign IIII208 = \DFF_4.D ;
  assign IIII285 = \DFF_5.D ;
  assign IIII320 = \DFF_6.D ;
  assign IIII327 = \DFF_7.D ;
  assign IIII334 = \DFF_8.D ;
  assign IIII341 = \DFF_9.D ;
  assign IIII348 = \DFF_10.D ;
  assign IIII398 = G86BF;
  assign IIII406 = G87BF;
  assign IIII414 = G88BF;
  assign IIII422 = G89BF;
  assign IIII476 = \DFF_4.D ;
endmodule
