
module s953(GND, VDD, CK, ActBmHS1, ActRtHS1, DumpIIHS1, FullIIHS1, FullOHS1, GoBmHS1, GoRtHS1, IInDoneHS1, LdProgHS1, LoadIIHHS1, LoadOHHS1, LxHIInHS1, Mode0HS1, Mode1HS1, Mode2HS1, NewLineHS1, NewTrHS1, OutAvHS1, OutputHS1, Prog_0, Prog_1, Prog_2, Rdy1BmHS1, Rdy1RtHS1, Rdy2BmHS1, Rdy2RtHS1, ReRtTSHS1, ReWhBufHS1, RtTSHS1, SeFullIIHS1, SeFullOHS1, SeOutAvHS1, ShftIIRHS1, ShftORHS1, TgWhBufHS1, TpArrayHS1, TxHIInHS1, WantBmHS1, WantRtHS1);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  output ActBmHS1;
  output ActRtHS1;
  input CK;
  wire \DFF_0.CK ;
  wire \DFF_0.D ;
  wire \DFF_0.Q ;
  wire \DFF_1.CK ;
  wire \DFF_1.D ;
  wire \DFF_1.Q ;
  wire \DFF_10.CK ;
  wire \DFF_10.D ;
  wire \DFF_10.Q ;
  wire \DFF_11.CK ;
  wire \DFF_11.D ;
  wire \DFF_11.Q ;
  wire \DFF_12.CK ;
  wire \DFF_12.D ;
  wire \DFF_12.Q ;
  wire \DFF_13.CK ;
  wire \DFF_13.D ;
  wire \DFF_13.Q ;
  wire \DFF_14.CK ;
  wire \DFF_14.D ;
  wire \DFF_14.Q ;
  wire \DFF_15.CK ;
  wire \DFF_15.D ;
  wire \DFF_15.Q ;
  wire \DFF_16.CK ;
  wire \DFF_16.D ;
  wire \DFF_16.Q ;
  wire \DFF_17.CK ;
  wire \DFF_17.D ;
  wire \DFF_17.Q ;
  wire \DFF_18.CK ;
  wire \DFF_18.D ;
  wire \DFF_18.Q ;
  wire \DFF_19.CK ;
  wire \DFF_19.D ;
  wire \DFF_19.Q ;
  wire \DFF_2.CK ;
  wire \DFF_2.D ;
  wire \DFF_2.Q ;
  wire \DFF_20.CK ;
  wire \DFF_20.D ;
  wire \DFF_20.Q ;
  wire \DFF_21.CK ;
  wire \DFF_21.D ;
  wire \DFF_21.Q ;
  wire \DFF_22.CK ;
  wire \DFF_22.D ;
  wire \DFF_22.Q ;
  wire \DFF_23.CK ;
  wire \DFF_23.D ;
  wire \DFF_23.Q ;
  wire \DFF_24.CK ;
  wire \DFF_24.D ;
  wire \DFF_24.Q ;
  wire \DFF_25.CK ;
  wire \DFF_25.D ;
  wire \DFF_25.Q ;
  wire \DFF_26.CK ;
  wire \DFF_26.D ;
  wire \DFF_26.Q ;
  wire \DFF_27.CK ;
  wire \DFF_27.D ;
  wire \DFF_27.Q ;
  wire \DFF_28.CK ;
  wire \DFF_28.D ;
  wire \DFF_28.Q ;
  wire \DFF_3.CK ;
  wire \DFF_3.D ;
  wire \DFF_3.Q ;
  wire \DFF_4.CK ;
  wire \DFF_4.D ;
  wire \DFF_4.Q ;
  wire \DFF_5.CK ;
  wire \DFF_5.D ;
  wire \DFF_5.Q ;
  wire \DFF_6.CK ;
  wire \DFF_6.D ;
  wire \DFF_6.Q ;
  wire \DFF_7.CK ;
  wire \DFF_7.D ;
  wire \DFF_7.Q ;
  wire \DFF_8.CK ;
  wire \DFF_8.D ;
  wire \DFF_8.Q ;
  wire \DFF_9.CK ;
  wire \DFF_9.D ;
  wire \DFF_9.Q ;
  output DumpIIHS1;
  input FullIIHS1;
  input FullOHS1;
  input GND;
  output GoBmHS1;
  output GoRtHS1;
  wire II10;
  wire II11;
  wire II12;
  wire II13;
  wire II14;
  wire II15;
  wire II16;
  wire II17;
  wire II18;
  wire II19;
  wire II2;
  wire II20;
  wire II21;
  wire II22;
  wire II23;
  wire II24;
  wire II25;
  wire II26;
  wire II27;
  wire II28;
  wire II29;
  wire II3;
  wire II30;
  wire II322;
  wire II4;
  wire II414;
  wire II5;
  wire II6;
  wire II7;
  wire II8;
  wire II9;
  input IInDoneHS1;
  output LdProgHS1;
  output LoadIIHHS1;
  output LoadOHHS1;
  output LxHIInHS1;
  output Mode0HS1;
  output Mode1HS1;
  output Mode2HS1;
  output NewLineHS1;
  output NewTrHS1;
  input OutAvHS1;
  input OutputHS1;
  input Prog_0;
  input Prog_1;
  input Prog_2;
  input Rdy1BmHS1;
  input Rdy1RtHS1;
  input Rdy2BmHS1;
  input Rdy2RtHS1;
  output ReRtTSHS1;
  output ReWhBufHS1;
  input RtTSHS1;
  output SeFullIIHS1;
  output SeFullOHS1;
  output SeOutAvHS1;
  output ShftIIRHS1;
  output ShftORHS1;
  wire State_0;
  wire State_1;
  wire State_2;
  wire State_3;
  wire State_4;
  wire State_5;
  output TgWhBufHS1;
  input TpArrayHS1;
  output TxHIInHS1;
  input VDD;
  input WantBmHS1;
  input WantRtHS1;
  al_and3fft _199_ (
    .a(Prog_2),
    .b(\DFF_1.Q ),
    .c(Prog_0),
    .y(_156_)
  );
  al_nand3fft _200_ (
    .a(\DFF_3.Q ),
    .b(\DFF_2.Q ),
    .c(\DFF_0.Q ),
    .y(_157_)
  );
  al_and2ft _201_ (
    .a(\DFF_4.Q ),
    .b(\DFF_5.Q ),
    .y(_158_)
  );
  al_and3ftt _202_ (
    .a(_157_),
    .b(_156_),
    .c(_158_),
    .y(_159_)
  );
  al_or2 _203_ (
    .a(\DFF_5.Q ),
    .b(\DFF_4.Q ),
    .y(_160_)
  );
  al_nor3ftt _204_ (
    .a(\DFF_1.Q ),
    .b(_157_),
    .c(_160_),
    .y(\DFF_14.D )
  );
  al_inv _205_ (
    .a(\DFF_3.Q ),
    .y(_161_)
  );
  al_and2ft _206_ (
    .a(\DFF_2.Q ),
    .b(\DFF_0.Q ),
    .y(_162_)
  );
  al_and3ftt _207_ (
    .a(\DFF_5.Q ),
    .b(\DFF_4.Q ),
    .c(_162_),
    .y(_163_)
  );
  al_ao21ftf _208_ (
    .a(_156_),
    .b(_161_),
    .c(_163_),
    .y(_164_)
  );
  al_nand3fft _209_ (
    .a(_159_),
    .b(\DFF_14.D ),
    .c(_164_),
    .y(\DFF_6.D )
  );
  al_nand2 _210_ (
    .a(Prog_0),
    .b(\DFF_14.D ),
    .y(_165_)
  );
  al_and2ft _211_ (
    .a(\DFF_1.Q ),
    .b(\DFF_3.Q ),
    .y(_166_)
  );
  al_or3 _212_ (
    .a(Prog_0),
    .b(Prog_2),
    .c(\DFF_1.Q ),
    .y(_167_)
  );
  al_ao21ftf _213_ (
    .a(_166_),
    .b(_167_),
    .c(_163_),
    .y(_168_)
  );
  al_nand3ftt _214_ (
    .a(_159_),
    .b(_168_),
    .c(_165_),
    .y(\DFF_12.D )
  );
  al_nor2 _215_ (
    .a(\DFF_1.Q ),
    .b(\DFF_0.Q ),
    .y(_169_)
  );
  al_and3fft _216_ (
    .a(\DFF_1.Q ),
    .b(\DFF_0.Q ),
    .c(\DFF_2.Q ),
    .y(_170_)
  );
  al_nand3ftt _217_ (
    .a(\DFF_3.Q ),
    .b(\DFF_5.Q ),
    .c(_170_),
    .y(_171_)
  );
  al_aoi21ftf _218_ (
    .a(_160_),
    .b(_169_),
    .c(_171_),
    .y(_172_)
  );
  al_and3fft _219_ (
    .a(\DFF_3.Q ),
    .b(\DFF_2.Q ),
    .c(\DFF_0.Q ),
    .y(_173_)
  );
  al_and2ft _220_ (
    .a(\DFF_1.Q ),
    .b(_173_),
    .y(_174_)
  );
  al_nand3ftt _221_ (
    .a(Rdy1BmHS1),
    .b(\DFF_5.Q ),
    .c(_174_),
    .y(_175_)
  );
  al_nand2 _222_ (
    .a(Rdy2RtHS1),
    .b(Prog_0),
    .y(_176_)
  );
  al_or2 _223_ (
    .a(Rdy1BmHS1),
    .b(Prog_0),
    .y(_177_)
  );
  al_ao21 _224_ (
    .a(_177_),
    .b(_176_),
    .c(FullIIHS1),
    .y(_178_)
  );
  al_nand2ft _225_ (
    .a(Prog_0),
    .b(Rdy2BmHS1),
    .y(_179_)
  );
  al_nand2ft _226_ (
    .a(Rdy1RtHS1),
    .b(Prog_0),
    .y(_180_)
  );
  al_ao21 _227_ (
    .a(_179_),
    .b(_180_),
    .c(FullOHS1),
    .y(_181_)
  );
  al_nand3fft _228_ (
    .a(Prog_2),
    .b(\DFF_5.Q ),
    .c(_173_),
    .y(_182_)
  );
  al_ao21 _229_ (
    .a(_181_),
    .b(_178_),
    .c(_182_),
    .y(_183_)
  );
  al_nand3 _230_ (
    .a(_172_),
    .b(_175_),
    .c(_183_),
    .y(\DFF_19.D )
  );
  al_nand3fft _231_ (
    .a(Rdy1BmHS1),
    .b(Rdy1RtHS1),
    .c(_174_),
    .y(_184_)
  );
  al_or2 _232_ (
    .a(Prog_2),
    .b(\DFF_5.Q ),
    .y(_185_)
  );
  al_oai21ttf _233_ (
    .a(FullIIHS1),
    .b(FullOHS1),
    .c(\DFF_1.Q ),
    .y(_186_)
  );
  al_or3fft _234_ (
    .a(_185_),
    .b(_173_),
    .c(_186_),
    .y(_187_)
  );
  al_nand3ftt _235_ (
    .a(\DFF_4.Q ),
    .b(\DFF_5.Q ),
    .c(_162_),
    .y(_188_)
  );
  al_and2 _236_ (
    .a(Rdy1BmHS1),
    .b(Rdy2BmHS1),
    .y(_189_)
  );
  al_nand3fft _237_ (
    .a(Prog_0),
    .b(\DFF_4.Q ),
    .c(_173_),
    .y(_190_)
  );
  al_ao21 _238_ (
    .a(_190_),
    .b(_188_),
    .c(_189_),
    .y(_191_)
  );
  al_nand3 _239_ (
    .a(_187_),
    .b(_184_),
    .c(_191_),
    .y(_192_)
  );
  al_nand2 _240_ (
    .a(Rdy1RtHS1),
    .b(Rdy2RtHS1),
    .y(_193_)
  );
  al_nand3ftt _241_ (
    .a(\DFF_5.Q ),
    .b(Prog_0),
    .c(_173_),
    .y(_194_)
  );
  al_oa21ftt _242_ (
    .a(_194_),
    .b(_163_),
    .c(_193_),
    .y(_195_)
  );
  al_and3ftt _243_ (
    .a(\DFF_5.Q ),
    .b(\DFF_3.Q ),
    .c(_169_),
    .y(_196_)
  );
  al_and3fft _244_ (
    .a(\DFF_4.Q ),
    .b(\DFF_2.Q ),
    .c(RtTSHS1),
    .y(_197_)
  );
  al_and2 _245_ (
    .a(_197_),
    .b(_196_),
    .y(\DFF_11.D )
  );
  al_oai21 _246_ (
    .a(Prog_1),
    .b(Prog_2),
    .c(\DFF_11.D ),
    .y(_198_)
  );
  al_or3fft _247_ (
    .a(\DFF_1.Q ),
    .b(_173_),
    .c(_160_),
    .y(_000_)
  );
  al_and2ft _248_ (
    .a(\DFF_4.Q ),
    .b(_173_),
    .y(_001_)
  );
  al_and2ft _249_ (
    .a(\DFF_5.Q ),
    .b(Prog_2),
    .y(_002_)
  );
  al_aoi21ttf _250_ (
    .a(_002_),
    .b(_001_),
    .c(_000_),
    .y(_003_)
  );
  al_nor2 _251_ (
    .a(Prog_2),
    .b(\DFF_1.Q ),
    .y(_004_)
  );
  al_nand2ft _252_ (
    .a(\DFF_2.Q ),
    .b(\DFF_0.Q ),
    .y(_005_)
  );
  al_and2 _253_ (
    .a(\DFF_5.Q ),
    .b(\DFF_4.Q ),
    .y(_006_)
  );
  al_and3fft _254_ (
    .a(_005_),
    .b(_006_),
    .c(_160_),
    .y(_007_)
  );
  al_ao21ftf _255_ (
    .a(_004_),
    .b(_161_),
    .c(_007_),
    .y(_008_)
  );
  al_and3 _256_ (
    .a(_003_),
    .b(_008_),
    .c(_198_),
    .y(_009_)
  );
  al_nand3fft _257_ (
    .a(_192_),
    .b(_195_),
    .c(_009_),
    .y(\DFF_0.D )
  );
  al_and3ftt _258_ (
    .a(_005_),
    .b(_004_),
    .c(_158_),
    .y(_010_)
  );
  al_or2 _259_ (
    .a(Prog_2),
    .b(\DFF_1.Q ),
    .y(_011_)
  );
  al_and2ft _260_ (
    .a(\DFF_5.Q ),
    .b(\DFF_4.Q ),
    .y(_012_)
  );
  al_nand3fft _261_ (
    .a(_157_),
    .b(_011_),
    .c(_012_),
    .y(_013_)
  );
  al_oai21ftf _262_ (
    .a(_013_),
    .b(_010_),
    .c(Prog_0),
    .y(_014_)
  );
  al_and2ft _263_ (
    .a(\DFF_3.Q ),
    .b(_170_),
    .y(_015_)
  );
  al_and3ftt _264_ (
    .a(\DFF_5.Q ),
    .b(\DFF_3.Q ),
    .c(_170_),
    .y(_016_)
  );
  al_ao21ftt _265_ (
    .a(_012_),
    .b(_015_),
    .c(_016_),
    .y(\DFF_10.D )
  );
  al_oa21ftt _266_ (
    .a(\DFF_3.Q ),
    .b(_188_),
    .c(_000_),
    .y(_017_)
  );
  al_nand3ftt _267_ (
    .a(\DFF_10.D ),
    .b(_017_),
    .c(_014_),
    .y(\DFF_7.D )
  );
  al_nor2 _268_ (
    .a(\DFF_4.Q ),
    .b(\DFF_3.Q ),
    .y(_018_)
  );
  al_nand3fft _269_ (
    .a(\DFF_1.Q ),
    .b(\DFF_0.Q ),
    .c(_018_),
    .y(_019_)
  );
  al_or2 _270_ (
    .a(FullIIHS1),
    .b(FullOHS1),
    .y(_020_)
  );
  al_nand3fft _271_ (
    .a(\DFF_5.Q ),
    .b(_020_),
    .c(_189_),
    .y(_021_)
  );
  al_or3 _272_ (
    .a(\DFF_2.Q ),
    .b(_019_),
    .c(_021_),
    .y(_022_)
  );
  al_nand3ftt _273_ (
    .a(\DFF_4.Q ),
    .b(\DFF_5.Q ),
    .c(_173_),
    .y(_023_)
  );
  al_and2ft _274_ (
    .a(Rdy2BmHS1),
    .b(Rdy1BmHS1),
    .y(_024_)
  );
  al_oai21 _275_ (
    .a(Prog_2),
    .b(\DFF_1.Q ),
    .c(_186_),
    .y(_025_)
  );
  al_or3ftt _276_ (
    .a(_024_),
    .b(_023_),
    .c(_025_),
    .y(_026_)
  );
  al_and3fft _277_ (
    .a(FullIIHS1),
    .b(\DFF_1.Q ),
    .c(_173_),
    .y(_027_)
  );
  al_or3 _278_ (
    .a(Rdy1BmHS1),
    .b(Rdy1RtHS1),
    .c(FullOHS1),
    .y(_028_)
  );
  al_and3ftt _279_ (
    .a(_028_),
    .b(_006_),
    .c(_027_),
    .y(_029_)
  );
  al_nor3fft _280_ (
    .a(_026_),
    .b(_022_),
    .c(_029_),
    .y(_030_)
  );
  al_nand2 _281_ (
    .a(FullIIHS1),
    .b(FullOHS1),
    .y(_031_)
  );
  al_inv _282_ (
    .a(Prog_0),
    .y(_032_)
  );
  al_or3 _283_ (
    .a(Prog_2),
    .b(\DFF_5.Q ),
    .c(\DFF_1.Q ),
    .y(_033_)
  );
  al_and3ftt _284_ (
    .a(_033_),
    .b(_032_),
    .c(_001_),
    .y(_034_)
  );
  al_nor2 _285_ (
    .a(Rdy1BmHS1),
    .b(Rdy2BmHS1),
    .y(_035_)
  );
  al_nor2 _286_ (
    .a(_035_),
    .b(_189_),
    .y(_036_)
  );
  al_nand3 _287_ (
    .a(_031_),
    .b(_036_),
    .c(_034_),
    .y(_037_)
  );
  al_nand3ftt _288_ (
    .a(\DFF_4.Q ),
    .b(Prog_2),
    .c(_173_),
    .y(_038_)
  );
  al_oa21ftt _289_ (
    .a(Rdy1RtHS1),
    .b(Rdy2RtHS1),
    .c(WantRtHS1),
    .y(_039_)
  );
  al_or3 _290_ (
    .a(FullIIHS1),
    .b(FullOHS1),
    .c(\DFF_1.Q ),
    .y(_040_)
  );
  al_and3fft _291_ (
    .a(Rdy2BmHS1),
    .b(_040_),
    .c(Rdy1BmHS1),
    .y(_041_)
  );
  al_nand3fft _292_ (
    .a(_039_),
    .b(_038_),
    .c(_041_),
    .y(_042_)
  );
  al_or2ft _293_ (
    .a(WantBmHS1),
    .b(_042_),
    .y(_043_)
  );
  al_nand3 _294_ (
    .a(_037_),
    .b(_043_),
    .c(_030_),
    .y(\DFF_9.D )
  );
  al_nand3fft _295_ (
    .a(Rdy2BmHS1),
    .b(_005_),
    .c(_158_),
    .y(_044_)
  );
  al_aoi21ftf _296_ (
    .a(Rdy2RtHS1),
    .b(_163_),
    .c(_044_),
    .y(_045_)
  );
  al_ao21ftf _297_ (
    .a(_161_),
    .b(_007_),
    .c(_045_),
    .y(_046_)
  );
  al_nor2 _298_ (
    .a(Prog_0),
    .b(Prog_1),
    .y(_047_)
  );
  al_nand2 _299_ (
    .a(Prog_0),
    .b(Prog_1),
    .y(_048_)
  );
  al_nor3fft _300_ (
    .a(Rdy2BmHS1),
    .b(_048_),
    .c(_047_),
    .y(_049_)
  );
  al_oa21ftt _301_ (
    .a(Rdy1BmHS1),
    .b(Rdy2BmHS1),
    .c(WantBmHS1),
    .y(_050_)
  );
  al_ao21 _302_ (
    .a(_176_),
    .b(_039_),
    .c(_050_),
    .y(_051_)
  );
  al_ao21ftf _303_ (
    .a(_039_),
    .b(_049_),
    .c(_051_),
    .y(_052_)
  );
  al_and3ftt _304_ (
    .a(_040_),
    .b(_002_),
    .c(_001_),
    .y(_053_)
  );
  al_and2ft _305_ (
    .a(IInDoneHS1),
    .b(\DFF_14.D ),
    .y(_054_)
  );
  al_aoi21 _306_ (
    .a(_053_),
    .b(_052_),
    .c(_054_),
    .y(_055_)
  );
  al_ao21ttf _307_ (
    .a(\DFF_1.Q ),
    .b(_046_),
    .c(_055_),
    .y(\DFF_1.D )
  );
  al_and3 _308_ (
    .a(Rdy1RtHS1),
    .b(_173_),
    .c(_002_),
    .y(_056_)
  );
  al_nand3fft _309_ (
    .a(Rdy2RtHS1),
    .b(_040_),
    .c(_056_),
    .y(_057_)
  );
  al_nand3fft _310_ (
    .a(\DFF_4.Q ),
    .b(_157_),
    .c(_002_),
    .y(_058_)
  );
  al_or3 _311_ (
    .a(WantRtHS1),
    .b(_040_),
    .c(_058_),
    .y(_059_)
  );
  al_aoi21 _312_ (
    .a(_059_),
    .b(_057_),
    .c(WantBmHS1),
    .y(_060_)
  );
  al_nor2 _313_ (
    .a(Rdy1RtHS1),
    .b(Rdy2RtHS1),
    .y(_061_)
  );
  al_nand2ft _314_ (
    .a(_061_),
    .b(_193_),
    .y(_062_)
  );
  al_inv _315_ (
    .a(FullOHS1),
    .y(_063_)
  );
  al_and3ftt _316_ (
    .a(_033_),
    .b(_063_),
    .c(_001_),
    .y(_064_)
  );
  al_nand3fft _317_ (
    .a(_032_),
    .b(_062_),
    .c(_064_),
    .y(_065_)
  );
  al_nand3fft _318_ (
    .a(\DFF_5.Q ),
    .b(\DFF_4.Q ),
    .c(\DFF_3.Q ),
    .y(_066_)
  );
  al_nand3ftt _319_ (
    .a(\DFF_3.Q ),
    .b(TpArrayHS1),
    .c(_006_),
    .y(_067_)
  );
  al_ao21ttf _320_ (
    .a(_066_),
    .b(_067_),
    .c(_170_),
    .y(_068_)
  );
  al_nand3ftt _321_ (
    .a(_029_),
    .b(_068_),
    .c(_065_),
    .y(_069_)
  );
  al_nand3 _322_ (
    .a(_063_),
    .b(_036_),
    .c(_034_),
    .y(_070_)
  );
  al_and2ft _323_ (
    .a(Rdy2RtHS1),
    .b(Rdy1RtHS1),
    .y(_071_)
  );
  al_nand3ftt _324_ (
    .a(Rdy2BmHS1),
    .b(Rdy1BmHS1),
    .c(_158_),
    .y(_072_)
  );
  al_ao21ttf _325_ (
    .a(_012_),
    .b(_071_),
    .c(_072_),
    .y(_073_)
  );
  al_and2ft _326_ (
    .a(FullOHS1),
    .b(Prog_2),
    .y(_074_)
  );
  al_and3 _327_ (
    .a(_027_),
    .b(_074_),
    .c(_073_),
    .y(_075_)
  );
  al_nor3fft _328_ (
    .a(_042_),
    .b(_070_),
    .c(_075_),
    .y(_076_)
  );
  al_nand3fft _329_ (
    .a(_060_),
    .b(_069_),
    .c(_076_),
    .y(\DFF_20.D )
  );
  al_and3 _330_ (
    .a(Rdy2RtHS1),
    .b(WantRtHS1),
    .c(_053_),
    .y(_077_)
  );
  al_or2 _331_ (
    .a(WantBmHS1),
    .b(Prog_0),
    .y(_078_)
  );
  al_nand2ft _332_ (
    .a(_047_),
    .b(_048_),
    .y(_079_)
  );
  al_nand2 _333_ (
    .a(Rdy2BmHS1),
    .b(WantBmHS1),
    .y(_080_)
  );
  al_and3fft _334_ (
    .a(_080_),
    .b(_059_),
    .c(_079_),
    .y(_081_)
  );
  al_ao21ftt _335_ (
    .a(_078_),
    .b(_077_),
    .c(_081_),
    .y(\DFF_28.D )
  );
  al_or3 _336_ (
    .a(\DFF_4.Q ),
    .b(_157_),
    .c(_033_),
    .y(_082_)
  );
  al_mux2l _337_ (
    .a(_024_),
    .b(_071_),
    .s(_032_),
    .y(_083_)
  );
  al_and2ft _338_ (
    .a(FullIIHS1),
    .b(FullOHS1),
    .y(_084_)
  );
  al_nand3ftt _339_ (
    .a(_082_),
    .b(_084_),
    .c(_083_),
    .y(_085_)
  );
  al_nand3fft _340_ (
    .a(_157_),
    .b(_186_),
    .c(_006_),
    .y(_086_)
  );
  al_nand3ftt _341_ (
    .a(IInDoneHS1),
    .b(\DFF_4.Q ),
    .c(_016_),
    .y(_087_)
  );
  al_nand3 _342_ (
    .a(_086_),
    .b(_087_),
    .c(_085_),
    .y(_088_)
  );
  al_and3fft _343_ (
    .a(FullIIHS1),
    .b(FullOHS1),
    .c(Prog_2),
    .y(_089_)
  );
  al_nand2ft _344_ (
    .a(Prog_2),
    .b(IInDoneHS1),
    .y(_090_)
  );
  al_nand3fft _345_ (
    .a(\DFF_1.Q ),
    .b(_089_),
    .c(_090_),
    .y(_091_)
  );
  al_ao21ttf _346_ (
    .a(Rdy1RtHS1),
    .b(Rdy2RtHS1),
    .c(_011_),
    .y(_092_)
  );
  al_nand3 _347_ (
    .a(_161_),
    .b(_092_),
    .c(_091_),
    .y(_093_)
  );
  al_nand2 _348_ (
    .a(_163_),
    .b(_093_),
    .y(_094_)
  );
  al_and3ftt _349_ (
    .a(\DFF_2.Q ),
    .b(_012_),
    .c(_166_),
    .y(_095_)
  );
  al_aoi21ttf _350_ (
    .a(_193_),
    .b(_095_),
    .c(_171_),
    .y(_096_)
  );
  al_and2ft _351_ (
    .a(Rdy1BmHS1),
    .b(Rdy2BmHS1),
    .y(_097_)
  );
  al_or3ftt _352_ (
    .a(_097_),
    .b(_023_),
    .c(_025_),
    .y(_098_)
  );
  al_nand3 _353_ (
    .a(_096_),
    .b(_098_),
    .c(_094_),
    .y(_099_)
  );
  al_nand3fft _354_ (
    .a(\DFF_4.Q ),
    .b(_040_),
    .c(_056_),
    .y(_100_)
  );
  al_ao21ftf _355_ (
    .a(Rdy2RtHS1),
    .b(WantRtHS1),
    .c(_053_),
    .y(_101_)
  );
  al_ao21 _356_ (
    .a(_100_),
    .b(_101_),
    .c(_080_),
    .y(_102_)
  );
  al_nand3fft _357_ (
    .a(_088_),
    .b(_099_),
    .c(_102_),
    .y(\DFF_4.D )
  );
  al_nand2 _358_ (
    .a(OutputHS1),
    .b(\DFF_14.D ),
    .y(_103_)
  );
  al_aoi21 _359_ (
    .a(_166_),
    .b(_007_),
    .c(_010_),
    .y(_104_)
  );
  al_ao21ttf _360_ (
    .a(_103_),
    .b(_104_),
    .c(IInDoneHS1),
    .y(_105_)
  );
  al_and3fft _361_ (
    .a(_033_),
    .b(_190_),
    .c(_097_),
    .y(_106_)
  );
  al_aoi21ftt _362_ (
    .a(FullOHS1),
    .b(_106_),
    .c(_029_),
    .y(_107_)
  );
  al_and3fft _363_ (
    .a(FullOHS1),
    .b(_082_),
    .c(Prog_0),
    .y(_108_)
  );
  al_and2ft _364_ (
    .a(Rdy1RtHS1),
    .b(Rdy2RtHS1),
    .y(_109_)
  );
  al_aoi21ttf _365_ (
    .a(_109_),
    .b(_108_),
    .c(_068_),
    .y(_110_)
  );
  al_nand3 _366_ (
    .a(_107_),
    .b(_110_),
    .c(_105_),
    .y(\DFF_23.D )
  );
  al_nor2 _367_ (
    .a(FullIIHS1),
    .b(OutAvHS1),
    .y(\DFF_26.D )
  );
  al_and2ft _368_ (
    .a(OutAvHS1),
    .b(FullIIHS1),
    .y(\DFF_25.D )
  );
  al_oa21ttf _369_ (
    .a(FullIIHS1),
    .b(FullOHS1),
    .c(OutAvHS1),
    .y(\DFF_22.D )
  );
  al_and3fft _370_ (
    .a(\DFF_3.Q ),
    .b(_160_),
    .c(_170_),
    .y(\DFF_27.D )
  );
  al_nand3ftt _371_ (
    .a(\DFF_5.Q ),
    .b(\DFF_4.Q ),
    .c(_173_),
    .y(_111_)
  );
  al_oai21ftt _372_ (
    .a(_004_),
    .b(_111_),
    .c(_000_),
    .y(\DFF_17.D )
  );
  al_ao21ftf _373_ (
    .a(_166_),
    .b(_011_),
    .c(_007_),
    .y(_112_)
  );
  al_ao21ftf _374_ (
    .a(_000_),
    .b(Prog_1),
    .c(_112_),
    .y(\DFF_13.D )
  );
  al_nand3ftt _375_ (
    .a(TpArrayHS1),
    .b(\DFF_5.Q ),
    .c(_015_),
    .y(_113_)
  );
  al_inv _376_ (
    .a(\DFF_2.Q ),
    .y(_114_)
  );
  al_ao21 _377_ (
    .a(_114_),
    .b(_021_),
    .c(_019_),
    .y(_115_)
  );
  al_nand2 _378_ (
    .a(\DFF_4.Q ),
    .b(_016_),
    .y(_116_)
  );
  al_aoi21ttf _379_ (
    .a(_158_),
    .b(_170_),
    .c(_116_),
    .y(_117_)
  );
  al_nand3 _380_ (
    .a(_113_),
    .b(_115_),
    .c(_117_),
    .y(\DFF_2.D )
  );
  al_nand3ftt _381_ (
    .a(\DFF_3.Q ),
    .b(_170_),
    .c(_006_),
    .y(_118_)
  );
  al_ao21ftf _382_ (
    .a(_197_),
    .b(_196_),
    .c(_118_),
    .y(_119_)
  );
  al_and3ftt _383_ (
    .a(IInDoneHS1),
    .b(\DFF_3.Q ),
    .c(_007_),
    .y(_120_)
  );
  al_or3ftt _384_ (
    .a(_071_),
    .b(_111_),
    .c(_025_),
    .y(_121_)
  );
  al_and3 _385_ (
    .a(_026_),
    .b(_022_),
    .c(_121_),
    .y(_122_)
  );
  al_nand3fft _386_ (
    .a(_119_),
    .b(_120_),
    .c(_122_),
    .y(\DFF_3.D )
  );
  al_aoi21ftf _387_ (
    .a(_012_),
    .b(_015_),
    .c(_000_),
    .y(_123_)
  );
  al_nand3 _388_ (
    .a(_116_),
    .b(_123_),
    .c(_104_),
    .y(\DFF_16.D )
  );
  al_nand3 _389_ (
    .a(_032_),
    .b(_031_),
    .c(_001_),
    .y(_124_)
  );
  al_ao21 _390_ (
    .a(_038_),
    .b(_124_),
    .c(Rdy2BmHS1),
    .y(_125_)
  );
  al_aoi21ttf _391_ (
    .a(FullIIHS1),
    .b(FullOHS1),
    .c(Prog_0),
    .y(_126_)
  );
  al_nand3fft _392_ (
    .a(Rdy2RtHS1),
    .b(\DFF_5.Q ),
    .c(_173_),
    .y(_127_)
  );
  al_oai21ttf _393_ (
    .a(Prog_2),
    .b(_126_),
    .c(_127_),
    .y(_128_)
  );
  al_nand3fft _394_ (
    .a(\DFF_2.Q ),
    .b(\DFF_1.Q ),
    .c(_002_),
    .y(_129_)
  );
  al_aoi21ftf _395_ (
    .a(_129_),
    .b(_018_),
    .c(_172_),
    .y(_130_)
  );
  al_nand3 _396_ (
    .a(_128_),
    .b(_130_),
    .c(_125_),
    .y(\DFF_18.D )
  );
  al_nand3 _397_ (
    .a(Prog_2),
    .b(_197_),
    .c(_196_),
    .y(_131_)
  );
  al_nor3fft _398_ (
    .a(_082_),
    .b(_131_),
    .c(_029_),
    .y(_132_)
  );
  al_nand3ftt _399_ (
    .a(_075_),
    .b(_022_),
    .c(_132_),
    .y(\DFF_15.D )
  );
  al_and3fft _400_ (
    .a(_040_),
    .b(_058_),
    .c(Rdy2RtHS1),
    .y(_133_)
  );
  al_nand3fft _401_ (
    .a(Rdy1BmHS1),
    .b(Rdy2BmHS1),
    .c(WantBmHS1),
    .y(_134_)
  );
  al_and3 _402_ (
    .a(WantRtHS1),
    .b(_134_),
    .c(_133_),
    .y(_135_)
  );
  al_ao21ttf _403_ (
    .a(Rdy1BmHS1),
    .b(Rdy2BmHS1),
    .c(_011_),
    .y(_136_)
  );
  al_nand3 _404_ (
    .a(_161_),
    .b(_136_),
    .c(_091_),
    .y(_137_)
  );
  al_and2ft _405_ (
    .a(_188_),
    .b(_137_),
    .y(_138_)
  );
  al_or3ftt _406_ (
    .a(_109_),
    .b(_111_),
    .c(_025_),
    .y(_139_)
  );
  al_aoi21ttf _407_ (
    .a(_083_),
    .b(_064_),
    .c(_139_),
    .y(_140_)
  );
  al_and3 _408_ (
    .a(_086_),
    .b(_115_),
    .c(_140_),
    .y(_141_)
  );
  al_nand3fft _409_ (
    .a(_135_),
    .b(_138_),
    .c(_141_),
    .y(\DFF_5.D )
  );
  al_and3fft _410_ (
    .a(_050_),
    .b(_057_),
    .c(WantRtHS1),
    .y(_142_)
  );
  al_nor3ftt _411_ (
    .a(_126_),
    .b(_082_),
    .c(_062_),
    .y(_143_)
  );
  al_nand2ft _412_ (
    .a(\DFF_2.Q ),
    .b(\DFF_4.Q ),
    .y(_144_)
  );
  al_nand3fft _413_ (
    .a(_144_),
    .b(_193_),
    .c(_196_),
    .y(_145_)
  );
  al_nor3ftt _414_ (
    .a(_145_),
    .b(_029_),
    .c(_143_),
    .y(_146_)
  );
  al_nand3ftt _415_ (
    .a(_142_),
    .b(_121_),
    .c(_146_),
    .y(\DFF_8.D )
  );
  al_mux2h _416_ (
    .a(_071_),
    .b(_036_),
    .s(_032_),
    .y(_147_)
  );
  al_and3ftt _417_ (
    .a(_082_),
    .b(_084_),
    .c(_147_),
    .y(_148_)
  );
  al_or3ftt _418_ (
    .a(FullOHS1),
    .b(Prog_2),
    .c(_180_),
    .y(_149_)
  );
  al_or3ftt _419_ (
    .a(WantRtHS1),
    .b(WantBmHS1),
    .c(Prog_0),
    .y(_150_)
  );
  al_ao21ftf _420_ (
    .a(_150_),
    .b(_074_),
    .c(_149_),
    .y(_151_)
  );
  al_and3fft _421_ (
    .a(\DFF_5.Q ),
    .b(\DFF_4.Q ),
    .c(Rdy2RtHS1),
    .y(_152_)
  );
  al_and3 _422_ (
    .a(_027_),
    .b(_152_),
    .c(_151_),
    .y(_153_)
  );
  al_or3 _423_ (
    .a(_153_),
    .b(_081_),
    .c(_148_),
    .y(\DFF_21.D )
  );
  al_and3fft _424_ (
    .a(_011_),
    .b(_111_),
    .c(IInDoneHS1),
    .y(_154_)
  );
  al_ao21 _425_ (
    .a(_084_),
    .b(_106_),
    .c(_154_),
    .y(_155_)
  );
  al_or3 _426_ (
    .a(_153_),
    .b(_155_),
    .c(_081_),
    .y(\DFF_24.D )
  );
  al_dffl _427_ (
    .clk(CK),
    .d(\DFF_0.D ),
    .q(\DFF_0.Q )
  );
  al_dffl _428_ (
    .clk(CK),
    .d(\DFF_1.D ),
    .q(\DFF_1.Q )
  );
  al_dffl _429_ (
    .clk(CK),
    .d(\DFF_2.D ),
    .q(\DFF_2.Q )
  );
  al_dffl _430_ (
    .clk(CK),
    .d(\DFF_3.D ),
    .q(\DFF_3.Q )
  );
  al_dffl _431_ (
    .clk(CK),
    .d(\DFF_4.D ),
    .q(\DFF_4.Q )
  );
  al_dffl _432_ (
    .clk(CK),
    .d(\DFF_5.D ),
    .q(\DFF_5.Q )
  );
  al_dffl _433_ (
    .clk(CK),
    .d(\DFF_6.D ),
    .q(\DFF_6.Q )
  );
  al_dffl _434_ (
    .clk(CK),
    .d(\DFF_7.D ),
    .q(\DFF_7.Q )
  );
  al_dffl _435_ (
    .clk(CK),
    .d(\DFF_8.D ),
    .q(\DFF_8.Q )
  );
  al_dffl _436_ (
    .clk(CK),
    .d(\DFF_9.D ),
    .q(\DFF_9.Q )
  );
  al_dffl _437_ (
    .clk(CK),
    .d(\DFF_10.D ),
    .q(\DFF_10.Q )
  );
  al_dffl _438_ (
    .clk(CK),
    .d(\DFF_11.D ),
    .q(\DFF_11.Q )
  );
  al_dffl _439_ (
    .clk(CK),
    .d(\DFF_12.D ),
    .q(\DFF_12.Q )
  );
  al_dffl _440_ (
    .clk(CK),
    .d(\DFF_13.D ),
    .q(\DFF_13.Q )
  );
  al_dffl _441_ (
    .clk(CK),
    .d(\DFF_14.D ),
    .q(\DFF_14.Q )
  );
  al_dffl _442_ (
    .clk(CK),
    .d(\DFF_15.D ),
    .q(\DFF_15.Q )
  );
  al_dffl _443_ (
    .clk(CK),
    .d(\DFF_16.D ),
    .q(\DFF_16.Q )
  );
  al_dffl _444_ (
    .clk(CK),
    .d(\DFF_17.D ),
    .q(\DFF_17.Q )
  );
  al_dffl _445_ (
    .clk(CK),
    .d(\DFF_18.D ),
    .q(\DFF_18.Q )
  );
  al_dffl _446_ (
    .clk(CK),
    .d(\DFF_19.D ),
    .q(\DFF_19.Q )
  );
  al_dffl _447_ (
    .clk(CK),
    .d(\DFF_20.D ),
    .q(\DFF_20.Q )
  );
  al_dffl _448_ (
    .clk(CK),
    .d(\DFF_21.D ),
    .q(\DFF_21.Q )
  );
  al_dffl _449_ (
    .clk(CK),
    .d(\DFF_22.D ),
    .q(\DFF_22.Q )
  );
  al_dffl _450_ (
    .clk(CK),
    .d(\DFF_23.D ),
    .q(\DFF_23.Q )
  );
  al_dffl _451_ (
    .clk(CK),
    .d(\DFF_24.D ),
    .q(\DFF_24.Q )
  );
  al_dffl _452_ (
    .clk(CK),
    .d(\DFF_25.D ),
    .q(\DFF_25.Q )
  );
  al_dffl _453_ (
    .clk(CK),
    .d(\DFF_26.D ),
    .q(\DFF_26.Q )
  );
  al_dffl _454_ (
    .clk(CK),
    .d(\DFF_27.D ),
    .q(\DFF_27.Q )
  );
  al_dffl _455_ (
    .clk(CK),
    .d(\DFF_28.D ),
    .q(\DFF_28.Q )
  );
  assign ActBmHS1 = \DFF_7.Q ;
  assign ActRtHS1 = \DFF_6.Q ;
  assign \DFF_0.CK  = CK;
  assign \DFF_1.CK  = CK;
  assign \DFF_10.CK  = CK;
  assign \DFF_11.CK  = CK;
  assign \DFF_12.CK  = CK;
  assign \DFF_13.CK  = CK;
  assign \DFF_14.CK  = CK;
  assign \DFF_15.CK  = CK;
  assign \DFF_16.CK  = CK;
  assign \DFF_17.CK  = CK;
  assign \DFF_18.CK  = CK;
  assign \DFF_19.CK  = CK;
  assign \DFF_2.CK  = CK;
  assign \DFF_20.CK  = CK;
  assign \DFF_21.CK  = CK;
  assign \DFF_22.CK  = CK;
  assign \DFF_23.CK  = CK;
  assign \DFF_24.CK  = CK;
  assign \DFF_25.CK  = CK;
  assign \DFF_26.CK  = CK;
  assign \DFF_27.CK  = CK;
  assign \DFF_28.CK  = CK;
  assign \DFF_3.CK  = CK;
  assign \DFF_4.CK  = CK;
  assign \DFF_5.CK  = CK;
  assign \DFF_6.CK  = CK;
  assign \DFF_7.CK  = CK;
  assign \DFF_8.CK  = CK;
  assign \DFF_9.CK  = CK;
  assign DumpIIHS1 = \DFF_28.Q ;
  assign GoBmHS1 = \DFF_9.Q ;
  assign GoRtHS1 = \DFF_8.Q ;
  assign II10 = \DFF_8.D ;
  assign II11 = \DFF_9.D ;
  assign II12 = \DFF_10.D ;
  assign II13 = \DFF_11.D ;
  assign II14 = \DFF_12.D ;
  assign II15 = \DFF_13.D ;
  assign II16 = \DFF_14.D ;
  assign II17 = \DFF_15.D ;
  assign II18 = \DFF_16.D ;
  assign II19 = \DFF_17.D ;
  assign II2 = \DFF_0.D ;
  assign II20 = \DFF_18.D ;
  assign II21 = \DFF_19.D ;
  assign II22 = \DFF_20.D ;
  assign II23 = \DFF_21.D ;
  assign II24 = \DFF_22.D ;
  assign II25 = \DFF_23.D ;
  assign II26 = \DFF_24.D ;
  assign II27 = \DFF_25.D ;
  assign II28 = \DFF_26.D ;
  assign II29 = \DFF_27.D ;
  assign II3 = \DFF_1.D ;
  assign II30 = \DFF_28.D ;
  assign II322 = \DFF_14.D ;
  assign II4 = \DFF_2.D ;
  assign II414 = \DFF_11.D ;
  assign II5 = \DFF_3.D ;
  assign II6 = \DFF_4.D ;
  assign II7 = \DFF_5.D ;
  assign II8 = \DFF_6.D ;
  assign II9 = \DFF_7.D ;
  assign LdProgHS1 = \DFF_27.Q ;
  assign LoadIIHHS1 = \DFF_21.Q ;
  assign LoadOHHS1 = \DFF_20.Q ;
  assign LxHIInHS1 = \DFF_18.Q ;
  assign Mode0HS1 = \DFF_12.Q ;
  assign Mode1HS1 = \DFF_13.Q ;
  assign Mode2HS1 = \DFF_14.Q ;
  assign NewLineHS1 = \DFF_15.Q ;
  assign NewTrHS1 = \DFF_10.Q ;
  assign ReRtTSHS1 = \DFF_11.Q ;
  assign ReWhBufHS1 = \DFF_26.Q ;
  assign SeFullIIHS1 = \DFF_24.Q ;
  assign SeFullOHS1 = \DFF_23.Q ;
  assign SeOutAvHS1 = \DFF_22.Q ;
  assign ShftIIRHS1 = \DFF_17.Q ;
  assign ShftORHS1 = \DFF_16.Q ;
  assign State_0 = \DFF_5.Q ;
  assign State_1 = \DFF_4.Q ;
  assign State_2 = \DFF_3.Q ;
  assign State_3 = \DFF_2.Q ;
  assign State_4 = \DFF_1.Q ;
  assign State_5 = \DFF_0.Q ;
  assign TgWhBufHS1 = \DFF_25.Q ;
  assign TxHIInHS1 = \DFF_19.Q ;
endmodule
