
module c5315(N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, N106, N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N140, N141, N145, N146, N149, N152, N155, N158, N161, N164, N167, N170, N173, N176, N179, N182, N185, N188, N191, N194, N197, N200, N203, N206, N209, N210, N217, N218, N225, N226, N233, N234, N241, N242, N245, N248, N251, N254, N257, N264, N265, N272, N273, N280, N281, N288, N289, N292, N293, N299, N302, N307, N308, N315, N316, N323, N324, N331, N332, N335, N338, N341, N348, N351, N358, N361, N366, N369, N372, N373, N374, N386, N389, N400, N411, N422, N435, N446, N457, N468, N479, N490, N503, N514, N523, N534, N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, N610, N613, N616, N619, N625, N631, N709, N816, N1066, N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1147, N1152, N1153, N1154, N1155, N1972, N2054, N2060, N2061, N2139, N2142, N2309, N2387, N2527, N2584, N2590, N2623, N3357, N3358, N3359, N3360, N3604, N3613, N4272, N4275, N4278, N4279, N4737, N4738, N4739, N4740, N5240, N5388, N6641, N6643, N6646, N6648, N6716, N6877, N6924, N6925, N6926, N6927, N7015, N7363, N7365, N7432, N7449, N7465, N7466, N7467, N7469, N7470, N7471, N7472, N7473, N7474, N7476, N7503, N7504, N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520, N7521, N7522, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607, N7626, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706, N7707, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7754, N7755, N7756, N7757, N7758, N7759, N7760, N7761, N8075, N8076, N8123, N8124, N8127, N8128);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  input N1;
  input N100;
  input N103;
  input N106;
  output N1066;
  input N109;
  input N11;
  input N112;
  input N113;
  output N1137;
  output N1138;
  output N1139;
  input N114;
  output N1140;
  output N1141;
  output N1142;
  output N1143;
  output N1144;
  output N1145;
  output N1147;
  input N115;
  output N1152;
  output N1153;
  output N1154;
  output N1155;
  input N116;
  wire N1161;
  input N117;
  wire N1173;
  input N118;
  wire N1185;
  input N119;
  wire N1197;
  input N120;
  wire N1209;
  input N121;
  wire N1213;
  wire N1216;
  input N122;
  wire N1223;
  input N123;
  wire N1235;
  wire N1247;
  wire N1259;
  input N126;
  input N127;
  wire N1271;
  input N128;
  wire N1280;
  input N129;
  wire N1292;
  input N130;
  wire N1303;
  input N131;
  wire N1315;
  input N132;
  wire N1327;
  wire N1339;
  input N135;
  wire N1351;
  input N136;
  wire N1363;
  input N137;
  wire N1375;
  wire N1378;
  wire N1381;
  wire N1384;
  wire N1387;
  wire N1390;
  wire N1393;
  wire N1396;
  input N14;
  input N140;
  input N141;
  wire N1415;
  wire N1418;
  wire N1421;
  wire N1424;
  wire N1427;
  wire N1430;
  wire N1433;
  wire N1436;
  input N145;
  wire N1455;
  input N146;
  wire N1462;
  wire N1469;
  wire N1479;
  wire N1482;
  input N149;
  wire N1492;
  wire N1495;
  wire N1498;
  wire N1501;
  wire N1504;
  wire N1507;
  wire N1510;
  wire N1513;
  wire N1516;
  wire N1519;
  input N152;
  wire N1522;
  wire N1525;
  wire N1542;
  wire N1545;
  wire N1548;
  input N155;
  wire N1551;
  wire N1554;
  wire N1557;
  wire N1560;
  wire N1563;
  wire N1566;
  wire N1573;
  input N158;
  wire N1580;
  wire N1594;
  wire N1597;
  wire N1600;
  wire N1603;
  wire N1606;
  wire N1609;
  input N161;
  wire N1612;
  wire N1615;
  wire N1618;
  wire N1621;
  wire N1624;
  wire N1627;
  wire N1630;
  wire N1633;
  wire N1636;
  wire N1639;
  input N164;
  wire N1642;
  wire N1645;
  wire N1648;
  wire N1651;
  wire N1654;
  wire N1657;
  wire N1663;
  input N167;
  wire N1675;
  wire N1685;
  wire N1697;
  input N17;
  input N170;
  wire N1709;
  wire N1721;
  wire N1727;
  input N173;
  wire N1731;
  wire N1743;
  input N176;
  wire N1761;
  wire N1769;
  wire N1777;
  wire N1785;
  input N179;
  wire N1793;
  wire N1800;
  wire N1807;
  wire N1814;
  input N182;
  wire N1821;
  wire N1824;
  wire N1827;
  wire N1830;
  wire N1833;
  wire N1836;
  wire N1839;
  wire N1842;
  wire N1845;
  wire N1848;
  input N185;
  wire N1851;
  wire N1854;
  wire N1857;
  wire N1860;
  wire N1863;
  wire N1866;
  wire N1869;
  wire N1872;
  wire N1875;
  wire N1878;
  input N188;
  wire N1881;
  wire N1884;
  wire N1887;
  wire N1890;
  wire N1893;
  wire N1896;
  wire N1899;
  wire N1902;
  wire N1905;
  wire N1908;
  input N191;
  wire N1911;
  wire N1914;
  wire N1917;
  wire N1920;
  wire N1923;
  wire N1926;
  wire N1929;
  wire N1932;
  wire N1935;
  wire N1938;
  input N194;
  wire N1941;
  wire N1944;
  wire N1947;
  wire N1950;
  wire N1953;
  wire N1956;
  wire N1959;
  wire N1962;
  wire N1965;
  wire N1968;
  input N197;
  output N1972;
  input N20;
  input N200;
  input N203;
  output N2054;
  input N206;
  output N2060;
  output N2061;
  input N209;
  input N210;
  output N2139;
  output N2142;
  input N217;
  input N218;
  input N225;
  input N226;
  input N23;
  output N2309;
  input N233;
  input N234;
  output N2387;
  input N24;
  input N241;
  input N242;
  input N245;
  input N248;
  input N25;
  input N251;
  output N2527;
  input N254;
  input N257;
  output N2584;
  output N2590;
  input N26;
  output N2623;
  input N264;
  wire N2647;
  input N265;
  wire N2675;
  input N27;
  wire N2704;
  input N272;
  wire N2722;
  input N273;
  wire N2750;
  input N280;
  input N281;
  wire N2877;
  input N288;
  input N289;
  wire N2891;
  input N292;
  input N293;
  wire N2964;
  input N299;
  wire N3000;
  wire N3003;
  wire N3007;
  wire N3010;
  input N302;
  input N307;
  input N308;
  input N31;
  input N315;
  input N316;
  wire N3191;
  wire N3200;
  input N323;
  input N324;
  input N331;
  input N332;
  input N335;
  output N3357;
  output N3358;
  output N3359;
  output N3360;
  input N338;
  input N34;
  input N341;
  input N348;
  input N351;
  input N358;
  output N3604;
  input N361;
  output N3613;
  input N366;
  input N369;
  input N37;
  input N372;
  input N373;
  input N374;
  wire N3779;
  wire N3780;
  input N386;
  input N389;
  input N4;
  input N40;
  input N400;
  input N411;
  input N422;
  output N4272;
  output N4275;
  output N4278;
  output N4279;
  input N43;
  input N435;
  input N446;
  input N457;
  input N46;
  input N468;
  output N4737;
  output N4738;
  output N4739;
  output N4740;
  input N479;
  input N49;
  input N490;
  input N503;
  input N514;
  input N52;
  input N523;
  output N5240;
  input N53;
  input N534;
  output N5388;
  input N54;
  input N545;
  input N549;
  input N552;
  input N556;
  input N559;
  input N562;
  input N566;
  input N571;
  input N574;
  input N577;
  input N580;
  input N583;
  input N588;
  input N591;
  input N592;
  input N595;
  input N596;
  input N597;
  input N598;
  input N599;
  input N603;
  input N607;
  input N61;
  input N610;
  input N613;
  input N616;
  input N619;
  input N625;
  input N631;
  input N64;
  wire N6466;
  output N6641;
  output N6643;
  output N6646;
  output N6648;
  input N67;
  output N6716;
  wire N6724;
  output N6877;
  output N6924;
  output N6925;
  output N6926;
  output N6927;
  input N70;
  output N7015;
  output N709;
  input N73;
  output N7363;
  output N7365;
  wire N7394;
  wire N7397;
  wire N7431;
  output N7432;
  output N7449;
  output N7465;
  output N7466;
  output N7467;
  output N7469;
  output N7470;
  output N7471;
  output N7472;
  output N7473;
  output N7474;
  output N7476;
  output N7503;
  output N7504;
  output N7506;
  output N7511;
  output N7515;
  output N7516;
  output N7517;
  output N7518;
  output N7519;
  output N7520;
  output N7521;
  output N7522;
  input N76;
  output N7600;
  output N7601;
  output N7602;
  output N7603;
  output N7604;
  output N7605;
  output N7606;
  output N7607;
  output N7626;
  output N7698;
  output N7699;
  output N7700;
  output N7701;
  output N7702;
  output N7703;
  output N7704;
  output N7705;
  output N7706;
  output N7707;
  output N7735;
  output N7736;
  output N7737;
  output N7738;
  output N7739;
  output N7740;
  output N7741;
  output N7742;
  output N7754;
  output N7755;
  output N7756;
  output N7757;
  output N7758;
  output N7759;
  output N7760;
  output N7761;
  input N79;
  input N80;
  output N8075;
  output N8076;
  input N81;
  output N8123;
  output N8124;
  output N8127;
  output N8128;
  output N816;
  input N82;
  input N83;
  input N86;
  input N87;
  input N88;
  input N91;
  input N94;
  input N97;
  al_inv _0751_ (
    .a(N348),
    .y(N1138)
  );
  al_inv _0752_ (
    .a(N366),
    .y(N1139)
  );
  al_inv _0753_ (
    .a(N545),
    .y(N1137)
  );
  al_inv _0754_ (
    .a(N338),
    .y(N1144)
  );
  al_inv _0755_ (
    .a(N358),
    .y(N1145)
  );
  al_inv _0756_ (
    .a(N245),
    .y(N1152)
  );
  al_inv _0757_ (
    .a(N552),
    .y(N1153)
  );
  al_inv _0758_ (
    .a(N562),
    .y(N1154)
  );
  al_inv _0759_ (
    .a(N559),
    .y(N1155)
  );
  al_nand2ft _0760_ (
    .a(N591),
    .b(N27),
    .y(N2060)
  );
  al_nand2 _0761_ (
    .a(N386),
    .b(N556),
    .y(N2061)
  );
  al_inv _0762_ (
    .a(N549),
    .y(N1141)
  );
  al_nand3 _0763_ (
    .a(N27),
    .b(N31),
    .c(N140),
    .y(N2590)
  );
  al_and2 _0764_ (
    .a(N27),
    .b(N31),
    .y(_0108_)
  );
  al_inv _0765_ (
    .a(_0108_),
    .y(N2623)
  );
  al_inv _0766_ (
    .a(N299),
    .y(N3613)
  );
  al_mux2l _0767_ (
    .a(N87),
    .b(N86),
    .s(N588),
    .y(_0109_)
  );
  al_nand3 _0768_ (
    .a(N27),
    .b(N31),
    .c(_0109_),
    .y(N4272)
  );
  al_mux2l _0769_ (
    .a(N34),
    .b(N88),
    .s(N588),
    .y(_0110_)
  );
  al_nand3 _0770_ (
    .a(N27),
    .b(N31),
    .c(_0110_),
    .y(N4275)
  );
  al_nand3 _0771_ (
    .a(N27),
    .b(N31),
    .c(N83),
    .y(N4279)
  );
  al_and2ft _0772_ (
    .a(N293),
    .b(N302),
    .y(_0111_)
  );
  al_nand2ft _0773_ (
    .a(N302),
    .b(N293),
    .y(_0112_)
  );
  al_and2ft _0774_ (
    .a(N316),
    .b(N308),
    .y(_0113_)
  );
  al_nand2ft _0775_ (
    .a(N308),
    .b(N316),
    .y(_0114_)
  );
  al_nand2ft _0776_ (
    .a(_0113_),
    .b(_0114_),
    .y(_0115_)
  );
  al_or3ftt _0777_ (
    .a(_0112_),
    .b(_0111_),
    .c(_0115_),
    .y(_0116_)
  );
  al_aoi21ftf _0778_ (
    .a(_0111_),
    .b(_0112_),
    .c(_0115_),
    .y(_0117_)
  );
  al_nand2ft _0779_ (
    .a(_0117_),
    .b(_0116_),
    .y(_0118_)
  );
  al_nand2 _0780_ (
    .a(N324),
    .b(N361),
    .y(_0119_)
  );
  al_or2 _0781_ (
    .a(N324),
    .b(N361),
    .y(_0120_)
  );
  al_aoi21ttf _0782_ (
    .a(_0120_),
    .b(_0119_),
    .c(N369),
    .y(_0121_)
  );
  al_and3ftt _0783_ (
    .a(N369),
    .b(_0120_),
    .c(_0119_),
    .y(_0122_)
  );
  al_and2ft _0784_ (
    .a(N351),
    .b(N341),
    .y(_0123_)
  );
  al_nand2ft _0785_ (
    .a(N341),
    .b(N351),
    .y(_0124_)
  );
  al_nand2ft _0786_ (
    .a(_0123_),
    .b(_0124_),
    .y(_0125_)
  );
  al_or3 _0787_ (
    .a(_0122_),
    .b(_0125_),
    .c(_0121_),
    .y(_0126_)
  );
  al_oai21 _0788_ (
    .a(_0122_),
    .b(_0121_),
    .c(_0125_),
    .y(_0127_)
  );
  al_aoi21ttf _0789_ (
    .a(_0126_),
    .b(_0127_),
    .c(_0118_),
    .y(_0128_)
  );
  al_or3fft _0790_ (
    .a(_0126_),
    .b(_0127_),
    .c(_0118_),
    .y(_0129_)
  );
  al_nand2ft _0791_ (
    .a(_0128_),
    .b(_0129_),
    .y(N6716)
  );
  al_and2ft _0792_ (
    .a(N234),
    .b(N257),
    .y(_0130_)
  );
  al_nand2ft _0793_ (
    .a(N257),
    .b(N234),
    .y(_0131_)
  );
  al_nand2ft _0794_ (
    .a(_0130_),
    .b(_0131_),
    .y(_0132_)
  );
  al_nand2ft _0795_ (
    .a(N289),
    .b(N281),
    .y(_0133_)
  );
  al_nand2ft _0796_ (
    .a(N281),
    .b(N289),
    .y(_0134_)
  );
  al_nor3fft _0797_ (
    .a(_0133_),
    .b(_0134_),
    .c(_0132_),
    .y(_0135_)
  );
  al_ao21ttf _0798_ (
    .a(_0133_),
    .b(_0134_),
    .c(_0132_),
    .y(_0136_)
  );
  al_and2ft _0799_ (
    .a(N265),
    .b(N273),
    .y(_0137_)
  );
  al_nand2ft _0800_ (
    .a(N273),
    .b(N265),
    .y(_0138_)
  );
  al_nand2ft _0801_ (
    .a(_0137_),
    .b(_0138_),
    .y(_0139_)
  );
  al_oai21ftt _0802_ (
    .a(_0136_),
    .b(_0135_),
    .c(_0139_),
    .y(_0140_)
  );
  al_or3ftt _0803_ (
    .a(_0136_),
    .b(_0135_),
    .c(_0139_),
    .y(_0141_)
  );
  al_and2ft _0804_ (
    .a(N210),
    .b(N206),
    .y(_0142_)
  );
  al_nand2ft _0805_ (
    .a(N206),
    .b(N210),
    .y(_0143_)
  );
  al_and2ft _0806_ (
    .a(N226),
    .b(N218),
    .y(_0144_)
  );
  al_nand2ft _0807_ (
    .a(N218),
    .b(N226),
    .y(_0145_)
  );
  al_nand2ft _0808_ (
    .a(_0144_),
    .b(_0145_),
    .y(_0146_)
  );
  al_and3ftt _0809_ (
    .a(_0142_),
    .b(_0143_),
    .c(_0146_),
    .y(_0147_)
  );
  al_ao21ftt _0810_ (
    .a(_0142_),
    .b(_0143_),
    .c(_0146_),
    .y(_0148_)
  );
  al_nand2ft _0811_ (
    .a(_0147_),
    .b(_0148_),
    .y(_0149_)
  );
  al_nand3 _0812_ (
    .a(_0140_),
    .b(_0141_),
    .c(_0149_),
    .y(_0150_)
  );
  al_aoi21 _0813_ (
    .a(_0140_),
    .b(_0141_),
    .c(_0149_),
    .y(_0151_)
  );
  al_nand2ft _0814_ (
    .a(_0151_),
    .b(_0150_),
    .y(N6877)
  );
  al_and3ftt _0815_ (
    .a(N619),
    .b(N625),
    .c(N131),
    .y(_0152_)
  );
  al_inv _0816_ (
    .a(N619),
    .y(_0153_)
  );
  al_mux2l _0817_ (
    .a(N366),
    .b(N361),
    .s(N332),
    .y(_0154_)
  );
  al_or2ft _0818_ (
    .a(N54),
    .b(_0154_),
    .y(_0155_)
  );
  al_and2ft _0819_ (
    .a(N54),
    .b(_0154_),
    .y(_0156_)
  );
  al_oai21ftf _0820_ (
    .a(_0155_),
    .b(_0156_),
    .c(_0153_),
    .y(_0157_)
  );
  al_inv _0821_ (
    .a(N625),
    .y(_0158_)
  );
  al_mux2l _0822_ (
    .a(N248),
    .b(N251),
    .s(N361),
    .y(_0159_)
  );
  al_aoi21ftf _0823_ (
    .a(N619),
    .b(_0159_),
    .c(_0158_),
    .y(_0160_)
  );
  al_aoi21 _0824_ (
    .a(_0160_),
    .b(_0157_),
    .c(_0152_),
    .y(N7015)
  );
  al_and2ft _0825_ (
    .a(N619),
    .b(N625),
    .y(_0161_)
  );
  al_inv _0826_ (
    .a(_0161_),
    .y(_0162_)
  );
  al_inv _0827_ (
    .a(N54),
    .y(_0163_)
  );
  al_mux2l _0828_ (
    .a(N358),
    .b(N351),
    .s(N332),
    .y(_0164_)
  );
  al_or2 _0829_ (
    .a(N534),
    .b(_0164_),
    .y(_0165_)
  );
  al_nand2 _0830_ (
    .a(N534),
    .b(_0164_),
    .y(_0166_)
  );
  al_nand2 _0831_ (
    .a(_0166_),
    .b(_0165_),
    .y(_0167_)
  );
  al_ao21 _0832_ (
    .a(N534),
    .b(_0164_),
    .c(_0154_),
    .y(_0168_)
  );
  al_ao21ttf _0833_ (
    .a(_0166_),
    .b(_0165_),
    .c(_0154_),
    .y(_0169_)
  );
  al_ao21ftf _0834_ (
    .a(_0168_),
    .b(_0165_),
    .c(_0169_),
    .y(_0170_)
  );
  al_mux2h _0835_ (
    .a(_0167_),
    .b(_0170_),
    .s(_0163_),
    .y(_0171_)
  );
  al_inv _0836_ (
    .a(N534),
    .y(_0172_)
  );
  al_mux2l _0837_ (
    .a(N598),
    .b(N597),
    .s(N351),
    .y(_0173_)
  );
  al_inv _0838_ (
    .a(N595),
    .y(_0174_)
  );
  al_inv _0839_ (
    .a(N596),
    .y(_0175_)
  );
  al_mux2l _0840_ (
    .a(_0174_),
    .b(_0175_),
    .s(N351),
    .y(_0176_)
  );
  al_mux2h _0841_ (
    .a(_0173_),
    .b(_0176_),
    .s(_0172_),
    .y(_0177_)
  );
  al_mux2h _0842_ (
    .a(_0177_),
    .b(_0171_),
    .s(N619),
    .y(_0178_)
  );
  al_nand2 _0843_ (
    .a(_0158_),
    .b(_0178_),
    .y(_0179_)
  );
  al_ao21ftf _0844_ (
    .a(_0162_),
    .b(N129),
    .c(_0179_),
    .y(_0180_)
  );
  al_inv _0845_ (
    .a(_0180_),
    .y(N7363)
  );
  al_mux2l _0846_ (
    .a(N288),
    .b(N281),
    .s(N335),
    .y(_0181_)
  );
  al_nand2 _0847_ (
    .a(N374),
    .b(_0181_),
    .y(_0182_)
  );
  al_or2 _0848_ (
    .a(N374),
    .b(_0181_),
    .y(_0183_)
  );
  al_nand3 _0849_ (
    .a(N4),
    .b(_0182_),
    .c(_0183_),
    .y(_0184_)
  );
  al_aoi21 _0850_ (
    .a(_0182_),
    .b(_0183_),
    .c(N4),
    .y(_0185_)
  );
  al_or2ft _0851_ (
    .a(_0184_),
    .b(_0185_),
    .y(_0186_)
  );
  al_inv _0852_ (
    .a(N597),
    .y(_0187_)
  );
  al_inv _0853_ (
    .a(N598),
    .y(_0188_)
  );
  al_mux2l _0854_ (
    .a(_0188_),
    .b(_0187_),
    .s(N281),
    .y(_0189_)
  );
  al_mux2l _0855_ (
    .a(N595),
    .b(N596),
    .s(N281),
    .y(_0190_)
  );
  al_mux2h _0856_ (
    .a(_0190_),
    .b(_0189_),
    .s(N374),
    .y(_0191_)
  );
  al_aoi21 _0857_ (
    .a(_0153_),
    .b(_0191_),
    .c(N625),
    .y(_0192_)
  );
  al_ao21ftf _0858_ (
    .a(_0153_),
    .b(_0186_),
    .c(_0192_),
    .y(_0193_)
  );
  al_aoi21ftf _0859_ (
    .a(_0162_),
    .b(N117),
    .c(_0193_),
    .y(N7365)
  );
  al_inv _0860_ (
    .a(N331),
    .y(_0194_)
  );
  al_nand2ft _0861_ (
    .a(N338),
    .b(N332),
    .y(_0195_)
  );
  al_mux2l _0862_ (
    .a(N331),
    .b(N324),
    .s(N332),
    .y(_0196_)
  );
  al_mux2l _0863_ (
    .a(_0196_),
    .b(_0194_),
    .s(_0195_),
    .y(_0197_)
  );
  al_mux2l _0864_ (
    .a(N307),
    .b(N302),
    .s(N332),
    .y(_0198_)
  );
  al_mux2l _0865_ (
    .a(N299),
    .b(N293),
    .s(N332),
    .y(_0199_)
  );
  al_or2 _0866_ (
    .a(_0198_),
    .b(_0199_),
    .y(_0200_)
  );
  al_nand2 _0867_ (
    .a(_0198_),
    .b(_0199_),
    .y(_0201_)
  );
  al_and3ftt _0868_ (
    .a(_0197_),
    .b(_0200_),
    .c(_0201_),
    .y(_0202_)
  );
  al_ao21ttf _0869_ (
    .a(_0200_),
    .b(_0201_),
    .c(_0197_),
    .y(_0203_)
  );
  al_and2ft _0870_ (
    .a(_0202_),
    .b(_0203_),
    .y(_0204_)
  );
  al_mux2l _0871_ (
    .a(N323),
    .b(N316),
    .s(N332),
    .y(_0205_)
  );
  al_mux2l _0872_ (
    .a(N315),
    .b(N308),
    .s(N332),
    .y(_0206_)
  );
  al_and2ft _0873_ (
    .a(_0205_),
    .b(_0206_),
    .y(_0207_)
  );
  al_nand2ft _0874_ (
    .a(_0206_),
    .b(_0205_),
    .y(_0208_)
  );
  al_nand2ft _0875_ (
    .a(_0207_),
    .b(_0208_),
    .y(_0209_)
  );
  al_mux2l _0876_ (
    .a(N372),
    .b(N369),
    .s(N332),
    .y(_0210_)
  );
  al_mux2l _0877_ (
    .a(N348),
    .b(N341),
    .s(N332),
    .y(_0211_)
  );
  al_and2ft _0878_ (
    .a(_0211_),
    .b(_0210_),
    .y(_0212_)
  );
  al_nand2ft _0879_ (
    .a(_0210_),
    .b(_0211_),
    .y(_0213_)
  );
  al_nand3ftt _0880_ (
    .a(_0212_),
    .b(_0213_),
    .c(_0209_),
    .y(_0214_)
  );
  al_ao21ftt _0881_ (
    .a(_0212_),
    .b(_0213_),
    .c(_0209_),
    .y(_0215_)
  );
  al_nand2 _0882_ (
    .a(_0154_),
    .b(_0164_),
    .y(_0216_)
  );
  al_nor2 _0883_ (
    .a(_0154_),
    .b(_0164_),
    .y(_0217_)
  );
  al_and2ft _0884_ (
    .a(_0217_),
    .b(_0216_),
    .y(_0218_)
  );
  al_ao21 _0885_ (
    .a(_0214_),
    .b(_0215_),
    .c(_0218_),
    .y(_0219_)
  );
  al_nand3 _0886_ (
    .a(_0218_),
    .b(_0214_),
    .c(_0215_),
    .y(_0220_)
  );
  al_ao21 _0887_ (
    .a(_0220_),
    .b(_0219_),
    .c(_0204_),
    .y(_0221_)
  );
  al_and3 _0888_ (
    .a(_0204_),
    .b(_0220_),
    .c(_0219_),
    .y(_0222_)
  );
  al_nand2ft _0889_ (
    .a(_0222_),
    .b(_0221_),
    .y(N7474)
  );
  al_mux2l _0890_ (
    .a(N272),
    .b(N265),
    .s(N335),
    .y(_0223_)
  );
  al_mux2l _0891_ (
    .a(N280),
    .b(N273),
    .s(N335),
    .y(_0224_)
  );
  al_nand2 _0892_ (
    .a(_0181_),
    .b(_0224_),
    .y(_0225_)
  );
  al_or2 _0893_ (
    .a(_0181_),
    .b(_0224_),
    .y(_0226_)
  );
  al_and3 _0894_ (
    .a(_0223_),
    .b(_0226_),
    .c(_0225_),
    .y(_0227_)
  );
  al_ao21 _0895_ (
    .a(_0226_),
    .b(_0225_),
    .c(_0223_),
    .y(_0228_)
  );
  al_and2ft _0896_ (
    .a(_0227_),
    .b(_0228_),
    .y(_0229_)
  );
  al_mux2l _0897_ (
    .a(N209),
    .b(N206),
    .s(N335),
    .y(_0230_)
  );
  al_mux2l _0898_ (
    .a(N292),
    .b(N289),
    .s(N335),
    .y(_0231_)
  );
  al_nand2ft _0899_ (
    .a(_0231_),
    .b(_0230_),
    .y(_0232_)
  );
  al_nand2ft _0900_ (
    .a(_0230_),
    .b(_0231_),
    .y(_0233_)
  );
  al_mux2l _0901_ (
    .a(N264),
    .b(N257),
    .s(N335),
    .y(_0234_)
  );
  al_and3 _0902_ (
    .a(_0234_),
    .b(_0232_),
    .c(_0233_),
    .y(_0235_)
  );
  al_ao21 _0903_ (
    .a(_0232_),
    .b(_0233_),
    .c(_0234_),
    .y(_0236_)
  );
  al_nand2ft _0904_ (
    .a(_0235_),
    .b(_0236_),
    .y(_0237_)
  );
  al_mux2l _0905_ (
    .a(N241),
    .b(N234),
    .s(N335),
    .y(_0238_)
  );
  al_mux2l _0906_ (
    .a(N233),
    .b(N226),
    .s(N335),
    .y(_0239_)
  );
  al_and2ft _0907_ (
    .a(_0238_),
    .b(_0239_),
    .y(_0240_)
  );
  al_nand2ft _0908_ (
    .a(_0239_),
    .b(_0238_),
    .y(_0241_)
  );
  al_mux2l _0909_ (
    .a(N225),
    .b(N218),
    .s(N335),
    .y(_0242_)
  );
  al_mux2l _0910_ (
    .a(N217),
    .b(N210),
    .s(N335),
    .y(_0243_)
  );
  al_nand2 _0911_ (
    .a(_0242_),
    .b(_0243_),
    .y(_0244_)
  );
  al_nor2 _0912_ (
    .a(_0242_),
    .b(_0243_),
    .y(_0245_)
  );
  al_and2ft _0913_ (
    .a(_0245_),
    .b(_0244_),
    .y(_0246_)
  );
  al_nand3ftt _0914_ (
    .a(_0240_),
    .b(_0241_),
    .c(_0246_),
    .y(_0247_)
  );
  al_ao21ftt _0915_ (
    .a(_0240_),
    .b(_0241_),
    .c(_0246_),
    .y(_0248_)
  );
  al_ao21 _0916_ (
    .a(_0247_),
    .b(_0248_),
    .c(_0237_),
    .y(_0249_)
  );
  al_nand3 _0917_ (
    .a(_0247_),
    .b(_0237_),
    .c(_0248_),
    .y(_0250_)
  );
  al_aoi21 _0918_ (
    .a(_0249_),
    .b(_0250_),
    .c(_0229_),
    .y(_0251_)
  );
  al_nand3 _0919_ (
    .a(_0229_),
    .b(_0249_),
    .c(_0250_),
    .y(_0252_)
  );
  al_or2ft _0920_ (
    .a(_0252_),
    .b(_0251_),
    .y(N7476)
  );
  al_and2 _0921_ (
    .a(N479),
    .b(_0206_),
    .y(_0253_)
  );
  al_or2 _0922_ (
    .a(N479),
    .b(_0206_),
    .y(_0254_)
  );
  al_and2 _0923_ (
    .a(N490),
    .b(_0205_),
    .y(_0255_)
  );
  al_ao21 _0924_ (
    .a(_0255_),
    .b(_0254_),
    .c(_0253_),
    .y(_0256_)
  );
  al_nand2 _0925_ (
    .a(N479),
    .b(_0206_),
    .y(_0257_)
  );
  al_or2 _0926_ (
    .a(N490),
    .b(_0205_),
    .y(_0258_)
  );
  al_and2ft _0927_ (
    .a(_0255_),
    .b(_0258_),
    .y(_0259_)
  );
  al_and3 _0928_ (
    .a(_0257_),
    .b(_0254_),
    .c(_0259_),
    .y(_0260_)
  );
  al_and2 _0929_ (
    .a(N503),
    .b(_0196_),
    .y(_0261_)
  );
  al_nor2 _0930_ (
    .a(N503),
    .b(_0196_),
    .y(_0262_)
  );
  al_and3fft _0931_ (
    .a(N338),
    .b(N514),
    .c(N332),
    .y(_0263_)
  );
  al_oai21ftt _0932_ (
    .a(N332),
    .b(N338),
    .c(N514),
    .y(_0264_)
  );
  al_nand2 _0933_ (
    .a(N523),
    .b(_0211_),
    .y(_0265_)
  );
  al_or2 _0934_ (
    .a(N523),
    .b(_0211_),
    .y(_0266_)
  );
  al_nand3 _0935_ (
    .a(_0165_),
    .b(_0168_),
    .c(_0266_),
    .y(_0267_)
  );
  al_nand3 _0936_ (
    .a(_0264_),
    .b(_0265_),
    .c(_0267_),
    .y(_0268_)
  );
  al_nand3fft _0937_ (
    .a(_0262_),
    .b(_0263_),
    .c(_0268_),
    .y(_0269_)
  );
  al_and2ft _0938_ (
    .a(_0261_),
    .b(_0269_),
    .y(_0270_)
  );
  al_nand3ftt _0939_ (
    .a(_0154_),
    .b(_0166_),
    .c(_0165_),
    .y(_0271_)
  );
  al_and2ft _0940_ (
    .a(_0263_),
    .b(_0264_),
    .y(_0272_)
  );
  al_nand3 _0941_ (
    .a(_0265_),
    .b(_0266_),
    .c(_0272_),
    .y(_0273_)
  );
  al_or2 _0942_ (
    .a(_0261_),
    .b(_0262_),
    .y(_0274_)
  );
  al_or3 _0943_ (
    .a(_0271_),
    .b(_0274_),
    .c(_0273_),
    .y(_0275_)
  );
  al_ao21ftf _0944_ (
    .a(_0275_),
    .b(N54),
    .c(_0270_),
    .y(_0276_)
  );
  al_aoi21 _0945_ (
    .a(_0260_),
    .b(_0276_),
    .c(_0256_),
    .y(_0277_)
  );
  al_ao21ftf _0946_ (
    .a(_0198_),
    .b(_0277_),
    .c(_0199_),
    .y(_0278_)
  );
  al_aoi21ftf _0947_ (
    .a(_0200_),
    .b(_0277_),
    .c(_0278_),
    .y(N7432)
  );
  al_nand2ft _0948_ (
    .a(_0263_),
    .b(_0268_),
    .y(_0279_)
  );
  al_or2 _0949_ (
    .a(_0271_),
    .b(_0273_),
    .y(_0280_)
  );
  al_ao21ftf _0950_ (
    .a(_0280_),
    .b(N54),
    .c(_0279_),
    .y(_0281_)
  );
  al_or3 _0951_ (
    .a(_0261_),
    .b(_0262_),
    .c(_0281_),
    .y(_0282_)
  );
  al_and2 _0952_ (
    .a(_0274_),
    .b(_0281_),
    .y(_0283_)
  );
  al_and2ft _0953_ (
    .a(_0283_),
    .b(_0282_),
    .y(_0284_)
  );
  al_mux2l _0954_ (
    .a(_0188_),
    .b(_0187_),
    .s(N324),
    .y(_0285_)
  );
  al_mux2l _0955_ (
    .a(N595),
    .b(N596),
    .s(N324),
    .y(_0286_)
  );
  al_mux2h _0956_ (
    .a(_0286_),
    .b(_0285_),
    .s(N503),
    .y(_0287_)
  );
  al_ao21 _0957_ (
    .a(_0153_),
    .b(_0287_),
    .c(N625),
    .y(_0288_)
  );
  al_ao21 _0958_ (
    .a(N619),
    .b(_0284_),
    .c(_0288_),
    .y(_0289_)
  );
  al_aoi21ftf _0959_ (
    .a(_0162_),
    .b(N52),
    .c(_0289_),
    .y(N7465)
  );
  al_oa21ftt _0960_ (
    .a(_0163_),
    .b(_0168_),
    .c(_0165_),
    .y(_0290_)
  );
  al_oai21ftt _0961_ (
    .a(_0265_),
    .b(_0290_),
    .c(_0266_),
    .y(_0291_)
  );
  al_and2ft _0962_ (
    .a(_0272_),
    .b(_0291_),
    .y(_0292_)
  );
  al_or3ftt _0963_ (
    .a(_0264_),
    .b(_0263_),
    .c(_0291_),
    .y(_0293_)
  );
  al_nand2ft _0964_ (
    .a(_0292_),
    .b(_0293_),
    .y(_0294_)
  );
  al_mux2h _0965_ (
    .a(N595),
    .b(_0188_),
    .s(N514),
    .y(_0295_)
  );
  al_aoi21 _0966_ (
    .a(_0153_),
    .b(_0295_),
    .c(N625),
    .y(_0296_)
  );
  al_ao21ttf _0967_ (
    .a(N619),
    .b(_0294_),
    .c(_0296_),
    .y(_0297_)
  );
  al_ao21ftf _0968_ (
    .a(_0162_),
    .b(N130),
    .c(_0297_),
    .y(_0298_)
  );
  al_inv _0969_ (
    .a(_0298_),
    .y(N7466)
  );
  al_and3 _0970_ (
    .a(_0265_),
    .b(_0266_),
    .c(_0290_),
    .y(_0299_)
  );
  al_ao21 _0971_ (
    .a(_0265_),
    .b(_0266_),
    .c(_0290_),
    .y(_0300_)
  );
  al_nand2ft _0972_ (
    .a(_0299_),
    .b(_0300_),
    .y(_0301_)
  );
  al_mux2l _0973_ (
    .a(_0188_),
    .b(_0187_),
    .s(N341),
    .y(_0302_)
  );
  al_mux2l _0974_ (
    .a(N595),
    .b(N596),
    .s(N341),
    .y(_0303_)
  );
  al_mux2h _0975_ (
    .a(_0303_),
    .b(_0302_),
    .s(N523),
    .y(_0304_)
  );
  al_ao21 _0976_ (
    .a(_0153_),
    .b(_0304_),
    .c(N625),
    .y(_0305_)
  );
  al_ao21 _0977_ (
    .a(N619),
    .b(_0301_),
    .c(_0305_),
    .y(_0306_)
  );
  al_aoi21ftf _0978_ (
    .a(_0162_),
    .b(N119),
    .c(_0306_),
    .y(N7467)
  );
  al_and2 _0979_ (
    .a(N435),
    .b(_0238_),
    .y(_0307_)
  );
  al_or2 _0980_ (
    .a(N435),
    .b(_0238_),
    .y(_0308_)
  );
  al_nand2ft _0981_ (
    .a(_0307_),
    .b(_0308_),
    .y(_0309_)
  );
  al_or2 _0982_ (
    .a(N389),
    .b(_0234_),
    .y(_0310_)
  );
  al_and2 _0983_ (
    .a(N389),
    .b(_0234_),
    .y(_0311_)
  );
  al_inv _0984_ (
    .a(_0311_),
    .y(_0312_)
  );
  al_or2 _0985_ (
    .a(N400),
    .b(_0223_),
    .y(_0313_)
  );
  al_and2 _0986_ (
    .a(N400),
    .b(_0223_),
    .y(_0314_)
  );
  al_nand2ft _0987_ (
    .a(_0314_),
    .b(_0313_),
    .y(_0315_)
  );
  al_or2 _0988_ (
    .a(N411),
    .b(_0224_),
    .y(_0316_)
  );
  al_inv _0989_ (
    .a(N374),
    .y(_0317_)
  );
  al_nand2 _0990_ (
    .a(N411),
    .b(_0224_),
    .y(_0318_)
  );
  al_aoi21ftf _0991_ (
    .a(_0317_),
    .b(_0181_),
    .c(_0318_),
    .y(_0319_)
  );
  al_and3 _0992_ (
    .a(_0183_),
    .b(_0316_),
    .c(_0319_),
    .y(_0320_)
  );
  al_nand2ft _0993_ (
    .a(_0315_),
    .b(_0320_),
    .y(_0321_)
  );
  al_nand3 _0994_ (
    .a(N374),
    .b(_0181_),
    .c(_0316_),
    .y(_0322_)
  );
  al_inv _0995_ (
    .a(N400),
    .y(_0323_)
  );
  al_aoi21ftf _0996_ (
    .a(_0323_),
    .b(_0223_),
    .c(_0318_),
    .y(_0324_)
  );
  al_aoi21ttf _0997_ (
    .a(_0324_),
    .b(_0322_),
    .c(_0313_),
    .y(_0325_)
  );
  al_oa21ftf _0998_ (
    .a(N4),
    .b(_0321_),
    .c(_0325_),
    .y(_0326_)
  );
  al_ao21ttf _0999_ (
    .a(_0312_),
    .b(_0326_),
    .c(_0310_),
    .y(_0327_)
  );
  al_and2 _1000_ (
    .a(_0309_),
    .b(_0327_),
    .y(_0328_)
  );
  al_or3ftt _1001_ (
    .a(_0308_),
    .b(_0307_),
    .c(_0327_),
    .y(_0329_)
  );
  al_nand2ft _1002_ (
    .a(_0328_),
    .b(_0329_),
    .y(_0330_)
  );
  al_mux2l _1003_ (
    .a(_0188_),
    .b(_0187_),
    .s(N234),
    .y(_0331_)
  );
  al_mux2l _1004_ (
    .a(N595),
    .b(N596),
    .s(N234),
    .y(_0332_)
  );
  al_mux2h _1005_ (
    .a(_0332_),
    .b(_0331_),
    .s(N435),
    .y(_0333_)
  );
  al_ao21 _1006_ (
    .a(_0153_),
    .b(_0333_),
    .c(N625),
    .y(_0334_)
  );
  al_ao21 _1007_ (
    .a(N619),
    .b(_0330_),
    .c(_0334_),
    .y(_0335_)
  );
  al_aoi21ftf _1008_ (
    .a(_0162_),
    .b(N122),
    .c(_0335_),
    .y(N7470)
  );
  al_and2ft _1009_ (
    .a(_0311_),
    .b(_0310_),
    .y(_0336_)
  );
  al_and2ft _1010_ (
    .a(_0336_),
    .b(_0326_),
    .y(_0337_)
  );
  al_or3fft _1011_ (
    .a(_0310_),
    .b(_0312_),
    .c(_0326_),
    .y(_0338_)
  );
  al_nand2ft _1012_ (
    .a(_0337_),
    .b(_0338_),
    .y(_0339_)
  );
  al_mux2l _1013_ (
    .a(_0188_),
    .b(_0187_),
    .s(N257),
    .y(_0340_)
  );
  al_mux2l _1014_ (
    .a(N595),
    .b(N596),
    .s(N257),
    .y(_0341_)
  );
  al_mux2h _1015_ (
    .a(_0341_),
    .b(_0340_),
    .s(N389),
    .y(_0342_)
  );
  al_aoi21 _1016_ (
    .a(_0153_),
    .b(_0342_),
    .c(N625),
    .y(_0343_)
  );
  al_ao21ttf _1017_ (
    .a(N619),
    .b(_0339_),
    .c(_0343_),
    .y(_0344_)
  );
  al_ao21ftf _1018_ (
    .a(_0162_),
    .b(N128),
    .c(_0344_),
    .y(_0345_)
  );
  al_inv _1019_ (
    .a(_0345_),
    .y(N7471)
  );
  al_nor2 _1020_ (
    .a(N411),
    .b(_0224_),
    .y(_0346_)
  );
  al_ao21 _1021_ (
    .a(_0319_),
    .b(_0184_),
    .c(_0346_),
    .y(_0347_)
  );
  al_or2 _1022_ (
    .a(_0315_),
    .b(_0347_),
    .y(_0348_)
  );
  al_and2 _1023_ (
    .a(_0315_),
    .b(_0347_),
    .y(_0349_)
  );
  al_nand2ft _1024_ (
    .a(_0349_),
    .b(_0348_),
    .y(_0350_)
  );
  al_mux2l _1025_ (
    .a(_0188_),
    .b(_0187_),
    .s(N265),
    .y(_0351_)
  );
  al_mux2l _1026_ (
    .a(N595),
    .b(N596),
    .s(N265),
    .y(_0352_)
  );
  al_mux2h _1027_ (
    .a(_0352_),
    .b(_0351_),
    .s(N400),
    .y(_0353_)
  );
  al_aoi21 _1028_ (
    .a(_0153_),
    .b(_0353_),
    .c(N625),
    .y(_0354_)
  );
  al_ao21ttf _1029_ (
    .a(N619),
    .b(_0350_),
    .c(_0354_),
    .y(_0355_)
  );
  al_aoi21ftf _1030_ (
    .a(_0162_),
    .b(N127),
    .c(_0355_),
    .y(N7472)
  );
  al_aoi21ttf _1031_ (
    .a(N4),
    .b(_0183_),
    .c(_0182_),
    .y(_0356_)
  );
  al_aoi21ftf _1032_ (
    .a(_0346_),
    .b(_0318_),
    .c(_0356_),
    .y(_0357_)
  );
  al_or3fft _1033_ (
    .a(_0316_),
    .b(_0318_),
    .c(_0356_),
    .y(_0358_)
  );
  al_nand2ft _1034_ (
    .a(_0357_),
    .b(_0358_),
    .y(_0359_)
  );
  al_mux2l _1035_ (
    .a(_0188_),
    .b(_0187_),
    .s(N273),
    .y(_0360_)
  );
  al_mux2l _1036_ (
    .a(N595),
    .b(N596),
    .s(N273),
    .y(_0361_)
  );
  al_mux2h _1037_ (
    .a(_0361_),
    .b(_0360_),
    .s(N411),
    .y(_0362_)
  );
  al_ao21 _1038_ (
    .a(_0153_),
    .b(_0362_),
    .c(N625),
    .y(_0363_)
  );
  al_ao21 _1039_ (
    .a(N619),
    .b(_0359_),
    .c(_0363_),
    .y(_0364_)
  );
  al_ao21ftf _1040_ (
    .a(_0162_),
    .b(N126),
    .c(_0364_),
    .y(_0365_)
  );
  al_inv _1041_ (
    .a(_0365_),
    .y(N7473)
  );
  al_and3ftt _1042_ (
    .a(N619),
    .b(N625),
    .c(N123),
    .y(_0366_)
  );
  al_mux2l _1043_ (
    .a(N242),
    .b(N254),
    .s(N293),
    .y(_0367_)
  );
  al_oa21ttf _1044_ (
    .a(N619),
    .b(_0367_),
    .c(N625),
    .y(_0368_)
  );
  al_ao21ttf _1045_ (
    .a(N619),
    .b(N7432),
    .c(_0368_),
    .y(_0369_)
  );
  al_and2ft _1046_ (
    .a(_0366_),
    .b(_0369_),
    .y(N7699)
  );
  al_and3ftt _1047_ (
    .a(N619),
    .b(N625),
    .c(N121),
    .y(_0370_)
  );
  al_and2ft _1048_ (
    .a(_0198_),
    .b(_0277_),
    .y(_0371_)
  );
  al_or2ft _1049_ (
    .a(_0198_),
    .b(_0277_),
    .y(_0372_)
  );
  al_or3fft _1050_ (
    .a(N619),
    .b(_0372_),
    .c(_0371_),
    .y(_0373_)
  );
  al_mux2l _1051_ (
    .a(N248),
    .b(N251),
    .s(N302),
    .y(_0374_)
  );
  al_aoi21ftf _1052_ (
    .a(N619),
    .b(_0374_),
    .c(_0158_),
    .y(_0375_)
  );
  al_aoi21 _1053_ (
    .a(_0375_),
    .b(_0373_),
    .c(_0370_),
    .y(N7700)
  );
  al_oa21 _1054_ (
    .a(_0255_),
    .b(_0276_),
    .c(_0258_),
    .y(_0376_)
  );
  al_or3fft _1055_ (
    .a(_0257_),
    .b(_0254_),
    .c(_0376_),
    .y(_0377_)
  );
  al_aoi21ftf _1056_ (
    .a(_0253_),
    .b(_0254_),
    .c(_0376_),
    .y(_0378_)
  );
  al_and2ft _1057_ (
    .a(_0378_),
    .b(_0377_),
    .y(_0379_)
  );
  al_mux2l _1058_ (
    .a(N248),
    .b(N251),
    .s(N308),
    .y(_0380_)
  );
  al_inv _1059_ (
    .a(N242),
    .y(_0381_)
  );
  al_inv _1060_ (
    .a(N254),
    .y(_0382_)
  );
  al_mux2l _1061_ (
    .a(_0381_),
    .b(_0382_),
    .s(N308),
    .y(_0383_)
  );
  al_mux2l _1062_ (
    .a(_0380_),
    .b(_0383_),
    .s(N479),
    .y(_0384_)
  );
  al_ao21 _1063_ (
    .a(_0153_),
    .b(_0384_),
    .c(N625),
    .y(_0385_)
  );
  al_ao21 _1064_ (
    .a(N619),
    .b(_0379_),
    .c(_0385_),
    .y(_0386_)
  );
  al_aoi21ftf _1065_ (
    .a(_0162_),
    .b(N116),
    .c(_0386_),
    .y(N7701)
  );
  al_and2 _1066_ (
    .a(_0259_),
    .b(_0276_),
    .y(_0387_)
  );
  al_or2 _1067_ (
    .a(_0259_),
    .b(_0276_),
    .y(_0388_)
  );
  al_nand2ft _1068_ (
    .a(_0387_),
    .b(_0388_),
    .y(_0389_)
  );
  al_mux2l _1069_ (
    .a(N248),
    .b(N251),
    .s(N316),
    .y(_0390_)
  );
  al_mux2l _1070_ (
    .a(_0381_),
    .b(_0382_),
    .s(N316),
    .y(_0391_)
  );
  al_mux2l _1071_ (
    .a(_0390_),
    .b(_0391_),
    .s(N490),
    .y(_0392_)
  );
  al_ao21 _1072_ (
    .a(_0153_),
    .b(_0392_),
    .c(N625),
    .y(_0393_)
  );
  al_ao21 _1073_ (
    .a(N619),
    .b(_0389_),
    .c(_0393_),
    .y(_0394_)
  );
  al_aoi21ftf _1074_ (
    .a(_0162_),
    .b(N112),
    .c(_0394_),
    .y(N7702)
  );
  al_and3ftt _1075_ (
    .a(N619),
    .b(N625),
    .c(N115),
    .y(_0395_)
  );
  al_and2 _1076_ (
    .a(N446),
    .b(_0230_),
    .y(_0396_)
  );
  al_or2 _1077_ (
    .a(N446),
    .b(_0230_),
    .y(_0397_)
  );
  al_and2 _1078_ (
    .a(N457),
    .b(_0243_),
    .y(_0398_)
  );
  al_or2 _1079_ (
    .a(N457),
    .b(_0243_),
    .y(_0399_)
  );
  al_and2 _1080_ (
    .a(N468),
    .b(_0242_),
    .y(_0400_)
  );
  al_and2 _1081_ (
    .a(N422),
    .b(_0239_),
    .y(_0401_)
  );
  al_or2 _1082_ (
    .a(N468),
    .b(_0242_),
    .y(_0402_)
  );
  al_ao21 _1083_ (
    .a(_0401_),
    .b(_0402_),
    .c(_0400_),
    .y(_0403_)
  );
  al_aoi21 _1084_ (
    .a(_0399_),
    .b(_0403_),
    .c(_0398_),
    .y(_0404_)
  );
  al_and2ft _1085_ (
    .a(_0398_),
    .b(_0399_),
    .y(_0405_)
  );
  al_nand2ft _1086_ (
    .a(_0400_),
    .b(_0402_),
    .y(_0406_)
  );
  al_nor2 _1087_ (
    .a(N422),
    .b(_0239_),
    .y(_0407_)
  );
  al_nor2 _1088_ (
    .a(_0401_),
    .b(_0407_),
    .y(_0408_)
  );
  al_nand3ftt _1089_ (
    .a(_0406_),
    .b(_0405_),
    .c(_0408_),
    .y(_0409_)
  );
  al_and2 _1090_ (
    .a(N411),
    .b(_0224_),
    .y(_0410_)
  );
  al_nand3fft _1091_ (
    .a(_0314_),
    .b(_0410_),
    .c(_0322_),
    .y(_0411_)
  );
  al_nand3 _1092_ (
    .a(_0310_),
    .b(_0313_),
    .c(_0411_),
    .y(_0412_)
  );
  al_nand3fft _1093_ (
    .a(_0307_),
    .b(_0311_),
    .c(_0412_),
    .y(_0413_)
  );
  al_nand2 _1094_ (
    .a(_0308_),
    .b(_0413_),
    .y(_0414_)
  );
  al_and3fft _1095_ (
    .a(_0309_),
    .b(_0321_),
    .c(_0336_),
    .y(_0415_)
  );
  al_ao21ttf _1096_ (
    .a(N4),
    .b(_0415_),
    .c(_0414_),
    .y(_0416_)
  );
  al_ao21ftf _1097_ (
    .a(_0409_),
    .b(_0416_),
    .c(_0404_),
    .y(_0417_)
  );
  al_or3ftt _1098_ (
    .a(_0397_),
    .b(_0396_),
    .c(_0417_),
    .y(_0418_)
  );
  al_nand2ft _1099_ (
    .a(_0396_),
    .b(_0397_),
    .y(_0419_)
  );
  al_nand2 _1100_ (
    .a(_0419_),
    .b(_0417_),
    .y(_0420_)
  );
  al_nand3 _1101_ (
    .a(N619),
    .b(_0420_),
    .c(_0418_),
    .y(_0421_)
  );
  al_mux2l _1102_ (
    .a(N248),
    .b(N251),
    .s(N206),
    .y(_0422_)
  );
  al_mux2l _1103_ (
    .a(_0381_),
    .b(_0382_),
    .s(N206),
    .y(_0423_)
  );
  al_mux2l _1104_ (
    .a(_0422_),
    .b(_0423_),
    .s(N446),
    .y(_0424_)
  );
  al_aoi21 _1105_ (
    .a(_0153_),
    .b(_0424_),
    .c(N625),
    .y(_0425_)
  );
  al_aoi21 _1106_ (
    .a(_0425_),
    .b(_0421_),
    .c(_0395_),
    .y(N7704)
  );
  al_inv _1107_ (
    .a(_0403_),
    .y(_0426_)
  );
  al_nand2 _1108_ (
    .a(N468),
    .b(_0242_),
    .y(_0427_)
  );
  al_ao21ttf _1109_ (
    .a(_0427_),
    .b(_0407_),
    .c(_0402_),
    .y(_0428_)
  );
  al_mux2l _1110_ (
    .a(_0428_),
    .b(_0426_),
    .s(_0416_),
    .y(_0429_)
  );
  al_or2 _1111_ (
    .a(_0405_),
    .b(_0429_),
    .y(_0430_)
  );
  al_nand2 _1112_ (
    .a(_0405_),
    .b(_0429_),
    .y(_0431_)
  );
  al_nand3 _1113_ (
    .a(N619),
    .b(_0431_),
    .c(_0430_),
    .y(_0432_)
  );
  al_mux2l _1114_ (
    .a(_0188_),
    .b(_0187_),
    .s(N210),
    .y(_0433_)
  );
  al_mux2l _1115_ (
    .a(N595),
    .b(N596),
    .s(N210),
    .y(_0434_)
  );
  al_mux2h _1116_ (
    .a(_0434_),
    .b(_0433_),
    .s(N457),
    .y(_0435_)
  );
  al_aoi21 _1117_ (
    .a(_0153_),
    .b(_0435_),
    .c(N625),
    .y(_0436_)
  );
  al_nand2 _1118_ (
    .a(_0436_),
    .b(_0432_),
    .y(_0437_)
  );
  al_aoi21ftf _1119_ (
    .a(_0162_),
    .b(N114),
    .c(_0437_),
    .y(N7705)
  );
  al_and3ftt _1120_ (
    .a(N619),
    .b(N625),
    .c(N53),
    .y(_0438_)
  );
  al_nand2 _1121_ (
    .a(N422),
    .b(_0239_),
    .y(_0439_)
  );
  al_aoi21ttf _1122_ (
    .a(N4),
    .b(_0415_),
    .c(_0414_),
    .y(_0440_)
  );
  al_aoi21 _1123_ (
    .a(_0439_),
    .b(_0440_),
    .c(_0407_),
    .y(_0441_)
  );
  al_or3fft _1124_ (
    .a(_0427_),
    .b(_0402_),
    .c(_0441_),
    .y(_0442_)
  );
  al_nand2 _1125_ (
    .a(_0406_),
    .b(_0441_),
    .y(_0443_)
  );
  al_nand3 _1126_ (
    .a(N619),
    .b(_0443_),
    .c(_0442_),
    .y(_0444_)
  );
  al_mux2l _1127_ (
    .a(_0188_),
    .b(_0187_),
    .s(N218),
    .y(_0445_)
  );
  al_mux2l _1128_ (
    .a(N595),
    .b(N596),
    .s(N218),
    .y(_0446_)
  );
  al_mux2h _1129_ (
    .a(_0446_),
    .b(_0445_),
    .s(N468),
    .y(_0447_)
  );
  al_aoi21 _1130_ (
    .a(_0153_),
    .b(_0447_),
    .c(N625),
    .y(_0448_)
  );
  al_aoi21 _1131_ (
    .a(_0448_),
    .b(_0444_),
    .c(_0438_),
    .y(N7706)
  );
  al_and2 _1132_ (
    .a(_0408_),
    .b(_0416_),
    .y(_0449_)
  );
  al_nand2ft _1133_ (
    .a(_0408_),
    .b(_0440_),
    .y(_0450_)
  );
  al_nand2ft _1134_ (
    .a(_0449_),
    .b(_0450_),
    .y(_0451_)
  );
  al_inv _1135_ (
    .a(N422),
    .y(_0452_)
  );
  al_mux2l _1136_ (
    .a(N598),
    .b(N597),
    .s(N226),
    .y(_0453_)
  );
  al_mux2l _1137_ (
    .a(_0174_),
    .b(_0175_),
    .s(N226),
    .y(_0454_)
  );
  al_mux2h _1138_ (
    .a(_0453_),
    .b(_0454_),
    .s(_0452_),
    .y(_0455_)
  );
  al_oai21ftf _1139_ (
    .a(_0153_),
    .b(_0455_),
    .c(N625),
    .y(_0456_)
  );
  al_ao21 _1140_ (
    .a(N619),
    .b(_0451_),
    .c(_0456_),
    .y(_0457_)
  );
  al_aoi21ftf _1141_ (
    .a(_0162_),
    .b(N113),
    .c(_0457_),
    .y(N7707)
  );
  al_nand3 _1142_ (
    .a(_0427_),
    .b(_0402_),
    .c(_0419_),
    .y(_0458_)
  );
  al_nand3ftt _1143_ (
    .a(_0396_),
    .b(_0397_),
    .c(_0406_),
    .y(_0459_)
  );
  al_nand2 _1144_ (
    .a(N457),
    .b(_0243_),
    .y(_0460_)
  );
  al_ao21 _1145_ (
    .a(_0460_),
    .b(_0399_),
    .c(_0401_),
    .y(_0461_)
  );
  al_and3ftt _1146_ (
    .a(_0439_),
    .b(_0460_),
    .c(_0399_),
    .y(_0462_)
  );
  al_nand2ft _1147_ (
    .a(_0462_),
    .b(_0461_),
    .y(_0463_)
  );
  al_aoi21ttf _1148_ (
    .a(_0458_),
    .b(_0459_),
    .c(_0463_),
    .y(_0464_)
  );
  al_or3fft _1149_ (
    .a(_0458_),
    .b(_0459_),
    .c(_0463_),
    .y(_0465_)
  );
  al_nand2ft _1150_ (
    .a(_0464_),
    .b(_0465_),
    .y(_0466_)
  );
  al_nand3 _1151_ (
    .a(_0428_),
    .b(_0404_),
    .c(_0409_),
    .y(_0467_)
  );
  al_ao21 _1152_ (
    .a(_0404_),
    .b(_0409_),
    .c(_0428_),
    .y(_0468_)
  );
  al_ao21 _1153_ (
    .a(_0467_),
    .b(_0468_),
    .c(_0466_),
    .y(_0469_)
  );
  al_nand3 _1154_ (
    .a(_0467_),
    .b(_0468_),
    .c(_0466_),
    .y(_0470_)
  );
  al_nand3ftt _1155_ (
    .a(_0414_),
    .b(_0470_),
    .c(_0469_),
    .y(_0471_)
  );
  al_inv _1156_ (
    .a(N566),
    .y(_0472_)
  );
  al_ao21ftf _1157_ (
    .a(_0239_),
    .b(_0452_),
    .c(_0400_),
    .y(_0473_)
  );
  al_nand3fft _1158_ (
    .a(N422),
    .b(_0239_),
    .c(_0427_),
    .y(_0474_)
  );
  al_aoi21ftf _1159_ (
    .a(_0439_),
    .b(_0402_),
    .c(_0474_),
    .y(_0475_)
  );
  al_and3 _1160_ (
    .a(_0473_),
    .b(_0405_),
    .c(_0475_),
    .y(_0476_)
  );
  al_ao21 _1161_ (
    .a(_0473_),
    .b(_0475_),
    .c(_0405_),
    .y(_0477_)
  );
  al_nand2ft _1162_ (
    .a(_0476_),
    .b(_0477_),
    .y(_0478_)
  );
  al_ao21ttf _1163_ (
    .a(_0458_),
    .b(_0459_),
    .c(_0404_),
    .y(_0479_)
  );
  al_or3fft _1164_ (
    .a(_0458_),
    .b(_0459_),
    .c(_0404_),
    .y(_0480_)
  );
  al_or3fft _1165_ (
    .a(_0479_),
    .b(_0480_),
    .c(_0478_),
    .y(_0481_)
  );
  al_ao21ttf _1166_ (
    .a(_0479_),
    .b(_0480_),
    .c(_0478_),
    .y(_0482_)
  );
  al_nand3 _1167_ (
    .a(_0414_),
    .b(_0482_),
    .c(_0481_),
    .y(_0483_)
  );
  al_nand2 _1168_ (
    .a(_0472_),
    .b(_0483_),
    .y(_0484_)
  );
  al_ao21 _1169_ (
    .a(_0308_),
    .b(_0413_),
    .c(_0415_),
    .y(_0485_)
  );
  al_and3ftt _1170_ (
    .a(_0485_),
    .b(_0482_),
    .c(_0481_),
    .y(_0486_)
  );
  al_nand3 _1171_ (
    .a(_0485_),
    .b(_0470_),
    .c(_0469_),
    .y(_0487_)
  );
  al_nand3fft _1172_ (
    .a(_0472_),
    .b(_0486_),
    .c(_0487_),
    .y(_0488_)
  );
  al_ao21ftf _1173_ (
    .a(_0484_),
    .b(_0471_),
    .c(_0488_),
    .y(_0489_)
  );
  al_ao21ftt _1174_ (
    .a(_0315_),
    .b(_0320_),
    .c(_0325_),
    .y(_0490_)
  );
  al_mux2l _1175_ (
    .a(_0310_),
    .b(_0312_),
    .s(_0490_),
    .y(_0491_)
  );
  al_nand2ft _1176_ (
    .a(_0410_),
    .b(_0316_),
    .y(_0492_)
  );
  al_ao21ttf _1177_ (
    .a(_0182_),
    .b(_0183_),
    .c(_0492_),
    .y(_0493_)
  );
  al_nand2ft _1178_ (
    .a(_0320_),
    .b(_0493_),
    .y(_0494_)
  );
  al_mux2h _1179_ (
    .a(_0318_),
    .b(_0316_),
    .s(_0183_),
    .y(_0495_)
  );
  al_nand3ftt _1180_ (
    .a(_0307_),
    .b(_0308_),
    .c(_0495_),
    .y(_0496_)
  );
  al_ao21ftt _1181_ (
    .a(_0307_),
    .b(_0308_),
    .c(_0495_),
    .y(_0497_)
  );
  al_ao21 _1182_ (
    .a(_0496_),
    .b(_0497_),
    .c(_0494_),
    .y(_0498_)
  );
  al_nand3 _1183_ (
    .a(_0496_),
    .b(_0497_),
    .c(_0494_),
    .y(_0499_)
  );
  al_or3fft _1184_ (
    .a(_0499_),
    .b(_0498_),
    .c(_0491_),
    .y(_0500_)
  );
  al_ao21ttf _1185_ (
    .a(_0499_),
    .b(_0498_),
    .c(_0491_),
    .y(_0501_)
  );
  al_nand3 _1186_ (
    .a(N566),
    .b(_0501_),
    .c(_0500_),
    .y(_0502_)
  );
  al_mux2l _1187_ (
    .a(_0318_),
    .b(_0316_),
    .s(_0182_),
    .y(_0503_)
  );
  al_and3ftt _1188_ (
    .a(_0307_),
    .b(_0308_),
    .c(_0503_),
    .y(_0504_)
  );
  al_nand3ftt _1189_ (
    .a(_0319_),
    .b(_0322_),
    .c(_0309_),
    .y(_0505_)
  );
  al_nand2ft _1190_ (
    .a(_0504_),
    .b(_0505_),
    .y(_0506_)
  );
  al_ao21 _1191_ (
    .a(_0313_),
    .b(_0411_),
    .c(_0311_),
    .y(_0507_)
  );
  al_nand3 _1192_ (
    .a(_0412_),
    .b(_0507_),
    .c(_0494_),
    .y(_0508_)
  );
  al_ao21 _1193_ (
    .a(_0412_),
    .b(_0507_),
    .c(_0494_),
    .y(_0509_)
  );
  al_ao21 _1194_ (
    .a(_0508_),
    .b(_0509_),
    .c(_0506_),
    .y(_0510_)
  );
  al_nand3 _1195_ (
    .a(_0506_),
    .b(_0508_),
    .c(_0509_),
    .y(_0511_)
  );
  al_nand3 _1196_ (
    .a(_0472_),
    .b(_0511_),
    .c(_0510_),
    .y(_0512_)
  );
  al_and3ftt _1197_ (
    .a(_0311_),
    .b(_0310_),
    .c(_0315_),
    .y(_0513_)
  );
  al_ao21ftt _1198_ (
    .a(_0311_),
    .b(_0310_),
    .c(_0315_),
    .y(_0514_)
  );
  al_nand2ft _1199_ (
    .a(_0513_),
    .b(_0514_),
    .y(_0515_)
  );
  al_nand3 _1200_ (
    .a(_0515_),
    .b(_0512_),
    .c(_0502_),
    .y(_0516_)
  );
  al_ao21 _1201_ (
    .a(_0512_),
    .b(_0502_),
    .c(_0515_),
    .y(_0517_)
  );
  al_ao21 _1202_ (
    .a(_0517_),
    .b(_0516_),
    .c(_0489_),
    .y(_0518_)
  );
  al_and2 _1203_ (
    .a(_0516_),
    .b(_0517_),
    .y(_0519_)
  );
  al_aoi21 _1204_ (
    .a(_0489_),
    .b(_0519_),
    .c(_0153_),
    .y(_0520_)
  );
  al_mux2l _1205_ (
    .a(N248),
    .b(N251),
    .s(N281),
    .y(_0521_)
  );
  al_mux2l _1206_ (
    .a(_0381_),
    .b(_0382_),
    .s(N281),
    .y(_0522_)
  );
  al_mux2h _1207_ (
    .a(_0521_),
    .b(_0522_),
    .s(_0317_),
    .y(_0523_)
  );
  al_mux2l _1208_ (
    .a(N248),
    .b(N251),
    .s(N234),
    .y(_0524_)
  );
  al_mux2l _1209_ (
    .a(_0381_),
    .b(_0382_),
    .s(N234),
    .y(_0525_)
  );
  al_mux2l _1210_ (
    .a(_0524_),
    .b(_0525_),
    .s(N435),
    .y(_0526_)
  );
  al_nand2 _1211_ (
    .a(_0523_),
    .b(_0526_),
    .y(_0527_)
  );
  al_nor2 _1212_ (
    .a(_0523_),
    .b(_0526_),
    .y(_0528_)
  );
  al_nand2ft _1213_ (
    .a(_0528_),
    .b(_0527_),
    .y(_0529_)
  );
  al_mux2l _1214_ (
    .a(N248),
    .b(N251),
    .s(N273),
    .y(_0530_)
  );
  al_mux2l _1215_ (
    .a(_0381_),
    .b(_0382_),
    .s(N273),
    .y(_0531_)
  );
  al_mux2l _1216_ (
    .a(_0530_),
    .b(_0531_),
    .s(N411),
    .y(_0532_)
  );
  al_mux2l _1217_ (
    .a(N248),
    .b(N251),
    .s(N265),
    .y(_0533_)
  );
  al_mux2l _1218_ (
    .a(_0381_),
    .b(_0382_),
    .s(N265),
    .y(_0534_)
  );
  al_mux2h _1219_ (
    .a(_0533_),
    .b(_0534_),
    .s(_0323_),
    .y(_0535_)
  );
  al_nor2 _1220_ (
    .a(_0535_),
    .b(_0532_),
    .y(_0536_)
  );
  al_nand2 _1221_ (
    .a(_0535_),
    .b(_0532_),
    .y(_0537_)
  );
  al_mux2l _1222_ (
    .a(N248),
    .b(N251),
    .s(N257),
    .y(_0538_)
  );
  al_mux2l _1223_ (
    .a(_0381_),
    .b(_0382_),
    .s(N257),
    .y(_0539_)
  );
  al_mux2l _1224_ (
    .a(_0538_),
    .b(_0539_),
    .s(N389),
    .y(_0540_)
  );
  al_oai21ftt _1225_ (
    .a(_0537_),
    .b(_0536_),
    .c(_0540_),
    .y(_0541_)
  );
  al_and3fft _1226_ (
    .a(_0540_),
    .b(_0536_),
    .c(_0537_),
    .y(_0542_)
  );
  al_aoi21ftt _1227_ (
    .a(_0542_),
    .b(_0541_),
    .c(_0529_),
    .y(_0543_)
  );
  al_nand3ftt _1228_ (
    .a(_0542_),
    .b(_0529_),
    .c(_0541_),
    .y(_0544_)
  );
  al_mux2l _1229_ (
    .a(N248),
    .b(N251),
    .s(N210),
    .y(_0545_)
  );
  al_mux2l _1230_ (
    .a(_0381_),
    .b(_0382_),
    .s(N210),
    .y(_0546_)
  );
  al_mux2l _1231_ (
    .a(_0545_),
    .b(_0546_),
    .s(N457),
    .y(_0547_)
  );
  al_mux2l _1232_ (
    .a(N248),
    .b(N251),
    .s(N226),
    .y(_0548_)
  );
  al_nand2 _1233_ (
    .a(N422),
    .b(_0548_),
    .y(_0549_)
  );
  al_mux2l _1234_ (
    .a(N242),
    .b(N254),
    .s(N226),
    .y(_0550_)
  );
  al_aoi21ftf _1235_ (
    .a(_0550_),
    .b(_0452_),
    .c(_0549_),
    .y(_0551_)
  );
  al_or2ft _1236_ (
    .a(_0551_),
    .b(_0547_),
    .y(_0552_)
  );
  al_and2ft _1237_ (
    .a(_0551_),
    .b(_0547_),
    .y(_0553_)
  );
  al_nand2ft _1238_ (
    .a(_0553_),
    .b(_0552_),
    .y(_0554_)
  );
  al_mux2l _1239_ (
    .a(N248),
    .b(N251),
    .s(N218),
    .y(_0555_)
  );
  al_mux2l _1240_ (
    .a(_0381_),
    .b(_0382_),
    .s(N218),
    .y(_0556_)
  );
  al_mux2l _1241_ (
    .a(_0555_),
    .b(_0556_),
    .s(N468),
    .y(_0557_)
  );
  al_and2ft _1242_ (
    .a(_0424_),
    .b(_0557_),
    .y(_0558_)
  );
  al_nand2ft _1243_ (
    .a(_0557_),
    .b(_0424_),
    .y(_0559_)
  );
  al_aoi21ftf _1244_ (
    .a(_0558_),
    .b(_0559_),
    .c(_0554_),
    .y(_0560_)
  );
  al_or3ftt _1245_ (
    .a(_0559_),
    .b(_0558_),
    .c(_0554_),
    .y(_0561_)
  );
  al_nand2ft _1246_ (
    .a(_0560_),
    .b(_0561_),
    .y(_0562_)
  );
  al_or3ftt _1247_ (
    .a(_0544_),
    .b(_0543_),
    .c(_0562_),
    .y(_0563_)
  );
  al_ao21ftf _1248_ (
    .a(_0543_),
    .b(_0544_),
    .c(_0562_),
    .y(_0564_)
  );
  al_nand3 _1249_ (
    .a(_0153_),
    .b(_0564_),
    .c(_0563_),
    .y(_0565_)
  );
  al_nand2 _1250_ (
    .a(_0158_),
    .b(_0565_),
    .y(_0566_)
  );
  al_ao21 _1251_ (
    .a(_0518_),
    .b(_0520_),
    .c(_0566_),
    .y(_0567_)
  );
  al_nand2 _1252_ (
    .a(N625),
    .b(N97),
    .y(_0568_)
  );
  al_nand3 _1253_ (
    .a(N571),
    .b(_0568_),
    .c(_0567_),
    .y(_0569_)
  );
  al_inv _1254_ (
    .a(N571),
    .y(_0570_)
  );
  al_nand2ft _1255_ (
    .a(_0261_),
    .b(_0269_),
    .y(_0571_)
  );
  al_nand2 _1256_ (
    .a(_0198_),
    .b(_0256_),
    .y(_0572_)
  );
  al_aoi21ttf _1257_ (
    .a(_0198_),
    .b(_0260_),
    .c(_0572_),
    .y(_0573_)
  );
  al_nand3 _1258_ (
    .a(_0199_),
    .b(_0257_),
    .c(_0254_),
    .y(_0574_)
  );
  al_ao21 _1259_ (
    .a(_0257_),
    .b(_0254_),
    .c(_0199_),
    .y(_0575_)
  );
  al_nand3 _1260_ (
    .a(_0255_),
    .b(_0574_),
    .c(_0575_),
    .y(_0576_)
  );
  al_ao21ttf _1261_ (
    .a(_0257_),
    .b(_0254_),
    .c(_0199_),
    .y(_0577_)
  );
  al_nand3ftt _1262_ (
    .a(_0199_),
    .b(_0257_),
    .c(_0254_),
    .y(_0578_)
  );
  al_nand3ftt _1263_ (
    .a(_0255_),
    .b(_0578_),
    .c(_0577_),
    .y(_0579_)
  );
  al_ao21ttf _1264_ (
    .a(_0579_),
    .b(_0576_),
    .c(_0573_),
    .y(_0580_)
  );
  al_or3fft _1265_ (
    .a(_0579_),
    .b(_0576_),
    .c(_0573_),
    .y(_0581_)
  );
  al_nand3 _1266_ (
    .a(_0571_),
    .b(_0580_),
    .c(_0581_),
    .y(_0582_)
  );
  al_inv _1267_ (
    .a(N583),
    .y(_0583_)
  );
  al_nand3ftt _1268_ (
    .a(_0258_),
    .b(_0574_),
    .c(_0575_),
    .y(_0584_)
  );
  al_nand3 _1269_ (
    .a(_0258_),
    .b(_0578_),
    .c(_0577_),
    .y(_0585_)
  );
  al_nand3ftt _1270_ (
    .a(_0572_),
    .b(_0584_),
    .c(_0585_),
    .y(_0586_)
  );
  al_ao21ttf _1271_ (
    .a(_0585_),
    .b(_0584_),
    .c(_0572_),
    .y(_0587_)
  );
  al_nand3 _1272_ (
    .a(_0586_),
    .b(_0587_),
    .c(_0270_),
    .y(_0588_)
  );
  al_nand2 _1273_ (
    .a(_0583_),
    .b(_0588_),
    .y(_0589_)
  );
  al_and3ftt _1274_ (
    .a(_0261_),
    .b(_0275_),
    .c(_0269_),
    .y(_0590_)
  );
  al_and3 _1275_ (
    .a(_0586_),
    .b(_0587_),
    .c(_0590_),
    .y(_0591_)
  );
  al_nand3ftt _1276_ (
    .a(_0590_),
    .b(_0580_),
    .c(_0581_),
    .y(_0592_)
  );
  al_nand3fft _1277_ (
    .a(_0583_),
    .b(_0591_),
    .c(_0592_),
    .y(_0593_)
  );
  al_aoi21ftf _1278_ (
    .a(_0589_),
    .b(_0582_),
    .c(_0593_),
    .y(_0594_)
  );
  al_and2 _1279_ (
    .a(_0265_),
    .b(_0267_),
    .y(_0595_)
  );
  al_ao21ftf _1280_ (
    .a(_0154_),
    .b(_0165_),
    .c(_0166_),
    .y(_0596_)
  );
  al_nand3fft _1281_ (
    .a(_0261_),
    .b(_0262_),
    .c(_0596_),
    .y(_0597_)
  );
  al_oai21ttf _1282_ (
    .a(_0261_),
    .b(_0262_),
    .c(_0596_),
    .y(_0598_)
  );
  al_nand3 _1283_ (
    .a(_0597_),
    .b(_0598_),
    .c(_0595_),
    .y(_0599_)
  );
  al_ao21 _1284_ (
    .a(_0597_),
    .b(_0598_),
    .c(_0595_),
    .y(_0600_)
  );
  al_ao21ttf _1285_ (
    .a(_0600_),
    .b(_0599_),
    .c(_0279_),
    .y(_0601_)
  );
  al_nand3ftt _1286_ (
    .a(_0279_),
    .b(_0600_),
    .c(_0599_),
    .y(_0602_)
  );
  al_nand3 _1287_ (
    .a(_0583_),
    .b(_0602_),
    .c(_0601_),
    .y(_0603_)
  );
  al_aoi21ftf _1288_ (
    .a(_0263_),
    .b(_0268_),
    .c(_0280_),
    .y(_0604_)
  );
  al_mux2h _1289_ (
    .a(_0265_),
    .b(_0266_),
    .s(_0165_),
    .y(_0605_)
  );
  al_oai21ttf _1290_ (
    .a(_0261_),
    .b(_0262_),
    .c(_0605_),
    .y(_0606_)
  );
  al_nand3fft _1291_ (
    .a(_0261_),
    .b(_0262_),
    .c(_0605_),
    .y(_0607_)
  );
  al_ao21 _1292_ (
    .a(_0607_),
    .b(_0606_),
    .c(_0170_),
    .y(_0608_)
  );
  al_nand3 _1293_ (
    .a(_0170_),
    .b(_0606_),
    .c(_0607_),
    .y(_0609_)
  );
  al_ao21ttf _1294_ (
    .a(_0608_),
    .b(_0609_),
    .c(_0604_),
    .y(_0610_)
  );
  al_nand3ftt _1295_ (
    .a(_0604_),
    .b(_0609_),
    .c(_0608_),
    .y(_0611_)
  );
  al_nand3 _1296_ (
    .a(N583),
    .b(_0610_),
    .c(_0611_),
    .y(_0612_)
  );
  al_aoi21 _1297_ (
    .a(_0265_),
    .b(_0266_),
    .c(_0272_),
    .y(_0613_)
  );
  al_nor2ft _1298_ (
    .a(_0273_),
    .b(_0613_),
    .y(_0614_)
  );
  al_ao21 _1299_ (
    .a(_0603_),
    .b(_0612_),
    .c(_0614_),
    .y(_0615_)
  );
  al_nand3 _1300_ (
    .a(_0614_),
    .b(_0603_),
    .c(_0612_),
    .y(_0616_)
  );
  al_ao21 _1301_ (
    .a(_0616_),
    .b(_0615_),
    .c(_0594_),
    .y(_0617_)
  );
  al_nand3 _1302_ (
    .a(_0616_),
    .b(_0615_),
    .c(_0594_),
    .y(_0618_)
  );
  al_nand3 _1303_ (
    .a(N619),
    .b(_0618_),
    .c(_0617_),
    .y(_0619_)
  );
  al_nand2ft _1304_ (
    .a(N514),
    .b(N242),
    .y(_0620_)
  );
  al_ao21ftf _1305_ (
    .a(N248),
    .b(N514),
    .c(_0620_),
    .y(_0621_)
  );
  al_nor2 _1306_ (
    .a(_0159_),
    .b(_0621_),
    .y(_0622_)
  );
  al_nand2 _1307_ (
    .a(_0159_),
    .b(_0621_),
    .y(_0623_)
  );
  al_mux2l _1308_ (
    .a(N248),
    .b(N251),
    .s(N324),
    .y(_0624_)
  );
  al_mux2l _1309_ (
    .a(_0381_),
    .b(_0382_),
    .s(N324),
    .y(_0625_)
  );
  al_mux2l _1310_ (
    .a(_0624_),
    .b(_0625_),
    .s(N503),
    .y(_0626_)
  );
  al_and3ftt _1311_ (
    .a(_0622_),
    .b(_0623_),
    .c(_0626_),
    .y(_0627_)
  );
  al_ao21ftt _1312_ (
    .a(_0622_),
    .b(_0623_),
    .c(_0626_),
    .y(_0628_)
  );
  al_nand2ft _1313_ (
    .a(_0627_),
    .b(_0628_),
    .y(_0629_)
  );
  al_mux2l _1314_ (
    .a(N248),
    .b(N251),
    .s(N351),
    .y(_0630_)
  );
  al_mux2l _1315_ (
    .a(_0381_),
    .b(_0382_),
    .s(N351),
    .y(_0631_)
  );
  al_mux2h _1316_ (
    .a(_0630_),
    .b(_0631_),
    .s(_0172_),
    .y(_0632_)
  );
  al_mux2l _1317_ (
    .a(N248),
    .b(N251),
    .s(N341),
    .y(_0633_)
  );
  al_mux2l _1318_ (
    .a(_0381_),
    .b(_0382_),
    .s(N341),
    .y(_0634_)
  );
  al_mux2l _1319_ (
    .a(_0633_),
    .b(_0634_),
    .s(N523),
    .y(_0635_)
  );
  al_and2ft _1320_ (
    .a(_0632_),
    .b(_0635_),
    .y(_0636_)
  );
  al_nand2ft _1321_ (
    .a(_0635_),
    .b(_0632_),
    .y(_0637_)
  );
  al_ao21ftt _1322_ (
    .a(_0636_),
    .b(_0637_),
    .c(_0629_),
    .y(_0638_)
  );
  al_nand3ftt _1323_ (
    .a(_0636_),
    .b(_0637_),
    .c(_0629_),
    .y(_0639_)
  );
  al_nand2 _1324_ (
    .a(_0384_),
    .b(_0392_),
    .y(_0640_)
  );
  al_or2 _1325_ (
    .a(_0384_),
    .b(_0392_),
    .y(_0641_)
  );
  al_and2ft _1326_ (
    .a(_0367_),
    .b(_0374_),
    .y(_0642_)
  );
  al_nand2ft _1327_ (
    .a(_0374_),
    .b(_0367_),
    .y(_0643_)
  );
  al_nand2ft _1328_ (
    .a(_0642_),
    .b(_0643_),
    .y(_0644_)
  );
  al_ao21 _1329_ (
    .a(_0641_),
    .b(_0640_),
    .c(_0644_),
    .y(_0645_)
  );
  al_and3 _1330_ (
    .a(_0644_),
    .b(_0641_),
    .c(_0640_),
    .y(_0646_)
  );
  al_nand2ft _1331_ (
    .a(_0646_),
    .b(_0645_),
    .y(_0647_)
  );
  al_ao21 _1332_ (
    .a(_0638_),
    .b(_0639_),
    .c(_0647_),
    .y(_0648_)
  );
  al_nand3 _1333_ (
    .a(_0638_),
    .b(_0639_),
    .c(_0647_),
    .y(_0649_)
  );
  al_nand3 _1334_ (
    .a(_0153_),
    .b(_0649_),
    .c(_0648_),
    .y(_0650_)
  );
  al_and2 _1335_ (
    .a(_0158_),
    .b(_0650_),
    .y(_0651_)
  );
  al_and2 _1336_ (
    .a(N625),
    .b(N94),
    .y(_0652_)
  );
  al_aoi21 _1337_ (
    .a(_0651_),
    .b(_0619_),
    .c(_0652_),
    .y(_0653_)
  );
  al_aoi21 _1338_ (
    .a(_0570_),
    .b(_0653_),
    .c(N574),
    .y(_0654_)
  );
  al_and2ft _1339_ (
    .a(N571),
    .b(N574),
    .y(_0655_)
  );
  al_and3 _1340_ (
    .a(N571),
    .b(N574),
    .c(N179),
    .y(_0656_)
  );
  al_ao21 _1341_ (
    .a(N176),
    .b(_0655_),
    .c(_0656_),
    .y(_0657_)
  );
  al_ao21 _1342_ (
    .a(_0654_),
    .b(_0569_),
    .c(_0657_),
    .y(_0658_)
  );
  al_nand2 _1343_ (
    .a(N137),
    .b(_0658_),
    .y(N8127)
  );
  al_nand3 _1344_ (
    .a(N577),
    .b(_0568_),
    .c(_0567_),
    .y(_0659_)
  );
  al_inv _1345_ (
    .a(N577),
    .y(_0660_)
  );
  al_aoi21 _1346_ (
    .a(_0660_),
    .b(_0653_),
    .c(N580),
    .y(_0661_)
  );
  al_and2ft _1347_ (
    .a(N577),
    .b(N580),
    .y(_0662_)
  );
  al_and3 _1348_ (
    .a(N577),
    .b(N580),
    .c(N179),
    .y(_0663_)
  );
  al_ao21 _1349_ (
    .a(N176),
    .b(_0662_),
    .c(_0663_),
    .y(_0664_)
  );
  al_ao21 _1350_ (
    .a(_0661_),
    .b(_0659_),
    .c(_0664_),
    .y(_0665_)
  );
  al_nand2 _1351_ (
    .a(N137),
    .b(_0665_),
    .y(N8128)
  );
  al_and2 _1352_ (
    .a(N552),
    .b(N562),
    .y(N1140)
  );
  al_and2 _1353_ (
    .a(N373),
    .b(N1),
    .y(N1972)
  );
  al_and2 _1354_ (
    .a(N141),
    .b(N145),
    .y(N1147)
  );
  al_and2ft _1355_ (
    .a(N592),
    .b(N136),
    .y(N2054)
  );
  al_inv _1356_ (
    .a(N141),
    .y(_0666_)
  );
  al_nand2 _1357_ (
    .a(N588),
    .b(N25),
    .y(_0667_)
  );
  al_aoi21ftf _1358_ (
    .a(N588),
    .b(N24),
    .c(_0108_),
    .y(_0668_)
  );
  al_aoi21 _1359_ (
    .a(_0667_),
    .b(_0668_),
    .c(_0666_),
    .y(N4737)
  );
  al_nand2 _1360_ (
    .a(N588),
    .b(N81),
    .y(_0669_)
  );
  al_aoi21ftf _1361_ (
    .a(N588),
    .b(N26),
    .c(_0108_),
    .y(_0670_)
  );
  al_aoi21 _1362_ (
    .a(_0669_),
    .b(_0670_),
    .c(_0666_),
    .y(N4738)
  );
  al_nand2 _1363_ (
    .a(N588),
    .b(N23),
    .y(_0671_)
  );
  al_aoi21ftf _1364_ (
    .a(N588),
    .b(N79),
    .c(_0108_),
    .y(_0672_)
  );
  al_aoi21 _1365_ (
    .a(_0671_),
    .b(_0672_),
    .c(_0666_),
    .y(N4739)
  );
  al_nand2 _1366_ (
    .a(N588),
    .b(N80),
    .y(_0673_)
  );
  al_aoi21ftf _1367_ (
    .a(N588),
    .b(N82),
    .c(_0108_),
    .y(_0674_)
  );
  al_aoi21 _1368_ (
    .a(_0673_),
    .b(_0674_),
    .c(_0666_),
    .y(N4740)
  );
  al_nand2ft _1369_ (
    .a(_0177_),
    .b(_0287_),
    .y(_0675_)
  );
  al_and2 _1370_ (
    .a(_0159_),
    .b(_0295_),
    .y(_0676_)
  );
  al_and3 _1371_ (
    .a(_0642_),
    .b(_0676_),
    .c(_0304_),
    .y(_0677_)
  );
  al_nor3ftt _1372_ (
    .a(_0677_),
    .b(_0675_),
    .c(_0640_),
    .y(N5240)
  );
  al_and3ftt _1373_ (
    .a(_0455_),
    .b(_0435_),
    .c(_0447_),
    .y(_0678_)
  );
  al_and2 _1374_ (
    .a(_0191_),
    .b(_0333_),
    .y(_0679_)
  );
  al_and2 _1375_ (
    .a(_0362_),
    .b(_0424_),
    .y(_0680_)
  );
  al_and3 _1376_ (
    .a(_0342_),
    .b(_0353_),
    .c(_0680_),
    .y(_0681_)
  );
  al_and3 _1377_ (
    .a(_0678_),
    .b(_0679_),
    .c(_0681_),
    .y(N5388)
  );
  al_and3fft _1378_ (
    .a(_0419_),
    .b(_0409_),
    .c(_0415_),
    .y(N6641)
  );
  al_and3fft _1379_ (
    .a(_0200_),
    .b(_0275_),
    .c(_0260_),
    .y(N6643)
  );
  al_and3fft _1380_ (
    .a(_0396_),
    .b(_0409_),
    .c(_0397_),
    .y(_0682_)
  );
  al_oai21ftf _1381_ (
    .a(_0397_),
    .b(_0404_),
    .c(_0396_),
    .y(_0683_)
  );
  al_oai21ftf _1382_ (
    .a(_0682_),
    .b(_0414_),
    .c(_0683_),
    .y(N6924)
  );
  al_or3 _1383_ (
    .a(_0198_),
    .b(_0199_),
    .c(_0256_),
    .y(_0684_)
  );
  al_ao21 _1384_ (
    .a(_0260_),
    .b(_0571_),
    .c(_0684_),
    .y(N6925)
  );
  al_inv _1385_ (
    .a(N610),
    .y(_0685_)
  );
  al_ao21 _1386_ (
    .a(_0685_),
    .b(N7015),
    .c(N607),
    .y(_0686_)
  );
  al_ao21 _1387_ (
    .a(N610),
    .b(N7365),
    .c(_0686_),
    .y(_0687_)
  );
  al_and2ft _1388_ (
    .a(N610),
    .b(N607),
    .y(_0688_)
  );
  al_and3 _1389_ (
    .a(N610),
    .b(N607),
    .c(N61),
    .y(_0689_)
  );
  al_aoi21 _1390_ (
    .a(N11),
    .b(_0688_),
    .c(_0689_),
    .y(_0690_)
  );
  al_nand2 _1391_ (
    .a(_0690_),
    .b(_0687_),
    .y(N7449)
  );
  al_inv _1392_ (
    .a(N613),
    .y(_0691_)
  );
  al_ao21 _1393_ (
    .a(_0691_),
    .b(N7015),
    .c(N616),
    .y(_0692_)
  );
  al_ao21 _1394_ (
    .a(N613),
    .b(N7365),
    .c(_0692_),
    .y(_0693_)
  );
  al_and3 _1395_ (
    .a(N613),
    .b(N616),
    .c(N61),
    .y(_0694_)
  );
  al_and2ft _1396_ (
    .a(N613),
    .b(N616),
    .y(_0695_)
  );
  al_aoi21 _1397_ (
    .a(N11),
    .b(_0695_),
    .c(_0694_),
    .y(_0696_)
  );
  al_nand2 _1398_ (
    .a(_0696_),
    .b(_0693_),
    .y(N7469)
  );
  al_and2 _1399_ (
    .a(_0443_),
    .b(_0442_),
    .y(_0697_)
  );
  al_nand3 _1400_ (
    .a(_0350_),
    .b(_0359_),
    .c(_0339_),
    .y(_0698_)
  );
  al_and3ftt _1401_ (
    .a(_0698_),
    .b(_0330_),
    .c(_0451_),
    .y(_0699_)
  );
  al_and3 _1402_ (
    .a(_0418_),
    .b(_0420_),
    .c(_0699_),
    .y(_0700_)
  );
  al_and3 _1403_ (
    .a(_0186_),
    .b(_0431_),
    .c(_0430_),
    .y(_0701_)
  );
  al_and3 _1404_ (
    .a(_0697_),
    .b(_0701_),
    .c(_0700_),
    .y(N7503)
  );
  al_aoi21ftt _1405_ (
    .a(_0156_),
    .b(_0155_),
    .c(_0167_),
    .y(_0702_)
  );
  al_and3 _1406_ (
    .a(_0301_),
    .b(_0702_),
    .c(_0294_),
    .y(_0703_)
  );
  al_and3 _1407_ (
    .a(_0284_),
    .b(_0703_),
    .c(_0389_),
    .y(_0704_)
  );
  al_and3ftt _1408_ (
    .a(_0371_),
    .b(_0372_),
    .c(_0704_),
    .y(_0705_)
  );
  al_and3 _1409_ (
    .a(N7432),
    .b(_0379_),
    .c(_0705_),
    .y(N7504)
  );
  al_inv _1410_ (
    .a(N137),
    .y(_0706_)
  );
  al_ao21 _1411_ (
    .a(_0570_),
    .b(N7015),
    .c(N574),
    .y(_0707_)
  );
  al_ao21 _1412_ (
    .a(N571),
    .b(N7365),
    .c(_0707_),
    .y(_0708_)
  );
  al_and3 _1413_ (
    .a(N571),
    .b(N574),
    .c(N185),
    .y(_0709_)
  );
  al_aoi21 _1414_ (
    .a(N182),
    .b(_0655_),
    .c(_0709_),
    .y(_0710_)
  );
  al_aoi21 _1415_ (
    .a(_0710_),
    .b(_0708_),
    .c(_0706_),
    .y(N7506)
  );
  al_ao21 _1416_ (
    .a(_0660_),
    .b(N7015),
    .c(N580),
    .y(_0711_)
  );
  al_ao21 _1417_ (
    .a(N577),
    .b(N7365),
    .c(_0711_),
    .y(_0712_)
  );
  al_and3 _1418_ (
    .a(N577),
    .b(N580),
    .c(N185),
    .y(_0713_)
  );
  al_aoi21 _1419_ (
    .a(N182),
    .b(_0662_),
    .c(_0713_),
    .y(_0714_)
  );
  al_aoi21 _1420_ (
    .a(_0714_),
    .b(_0712_),
    .c(_0706_),
    .y(N7511)
  );
  al_inv _1421_ (
    .a(N607),
    .y(_0715_)
  );
  al_mux2h _1422_ (
    .a(N7465),
    .b(N7470),
    .s(N610),
    .y(_0716_)
  );
  al_and3 _1423_ (
    .a(N610),
    .b(N607),
    .c(N37),
    .y(_0717_)
  );
  al_ao21 _1424_ (
    .a(N43),
    .b(_0688_),
    .c(_0717_),
    .y(_0718_)
  );
  al_oai21ftf _1425_ (
    .a(_0715_),
    .b(_0716_),
    .c(_0718_),
    .y(N7515)
  );
  al_mux2h _1426_ (
    .a(_0298_),
    .b(_0345_),
    .s(N610),
    .y(_0719_)
  );
  al_and3 _1427_ (
    .a(N610),
    .b(N607),
    .c(N20),
    .y(_0720_)
  );
  al_ao21 _1428_ (
    .a(N76),
    .b(_0688_),
    .c(_0720_),
    .y(_0721_)
  );
  al_ao21 _1429_ (
    .a(_0715_),
    .b(_0719_),
    .c(_0721_),
    .y(N7516)
  );
  al_nand2 _1430_ (
    .a(N610),
    .b(N7472),
    .y(_0722_)
  );
  al_aoi21 _1431_ (
    .a(_0685_),
    .b(N7467),
    .c(N607),
    .y(_0723_)
  );
  al_and3 _1432_ (
    .a(N610),
    .b(N607),
    .c(N17),
    .y(_0724_)
  );
  al_ao21 _1433_ (
    .a(N73),
    .b(_0688_),
    .c(_0724_),
    .y(_0725_)
  );
  al_ao21 _1434_ (
    .a(_0723_),
    .b(_0722_),
    .c(_0725_),
    .y(N7517)
  );
  al_mux2h _1435_ (
    .a(_0365_),
    .b(_0180_),
    .s(_0685_),
    .y(_0726_)
  );
  al_and3 _1436_ (
    .a(N610),
    .b(N607),
    .c(N70),
    .y(_0727_)
  );
  al_ao21 _1437_ (
    .a(N67),
    .b(_0688_),
    .c(_0727_),
    .y(_0728_)
  );
  al_ao21 _1438_ (
    .a(_0715_),
    .b(_0726_),
    .c(_0728_),
    .y(N7518)
  );
  al_inv _1439_ (
    .a(N616),
    .y(_0729_)
  );
  al_mux2h _1440_ (
    .a(N7465),
    .b(N7470),
    .s(N613),
    .y(_0730_)
  );
  al_and3 _1441_ (
    .a(N613),
    .b(N616),
    .c(N37),
    .y(_0731_)
  );
  al_ao21 _1442_ (
    .a(N43),
    .b(_0695_),
    .c(_0731_),
    .y(_0732_)
  );
  al_oai21ftf _1443_ (
    .a(_0729_),
    .b(_0730_),
    .c(_0732_),
    .y(N7519)
  );
  al_mux2h _1444_ (
    .a(_0298_),
    .b(_0345_),
    .s(N613),
    .y(_0733_)
  );
  al_and3 _1445_ (
    .a(N613),
    .b(N616),
    .c(N20),
    .y(_0734_)
  );
  al_ao21 _1446_ (
    .a(N76),
    .b(_0695_),
    .c(_0734_),
    .y(_0735_)
  );
  al_ao21 _1447_ (
    .a(_0729_),
    .b(_0733_),
    .c(_0735_),
    .y(N7520)
  );
  al_nand2 _1448_ (
    .a(N613),
    .b(N7472),
    .y(_0736_)
  );
  al_aoi21 _1449_ (
    .a(_0691_),
    .b(N7467),
    .c(N616),
    .y(_0737_)
  );
  al_and3 _1450_ (
    .a(N613),
    .b(N616),
    .c(N17),
    .y(_0738_)
  );
  al_ao21 _1451_ (
    .a(N73),
    .b(_0695_),
    .c(_0738_),
    .y(_0739_)
  );
  al_ao21 _1452_ (
    .a(_0737_),
    .b(_0736_),
    .c(_0739_),
    .y(N7521)
  );
  al_mux2h _1453_ (
    .a(_0365_),
    .b(_0180_),
    .s(_0691_),
    .y(_0740_)
  );
  al_and3 _1454_ (
    .a(N613),
    .b(N616),
    .c(N70),
    .y(_0741_)
  );
  al_ao21 _1455_ (
    .a(N67),
    .b(_0695_),
    .c(_0741_),
    .y(_0742_)
  );
  al_ao21 _1456_ (
    .a(_0729_),
    .b(_0740_),
    .c(_0742_),
    .y(N7522)
  );
  al_ao21 _1457_ (
    .a(_0570_),
    .b(N7465),
    .c(N574),
    .y(_0743_)
  );
  al_ao21 _1458_ (
    .a(N571),
    .b(N7470),
    .c(_0743_),
    .y(_0744_)
  );
  al_and3 _1459_ (
    .a(N571),
    .b(N574),
    .c(N170),
    .y(_0745_)
  );
  al_aoi21 _1460_ (
    .a(N200),
    .b(_0655_),
    .c(_0745_),
    .y(_0746_)
  );
  al_aoi21 _1461_ (
    .a(_0746_),
    .b(_0744_),
    .c(_0706_),
    .y(N7600)
  );
  al_inv _1462_ (
    .a(N574),
    .y(_0747_)
  );
  al_mux2h _1463_ (
    .a(_0365_),
    .b(_0180_),
    .s(_0570_),
    .y(_0748_)
  );
  al_nand2 _1464_ (
    .a(_0747_),
    .b(_0748_),
    .y(_0749_)
  );
  al_and3 _1465_ (
    .a(N571),
    .b(N574),
    .c(N158),
    .y(_0750_)
  );
  al_aoi21 _1466_ (
    .a(N188),
    .b(_0655_),
    .c(_0750_),
    .y(_0000_)
  );
  al_aoi21 _1467_ (
    .a(_0000_),
    .b(_0749_),
    .c(_0706_),
    .y(N7601)
  );
  al_aoi21 _1468_ (
    .a(_0570_),
    .b(N7467),
    .c(N574),
    .y(_0001_)
  );
  al_ao21ftf _1469_ (
    .a(_0570_),
    .b(N7472),
    .c(_0001_),
    .y(_0002_)
  );
  al_and3 _1470_ (
    .a(N571),
    .b(N574),
    .c(N152),
    .y(_0003_)
  );
  al_aoi21 _1471_ (
    .a(N155),
    .b(_0655_),
    .c(_0003_),
    .y(_0004_)
  );
  al_aoi21 _1472_ (
    .a(_0004_),
    .b(_0002_),
    .c(_0706_),
    .y(N7602)
  );
  al_mux2h _1473_ (
    .a(_0298_),
    .b(_0345_),
    .s(N571),
    .y(_0005_)
  );
  al_nand2 _1474_ (
    .a(_0747_),
    .b(_0005_),
    .y(_0006_)
  );
  al_and3 _1475_ (
    .a(N571),
    .b(N574),
    .c(N146),
    .y(_0007_)
  );
  al_aoi21 _1476_ (
    .a(N149),
    .b(_0655_),
    .c(_0007_),
    .y(_0008_)
  );
  al_aoi21 _1477_ (
    .a(_0008_),
    .b(_0006_),
    .c(_0706_),
    .y(N7603)
  );
  al_ao21 _1478_ (
    .a(_0660_),
    .b(N7465),
    .c(N580),
    .y(_0009_)
  );
  al_ao21 _1479_ (
    .a(N577),
    .b(N7470),
    .c(_0009_),
    .y(_0010_)
  );
  al_and3 _1480_ (
    .a(N577),
    .b(N580),
    .c(N170),
    .y(_0011_)
  );
  al_aoi21 _1481_ (
    .a(N200),
    .b(_0662_),
    .c(_0011_),
    .y(_0012_)
  );
  al_aoi21 _1482_ (
    .a(_0012_),
    .b(_0010_),
    .c(_0706_),
    .y(N7604)
  );
  al_inv _1483_ (
    .a(N580),
    .y(_0013_)
  );
  al_mux2h _1484_ (
    .a(_0365_),
    .b(_0180_),
    .s(_0660_),
    .y(_0014_)
  );
  al_nand2 _1485_ (
    .a(_0013_),
    .b(_0014_),
    .y(_0015_)
  );
  al_and3 _1486_ (
    .a(N577),
    .b(N580),
    .c(N158),
    .y(_0016_)
  );
  al_aoi21 _1487_ (
    .a(N188),
    .b(_0662_),
    .c(_0016_),
    .y(_0017_)
  );
  al_aoi21 _1488_ (
    .a(_0017_),
    .b(_0015_),
    .c(_0706_),
    .y(N7605)
  );
  al_aoi21 _1489_ (
    .a(_0660_),
    .b(N7467),
    .c(N580),
    .y(_0018_)
  );
  al_ao21ftf _1490_ (
    .a(_0660_),
    .b(N7472),
    .c(_0018_),
    .y(_0019_)
  );
  al_and3 _1491_ (
    .a(N577),
    .b(N580),
    .c(N152),
    .y(_0020_)
  );
  al_aoi21 _1492_ (
    .a(N155),
    .b(_0662_),
    .c(_0020_),
    .y(_0021_)
  );
  al_aoi21 _1493_ (
    .a(_0021_),
    .b(_0019_),
    .c(_0706_),
    .y(N7606)
  );
  al_mux2h _1494_ (
    .a(_0298_),
    .b(_0345_),
    .s(N577),
    .y(_0022_)
  );
  al_nand2 _1495_ (
    .a(_0013_),
    .b(_0022_),
    .y(_0023_)
  );
  al_and3 _1496_ (
    .a(N577),
    .b(N580),
    .c(N146),
    .y(_0024_)
  );
  al_aoi21 _1497_ (
    .a(N149),
    .b(_0662_),
    .c(_0024_),
    .y(_0025_)
  );
  al_aoi21 _1498_ (
    .a(_0025_),
    .b(_0023_),
    .c(_0706_),
    .y(N7607)
  );
  al_and2 _1499_ (
    .a(N135),
    .b(N631),
    .y(_0026_)
  );
  al_and2ft _1500_ (
    .a(N132),
    .b(_0199_),
    .y(_0027_)
  );
  al_or2ft _1501_ (
    .a(N132),
    .b(_0199_),
    .y(_0028_)
  );
  al_nand2ft _1502_ (
    .a(_0027_),
    .b(_0028_),
    .y(_0029_)
  );
  al_oai21ttf _1503_ (
    .a(N603),
    .b(_0367_),
    .c(N599),
    .y(_0030_)
  );
  al_ao21 _1504_ (
    .a(N603),
    .b(_0029_),
    .c(_0030_),
    .y(_0031_)
  );
  al_oa21 _1505_ (
    .a(N603),
    .b(N123),
    .c(N599),
    .y(_0032_)
  );
  al_ao21ttf _1506_ (
    .a(N603),
    .b(N7432),
    .c(_0032_),
    .y(_0033_)
  );
  al_aoi21 _1507_ (
    .a(_0031_),
    .b(_0033_),
    .c(_0026_),
    .y(N7626)
  );
  al_and2 _1508_ (
    .a(_0029_),
    .b(N7432),
    .y(_0034_)
  );
  al_or3ftt _1509_ (
    .a(_0028_),
    .b(_0027_),
    .c(N7432),
    .y(_0035_)
  );
  al_and2ft _1510_ (
    .a(_0034_),
    .b(_0035_),
    .y(N7698)
  );
  al_nand3 _1511_ (
    .a(N552),
    .b(N562),
    .c(N559),
    .y(_0036_)
  );
  al_nor3ftt _1512_ (
    .a(N245),
    .b(_0036_),
    .c(N2061),
    .y(_0037_)
  );
  al_and3fft _1513_ (
    .a(N6716),
    .b(N6877),
    .c(_0037_),
    .y(_0038_)
  );
  al_and3fft _1514_ (
    .a(N7474),
    .b(N7476),
    .c(_0038_),
    .y(N7703)
  );
  al_nand3fft _1515_ (
    .a(N613),
    .b(_0366_),
    .c(_0369_),
    .y(_0039_)
  );
  al_aoi21 _1516_ (
    .a(N613),
    .b(N7704),
    .c(N616),
    .y(_0040_)
  );
  al_and3 _1517_ (
    .a(N613),
    .b(N616),
    .c(N106),
    .y(_0041_)
  );
  al_ao21 _1518_ (
    .a(N109),
    .b(_0695_),
    .c(_0041_),
    .y(_0042_)
  );
  al_ao21 _1519_ (
    .a(_0039_),
    .b(_0040_),
    .c(_0042_),
    .y(N7735)
  );
  al_nand3fft _1520_ (
    .a(N610),
    .b(_0366_),
    .c(_0369_),
    .y(_0043_)
  );
  al_aoi21 _1521_ (
    .a(N610),
    .b(N7704),
    .c(N607),
    .y(_0044_)
  );
  al_and3 _1522_ (
    .a(N610),
    .b(N607),
    .c(N106),
    .y(_0045_)
  );
  al_ao21 _1523_ (
    .a(N109),
    .b(_0688_),
    .c(_0045_),
    .y(_0046_)
  );
  al_ao21 _1524_ (
    .a(_0043_),
    .b(_0044_),
    .c(_0046_),
    .y(N7736)
  );
  al_mux2h _1525_ (
    .a(N7700),
    .b(N7705),
    .s(N610),
    .y(_0047_)
  );
  al_and3 _1526_ (
    .a(N610),
    .b(N607),
    .c(N49),
    .y(_0048_)
  );
  al_ao21 _1527_ (
    .a(N46),
    .b(_0688_),
    .c(_0048_),
    .y(_0049_)
  );
  al_oai21ftf _1528_ (
    .a(_0715_),
    .b(_0047_),
    .c(_0049_),
    .y(N7737)
  );
  al_mux2h _1529_ (
    .a(N7706),
    .b(N7701),
    .s(_0685_),
    .y(_0050_)
  );
  al_and3 _1530_ (
    .a(N610),
    .b(N607),
    .c(N103),
    .y(_0051_)
  );
  al_ao21 _1531_ (
    .a(N100),
    .b(_0688_),
    .c(_0051_),
    .y(_0052_)
  );
  al_oai21ftf _1532_ (
    .a(_0715_),
    .b(_0050_),
    .c(_0052_),
    .y(N7738)
  );
  al_nand2 _1533_ (
    .a(N610),
    .b(N7707),
    .y(_0053_)
  );
  al_aoi21 _1534_ (
    .a(_0685_),
    .b(N7702),
    .c(N607),
    .y(_0054_)
  );
  al_and3 _1535_ (
    .a(N610),
    .b(N607),
    .c(N40),
    .y(_0055_)
  );
  al_ao21 _1536_ (
    .a(N91),
    .b(_0688_),
    .c(_0055_),
    .y(_0056_)
  );
  al_ao21 _1537_ (
    .a(_0053_),
    .b(_0054_),
    .c(_0056_),
    .y(N7739)
  );
  al_mux2h _1538_ (
    .a(N7700),
    .b(N7705),
    .s(N613),
    .y(_0057_)
  );
  al_and3 _1539_ (
    .a(N613),
    .b(N616),
    .c(N49),
    .y(_0058_)
  );
  al_ao21 _1540_ (
    .a(N46),
    .b(_0695_),
    .c(_0058_),
    .y(_0059_)
  );
  al_oai21ftf _1541_ (
    .a(_0729_),
    .b(_0057_),
    .c(_0059_),
    .y(N7740)
  );
  al_mux2h _1542_ (
    .a(N7706),
    .b(N7701),
    .s(_0691_),
    .y(_0060_)
  );
  al_and3 _1543_ (
    .a(N613),
    .b(N616),
    .c(N103),
    .y(_0061_)
  );
  al_ao21 _1544_ (
    .a(N100),
    .b(_0695_),
    .c(_0061_),
    .y(_0062_)
  );
  al_oai21ftf _1545_ (
    .a(_0729_),
    .b(_0060_),
    .c(_0062_),
    .y(N7741)
  );
  al_nand2 _1546_ (
    .a(N613),
    .b(N7707),
    .y(_0063_)
  );
  al_aoi21 _1547_ (
    .a(_0691_),
    .b(N7702),
    .c(N616),
    .y(_0064_)
  );
  al_and3 _1548_ (
    .a(N613),
    .b(N616),
    .c(N40),
    .y(_0065_)
  );
  al_ao21 _1549_ (
    .a(N91),
    .b(_0695_),
    .c(_0065_),
    .y(_0066_)
  );
  al_ao21 _1550_ (
    .a(_0063_),
    .b(_0064_),
    .c(_0066_),
    .y(N7742)
  );
  al_aoi21 _1551_ (
    .a(_0570_),
    .b(N7702),
    .c(N574),
    .y(_0067_)
  );
  al_ao21ftf _1552_ (
    .a(_0570_),
    .b(N7707),
    .c(_0067_),
    .y(_0068_)
  );
  al_and3 _1553_ (
    .a(N571),
    .b(N574),
    .c(N173),
    .y(_0069_)
  );
  al_aoi21 _1554_ (
    .a(N203),
    .b(_0655_),
    .c(_0069_),
    .y(_0070_)
  );
  al_aoi21 _1555_ (
    .a(_0070_),
    .b(_0068_),
    .c(_0706_),
    .y(N7754)
  );
  al_aoi21 _1556_ (
    .a(N571),
    .b(N7706),
    .c(N574),
    .y(_0071_)
  );
  al_ao21ttf _1557_ (
    .a(_0570_),
    .b(N7701),
    .c(_0071_),
    .y(_0072_)
  );
  al_and3 _1558_ (
    .a(N571),
    .b(N574),
    .c(N167),
    .y(_0073_)
  );
  al_aoi21 _1559_ (
    .a(N197),
    .b(_0655_),
    .c(_0073_),
    .y(_0074_)
  );
  al_aoi21 _1560_ (
    .a(_0074_),
    .b(_0072_),
    .c(_0706_),
    .y(N7755)
  );
  al_aoi21 _1561_ (
    .a(_0570_),
    .b(N7700),
    .c(N574),
    .y(_0075_)
  );
  al_ao21ftf _1562_ (
    .a(_0570_),
    .b(N7705),
    .c(_0075_),
    .y(_0076_)
  );
  al_and3 _1563_ (
    .a(N571),
    .b(N574),
    .c(N164),
    .y(_0077_)
  );
  al_aoi21 _1564_ (
    .a(N194),
    .b(_0655_),
    .c(_0077_),
    .y(_0078_)
  );
  al_aoi21 _1565_ (
    .a(_0078_),
    .b(_0076_),
    .c(_0706_),
    .y(N7756)
  );
  al_aoi21 _1566_ (
    .a(N571),
    .b(N7704),
    .c(N574),
    .y(_0079_)
  );
  al_ao21ftf _1567_ (
    .a(N571),
    .b(N7699),
    .c(_0079_),
    .y(_0080_)
  );
  al_and3 _1568_ (
    .a(N571),
    .b(N574),
    .c(N161),
    .y(_0081_)
  );
  al_aoi21 _1569_ (
    .a(N191),
    .b(_0655_),
    .c(_0081_),
    .y(_0082_)
  );
  al_aoi21 _1570_ (
    .a(_0082_),
    .b(_0080_),
    .c(_0706_),
    .y(N7757)
  );
  al_aoi21 _1571_ (
    .a(_0660_),
    .b(N7702),
    .c(N580),
    .y(_0083_)
  );
  al_ao21ftf _1572_ (
    .a(_0660_),
    .b(N7707),
    .c(_0083_),
    .y(_0084_)
  );
  al_and3 _1573_ (
    .a(N577),
    .b(N580),
    .c(N173),
    .y(_0085_)
  );
  al_aoi21 _1574_ (
    .a(N203),
    .b(_0662_),
    .c(_0085_),
    .y(_0086_)
  );
  al_aoi21 _1575_ (
    .a(_0086_),
    .b(_0084_),
    .c(_0706_),
    .y(N7758)
  );
  al_aoi21 _1576_ (
    .a(N577),
    .b(N7706),
    .c(N580),
    .y(_0087_)
  );
  al_ao21ttf _1577_ (
    .a(_0660_),
    .b(N7701),
    .c(_0087_),
    .y(_0088_)
  );
  al_and3 _1578_ (
    .a(N577),
    .b(N580),
    .c(N167),
    .y(_0089_)
  );
  al_aoi21 _1579_ (
    .a(N197),
    .b(_0662_),
    .c(_0089_),
    .y(_0090_)
  );
  al_aoi21 _1580_ (
    .a(_0090_),
    .b(_0088_),
    .c(_0706_),
    .y(N7759)
  );
  al_aoi21 _1581_ (
    .a(_0660_),
    .b(N7700),
    .c(N580),
    .y(_0091_)
  );
  al_ao21ftf _1582_ (
    .a(_0660_),
    .b(N7705),
    .c(_0091_),
    .y(_0092_)
  );
  al_and3 _1583_ (
    .a(N577),
    .b(N580),
    .c(N164),
    .y(_0093_)
  );
  al_aoi21 _1584_ (
    .a(N194),
    .b(_0662_),
    .c(_0093_),
    .y(_0094_)
  );
  al_aoi21 _1585_ (
    .a(_0094_),
    .b(_0092_),
    .c(_0706_),
    .y(N7760)
  );
  al_aoi21 _1586_ (
    .a(N577),
    .b(N7704),
    .c(N580),
    .y(_0095_)
  );
  al_ao21ftf _1587_ (
    .a(N577),
    .b(N7699),
    .c(_0095_),
    .y(_0096_)
  );
  al_and3 _1588_ (
    .a(N577),
    .b(N580),
    .c(N161),
    .y(_0097_)
  );
  al_aoi21 _1589_ (
    .a(N191),
    .b(_0662_),
    .c(_0097_),
    .y(_0098_)
  );
  al_aoi21 _1590_ (
    .a(_0098_),
    .b(_0096_),
    .c(_0706_),
    .y(N7761)
  );
  al_and3fft _1591_ (
    .a(N619),
    .b(N120),
    .c(N625),
    .y(_0099_)
  );
  al_aoi21 _1592_ (
    .a(_0651_),
    .b(_0619_),
    .c(_0099_),
    .y(N8075)
  );
  al_aoi21ftf _1593_ (
    .a(N118),
    .b(_0161_),
    .c(_0567_),
    .y(N8076)
  );
  al_nand3 _1594_ (
    .a(N610),
    .b(_0568_),
    .c(_0567_),
    .y(_0100_)
  );
  al_aoi21 _1595_ (
    .a(_0685_),
    .b(_0653_),
    .c(N607),
    .y(_0101_)
  );
  al_and3 _1596_ (
    .a(N610),
    .b(N607),
    .c(N64),
    .y(_0102_)
  );
  al_ao21 _1597_ (
    .a(N14),
    .b(_0688_),
    .c(_0102_),
    .y(_0103_)
  );
  al_ao21 _1598_ (
    .a(_0101_),
    .b(_0100_),
    .c(_0103_),
    .y(N8123)
  );
  al_nand3 _1599_ (
    .a(N613),
    .b(_0568_),
    .c(_0567_),
    .y(_0104_)
  );
  al_aoi21 _1600_ (
    .a(_0691_),
    .b(_0653_),
    .c(N616),
    .y(_0105_)
  );
  al_and3 _1601_ (
    .a(N613),
    .b(N616),
    .c(N64),
    .y(_0106_)
  );
  al_ao21 _1602_ (
    .a(N14),
    .b(_0695_),
    .c(_0106_),
    .y(_0107_)
  );
  al_ao21 _1603_ (
    .a(_0105_),
    .b(_0104_),
    .c(_0107_),
    .y(N8124)
  );
  al_and3fft _1604_ (
    .a(_0200_),
    .b(_0275_),
    .c(_0260_),
    .y(N6646)
  );
  al_and3fft _1605_ (
    .a(_0419_),
    .b(_0409_),
    .c(_0415_),
    .y(N6648)
  );
  al_oai21ftf _1606_ (
    .a(_0682_),
    .b(_0414_),
    .c(_0683_),
    .y(N6926)
  );
  al_ao21 _1607_ (
    .a(_0260_),
    .b(_0571_),
    .c(_0684_),
    .y(N6927)
  );
  assign N1066 = N592;
  assign N1142 = N1137;
  assign N1143 = N1137;
  assign N1161 = N571;
  assign N1173 = N574;
  assign N1185 = N571;
  assign N1197 = N574;
  assign N1209 = N137;
  assign N1213 = N137;
  assign N1216 = N141;
  assign N1223 = N577;
  assign N1235 = N580;
  assign N1247 = N577;
  assign N1259 = N580;
  assign N1271 = N254;
  assign N1280 = N251;
  assign N1292 = N251;
  assign N1303 = N248;
  assign N1315 = N248;
  assign N1327 = N610;
  assign N1339 = N607;
  assign N1351 = N613;
  assign N1363 = N616;
  assign N1375 = N210;
  assign N1378 = N210;
  assign N1381 = N218;
  assign N1384 = N218;
  assign N1387 = N226;
  assign N1390 = N226;
  assign N1393 = N234;
  assign N1396 = N234;
  assign N1415 = N257;
  assign N1418 = N257;
  assign N1421 = N265;
  assign N1424 = N265;
  assign N1427 = N273;
  assign N1430 = N273;
  assign N1433 = N281;
  assign N1436 = N281;
  assign N1455 = N335;
  assign N1462 = N335;
  assign N1469 = N206;
  assign N1479 = N1;
  assign N1482 = N588;
  assign N1492 = N293;
  assign N1495 = N302;
  assign N1498 = N308;
  assign N1501 = N308;
  assign N1504 = N316;
  assign N1507 = N316;
  assign N1510 = N324;
  assign N1513 = N324;
  assign N1516 = N341;
  assign N1519 = N341;
  assign N1522 = N351;
  assign N1525 = N351;
  assign N1542 = N257;
  assign N1545 = N257;
  assign N1548 = N265;
  assign N1551 = N265;
  assign N1554 = N273;
  assign N1557 = N273;
  assign N1560 = N281;
  assign N1563 = N281;
  assign N1566 = N332;
  assign N1573 = N332;
  assign N1580 = N549;
  assign N1594 = N324;
  assign N1597 = N324;
  assign N1600 = N341;
  assign N1603 = N341;
  assign N1606 = N351;
  assign N1609 = N351;
  assign N1612 = N293;
  assign N1615 = N302;
  assign N1618 = N308;
  assign N1621 = N308;
  assign N1624 = N316;
  assign N1627 = N316;
  assign N1630 = N361;
  assign N1633 = N361;
  assign N1636 = N210;
  assign N1639 = N210;
  assign N1642 = N218;
  assign N1645 = N218;
  assign N1648 = N226;
  assign N1651 = N226;
  assign N1654 = N234;
  assign N1657 = N234;
  assign N1663 = N242;
  assign N1675 = N242;
  assign N1685 = N254;
  assign N1697 = N610;
  assign N1709 = N607;
  assign N1721 = N625;
  assign N1727 = N619;
  assign N1731 = N613;
  assign N1743 = N616;
  assign N1761 = N619;
  assign N1769 = N625;
  assign N1777 = N619;
  assign N1785 = N625;
  assign N1793 = N619;
  assign N1800 = N625;
  assign N1807 = N619;
  assign N1814 = N625;
  assign N1821 = N299;
  assign N1824 = N446;
  assign N1827 = N457;
  assign N1830 = N468;
  assign N1833 = N422;
  assign N1836 = N435;
  assign N1839 = N389;
  assign N1842 = N400;
  assign N1845 = N411;
  assign N1848 = N374;
  assign N1851 = N4;
  assign N1854 = N446;
  assign N1857 = N457;
  assign N1860 = N468;
  assign N1863 = N435;
  assign N1866 = N389;
  assign N1869 = N400;
  assign N1872 = N411;
  assign N1875 = N422;
  assign N1878 = N374;
  assign N1881 = N479;
  assign N1884 = N490;
  assign N1887 = N503;
  assign N1890 = N514;
  assign N1893 = N523;
  assign N1896 = N534;
  assign N1899 = N54;
  assign N1902 = N479;
  assign N1905 = N503;
  assign N1908 = N514;
  assign N1911 = N523;
  assign N1914 = N534;
  assign N1917 = N490;
  assign N1920 = N361;
  assign N1923 = N369;
  assign N1926 = N341;
  assign N1929 = N351;
  assign N1932 = N308;
  assign N1935 = N316;
  assign N1938 = N293;
  assign N1941 = N302;
  assign N1944 = N281;
  assign N1947 = N289;
  assign N1950 = N265;
  assign N1953 = N273;
  assign N1956 = N234;
  assign N1959 = N257;
  assign N1962 = N218;
  assign N1965 = N226;
  assign N1968 = N210;
  assign N2139 = N137;
  assign N2142 = N141;
  assign N2309 = N1;
  assign N2387 = N549;
  assign N2527 = N299;
  assign N2584 = N1141;
  assign N2647 = N137;
  assign N2675 = N137;
  assign N2704 = N1;
  assign N2722 = N137;
  assign N2750 = N137;
  assign N2877 = N141;
  assign N2891 = N2623;
  assign N2964 = N588;
  assign N3000 = N206;
  assign N3003 = N206;
  assign N3007 = N206;
  assign N3010 = N206;
  assign N3191 = N299;
  assign N3200 = N206;
  assign N3357 = N1;
  assign N3358 = N1;
  assign N3359 = N1;
  assign N3360 = N1;
  assign N3604 = N299;
  assign N3779 = N324;
  assign N3780 = N324;
  assign N4278 = N4275;
  assign N6466 = N6716;
  assign N6724 = N6877;
  assign N709 = N141;
  assign N7394 = N7474;
  assign N7397 = N7476;
  assign N7431 = N7432;
  assign N816 = N293;
endmodule
