
module s1423(GND, VDD, CK, G0, G1, G10, G11, G12, G13, G14, G15, G16, G2, G3, G4, G5, G6, G7, G701BF, G702, G726, G727, G729, G8, G9);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  input CK;
  wire \DFF_0.CK ;
  wire \DFF_0.D ;
  wire \DFF_0.Q ;
  wire \DFF_1.CK ;
  wire \DFF_1.D ;
  wire \DFF_1.Q ;
  wire \DFF_10.CK ;
  wire \DFF_10.D ;
  wire \DFF_10.Q ;
  wire \DFF_11.CK ;
  wire \DFF_11.D ;
  wire \DFF_11.Q ;
  wire \DFF_12.CK ;
  wire \DFF_12.D ;
  wire \DFF_12.Q ;
  wire \DFF_13.CK ;
  wire \DFF_13.D ;
  wire \DFF_13.Q ;
  wire \DFF_14.CK ;
  wire \DFF_14.D ;
  wire \DFF_14.Q ;
  wire \DFF_15.CK ;
  wire \DFF_15.D ;
  wire \DFF_15.Q ;
  wire \DFF_16.CK ;
  wire \DFF_16.D ;
  wire \DFF_16.Q ;
  wire \DFF_17.CK ;
  wire \DFF_17.D ;
  wire \DFF_17.Q ;
  wire \DFF_18.CK ;
  wire \DFF_18.D ;
  wire \DFF_18.Q ;
  wire \DFF_19.CK ;
  wire \DFF_19.D ;
  wire \DFF_19.Q ;
  wire \DFF_2.CK ;
  wire \DFF_2.D ;
  wire \DFF_2.Q ;
  wire \DFF_20.CK ;
  wire \DFF_20.D ;
  wire \DFF_20.Q ;
  wire \DFF_21.CK ;
  wire \DFF_21.D ;
  wire \DFF_21.Q ;
  wire \DFF_22.CK ;
  wire \DFF_22.D ;
  wire \DFF_22.Q ;
  wire \DFF_23.CK ;
  wire \DFF_23.D ;
  wire \DFF_23.Q ;
  wire \DFF_24.CK ;
  wire \DFF_24.D ;
  wire \DFF_24.Q ;
  wire \DFF_25.CK ;
  wire \DFF_25.D ;
  wire \DFF_25.Q ;
  wire \DFF_26.CK ;
  wire \DFF_26.D ;
  wire \DFF_26.Q ;
  wire \DFF_27.CK ;
  wire \DFF_27.D ;
  wire \DFF_27.Q ;
  wire \DFF_28.CK ;
  wire \DFF_28.D ;
  wire \DFF_28.Q ;
  wire \DFF_29.CK ;
  wire \DFF_29.D ;
  wire \DFF_29.Q ;
  wire \DFF_3.CK ;
  wire \DFF_3.D ;
  wire \DFF_3.Q ;
  wire \DFF_30.CK ;
  wire \DFF_30.D ;
  wire \DFF_30.Q ;
  wire \DFF_31.CK ;
  wire \DFF_31.D ;
  wire \DFF_31.Q ;
  wire \DFF_32.CK ;
  wire \DFF_32.D ;
  wire \DFF_32.Q ;
  wire \DFF_33.CK ;
  wire \DFF_33.D ;
  wire \DFF_33.Q ;
  wire \DFF_34.CK ;
  wire \DFF_34.D ;
  wire \DFF_34.Q ;
  wire \DFF_35.CK ;
  wire \DFF_35.D ;
  wire \DFF_35.Q ;
  wire \DFF_36.CK ;
  wire \DFF_36.D ;
  wire \DFF_36.Q ;
  wire \DFF_37.CK ;
  wire \DFF_37.D ;
  wire \DFF_37.Q ;
  wire \DFF_38.CK ;
  wire \DFF_38.D ;
  wire \DFF_38.Q ;
  wire \DFF_39.CK ;
  wire \DFF_39.D ;
  wire \DFF_39.Q ;
  wire \DFF_4.CK ;
  wire \DFF_4.D ;
  wire \DFF_4.Q ;
  wire \DFF_40.CK ;
  wire \DFF_40.D ;
  wire \DFF_40.Q ;
  wire \DFF_41.CK ;
  wire \DFF_41.D ;
  wire \DFF_41.Q ;
  wire \DFF_42.CK ;
  wire \DFF_42.D ;
  wire \DFF_42.Q ;
  wire \DFF_43.CK ;
  wire \DFF_43.D ;
  wire \DFF_43.Q ;
  wire \DFF_44.CK ;
  wire \DFF_44.D ;
  wire \DFF_44.Q ;
  wire \DFF_45.CK ;
  wire \DFF_45.D ;
  wire \DFF_45.Q ;
  wire \DFF_46.CK ;
  wire \DFF_46.D ;
  wire \DFF_46.Q ;
  wire \DFF_47.CK ;
  wire \DFF_47.D ;
  wire \DFF_47.Q ;
  wire \DFF_48.CK ;
  wire \DFF_48.D ;
  wire \DFF_48.Q ;
  wire \DFF_49.CK ;
  wire \DFF_49.D ;
  wire \DFF_49.Q ;
  wire \DFF_5.CK ;
  wire \DFF_5.D ;
  wire \DFF_5.Q ;
  wire \DFF_50.CK ;
  wire \DFF_50.D ;
  wire \DFF_50.Q ;
  wire \DFF_51.CK ;
  wire \DFF_51.D ;
  wire \DFF_51.Q ;
  wire \DFF_52.CK ;
  wire \DFF_52.D ;
  wire \DFF_52.Q ;
  wire \DFF_53.CK ;
  wire \DFF_53.D ;
  wire \DFF_53.Q ;
  wire \DFF_54.CK ;
  wire \DFF_54.D ;
  wire \DFF_54.Q ;
  wire \DFF_55.CK ;
  wire \DFF_55.D ;
  wire \DFF_55.Q ;
  wire \DFF_56.CK ;
  wire \DFF_56.D ;
  wire \DFF_56.Q ;
  wire \DFF_57.CK ;
  wire \DFF_57.D ;
  wire \DFF_57.Q ;
  wire \DFF_58.CK ;
  wire \DFF_58.D ;
  wire \DFF_58.Q ;
  wire \DFF_59.CK ;
  wire \DFF_59.D ;
  wire \DFF_59.Q ;
  wire \DFF_6.CK ;
  wire \DFF_6.D ;
  wire \DFF_6.Q ;
  wire \DFF_60.CK ;
  wire \DFF_60.D ;
  wire \DFF_60.Q ;
  wire \DFF_61.CK ;
  wire \DFF_61.D ;
  wire \DFF_61.Q ;
  wire \DFF_62.CK ;
  wire \DFF_62.D ;
  wire \DFF_62.Q ;
  wire \DFF_63.CK ;
  wire \DFF_63.D ;
  wire \DFF_63.Q ;
  wire \DFF_64.CK ;
  wire \DFF_64.D ;
  wire \DFF_64.Q ;
  wire \DFF_65.CK ;
  wire \DFF_65.D ;
  wire \DFF_65.Q ;
  wire \DFF_66.CK ;
  wire \DFF_66.D ;
  wire \DFF_66.Q ;
  wire \DFF_67.CK ;
  wire \DFF_67.D ;
  wire \DFF_67.Q ;
  wire \DFF_68.CK ;
  wire \DFF_68.D ;
  wire \DFF_68.Q ;
  wire \DFF_69.CK ;
  wire \DFF_69.D ;
  wire \DFF_69.Q ;
  wire \DFF_7.CK ;
  wire \DFF_7.D ;
  wire \DFF_7.Q ;
  wire \DFF_70.CK ;
  wire \DFF_70.D ;
  wire \DFF_70.Q ;
  wire \DFF_71.CK ;
  wire \DFF_71.D ;
  wire \DFF_71.Q ;
  wire \DFF_72.CK ;
  wire \DFF_72.D ;
  wire \DFF_72.Q ;
  wire \DFF_73.CK ;
  wire \DFF_73.D ;
  wire \DFF_73.Q ;
  wire \DFF_8.CK ;
  wire \DFF_8.D ;
  wire \DFF_8.Q ;
  wire \DFF_9.CK ;
  wire \DFF_9.D ;
  wire \DFF_9.Q ;
  input G0;
  input G1;
  input G10;
  wire G108;
  wire G109;
  input G11;
  wire G112;
  wire G113;
  wire G117;
  wire G118;
  input G12;
  wire G124;
  wire G125;
  wire G128;
  wire G129;
  input G13;
  wire G139;
  input G14;
  wire G140;
  wire G143;
  wire G144;
  wire G148;
  wire G149;
  input G15;
  wire G153;
  wire G154;
  wire G158;
  wire G159;
  input G16;
  wire G165;
  wire G166;
  wire G174;
  wire G175;
  wire G179;
  wire G188;
  wire G189;
  wire G192;
  wire G193;
  wire G197;
  wire G198;
  input G2;
  wire G207;
  wire G208;
  wire G213;
  wire G214;
  wire G217;
  wire G218;
  wire G22;
  wire G23;
  wire G237;
  wire G24;
  wire G242;
  wire G247;
  wire G25;
  wire G252;
  wire G26;
  wire G260;
  wire G27;
  wire G28;
  wire G29;
  input G3;
  wire G30;
  wire G302;
  wire G303;
  wire G308;
  wire G309;
  wire G31;
  wire G314;
  wire G315;
  wire G32;
  wire G320;
  wire G321;
  wire G328;
  wire G328BF;
  wire G33;
  wire G332;
  wire G332BF;
  wire G34;
  wire G343;
  wire G347;
  wire G35;
  wire G351;
  wire G36;
  wire G360;
  wire G365;
  wire G37;
  wire G373;
  wire G379;
  wire G38;
  wire G384;
  wire G39;
  wire G392;
  wire G397;
  input G4;
  wire G40;
  wire G405;
  wire G407;
  wire G408;
  wire G41;
  wire G416;
  wire G42;
  wire G424;
  wire G426;
  wire G427;
  wire G43;
  wire G437;
  wire G438;
  wire G44;
  wire G440;
  wire G441;
  wire G446;
  wire G447;
  wire G45;
  wire G450;
  wire G451;
  wire G459;
  wire G46;
  wire G464;
  wire G469;
  wire G47;
  wire G477;
  wire G48;
  wire G486;
  wire G49;
  wire G494;
  wire G498;
  input G5;
  wire G50;
  wire G503;
  wire G504;
  wire G507;
  wire G51;
  wire G510;
  wire G52;
  wire G526;
  wire G53;
  wire G531;
  wire G536;
  wire G54;
  wire G541;
  wire G548;
  wire G55;
  wire G56;
  wire G565;
  wire G569;
  wire G57;
  wire G573;
  wire G577;
  wire G58;
  wire G59;
  wire G590;
  input G6;
  wire G60;
  wire G608;
  wire G61;
  wire G613;
  wire G617;
  wire G62;
  wire G620;
  wire G623;
  wire G626;
  wire G629;
  wire G63;
  wire G632;
  wire G635;
  wire G638;
  wire G64;
  wire G641;
  wire G644;
  wire G65;
  wire G656;
  wire G657;
  wire G659;
  wire G66;
  wire G662;
  wire G663;
  wire G668;
  wire G669;
  wire G67;
  wire G674;
  wire G675;
  wire G678;
  wire G68;
  wire G682;
  wire G687;
  wire G69;
  wire G693;
  wire G696;
  input G7;
  wire G70;
  wire G701;
  output G701BF;
  output G702;
  wire G704;
  wire G705;
  wire G706;
  wire G707;
  wire G71;
  wire G711;
  wire G713;
  wire G714;
  wire G715;
  wire G716;
  wire G717;
  wire G718;
  wire G719;
  wire G72;
  wire G720;
  wire G721;
  wire G722;
  wire G723;
  wire G724;
  wire G725;
  output G726;
  output G727;
  wire G728;
  output G729;
  wire G73;
  wire G74;
  wire G75;
  wire G76;
  wire G77;
  wire G78;
  wire G79;
  input G8;
  wire G80;
  wire G81;
  wire G82;
  wire G83;
  wire G84;
  wire G85;
  wire G86;
  wire G87;
  wire G88;
  wire G89;
  input G9;
  wire G90;
  wire G91;
  wire G92;
  wire G93;
  wire G94;
  wire G95;
  input GND;
  wire II1211;
  input VDD;
  al_and2 _233_ (
    .a(\DFF_28.Q ),
    .b(\DFF_25.Q ),
    .y(_000_)
  );
  al_and3 _234_ (
    .a(\DFF_27.Q ),
    .b(\DFF_26.Q ),
    .c(_000_),
    .y(_001_)
  );
  al_or3 _235_ (
    .a(\DFF_27.Q ),
    .b(\DFF_26.Q ),
    .c(\DFF_25.Q ),
    .y(_002_)
  );
  al_or3 _236_ (
    .a(G15),
    .b(\DFF_28.Q ),
    .c(_002_),
    .y(_003_)
  );
  al_nand2 _237_ (
    .a(\DFF_0.Q ),
    .b(_003_),
    .y(_004_)
  );
  al_ao21ftf _238_ (
    .a(G15),
    .b(_001_),
    .c(_004_),
    .y(\DFF_0.D )
  );
  al_mux2l _239_ (
    .a(\DFF_0.Q ),
    .b(\DFF_1.Q ),
    .s(G15),
    .y(\DFF_1.D )
  );
  al_inv _240_ (
    .a(G15),
    .y(G701BF)
  );
  al_inv _241_ (
    .a(G14),
    .y(_005_)
  );
  al_inv _242_ (
    .a(\DFF_61.Q ),
    .y(_006_)
  );
  al_nor2 _243_ (
    .a(\DFF_52.Q ),
    .b(\DFF_57.Q ),
    .y(_007_)
  );
  al_nand2 _244_ (
    .a(\DFF_52.Q ),
    .b(\DFF_57.Q ),
    .y(_008_)
  );
  al_nand2ft _245_ (
    .a(_007_),
    .b(_008_),
    .y(_009_)
  );
  al_nand2ft _246_ (
    .a(\DFF_53.Q ),
    .b(\DFF_58.Q ),
    .y(_010_)
  );
  al_nand2ft _247_ (
    .a(\DFF_58.Q ),
    .b(\DFF_53.Q ),
    .y(_011_)
  );
  al_and3 _248_ (
    .a(_010_),
    .b(_011_),
    .c(_009_),
    .y(_012_)
  );
  al_and2ft _249_ (
    .a(\DFF_59.Q ),
    .b(\DFF_54.Q ),
    .y(_013_)
  );
  al_and2ft _250_ (
    .a(\DFF_54.Q ),
    .b(\DFF_59.Q ),
    .y(_014_)
  );
  al_nor2 _251_ (
    .a(\DFF_55.Q ),
    .b(\DFF_60.Q ),
    .y(_015_)
  );
  al_nand2 _252_ (
    .a(\DFF_55.Q ),
    .b(\DFF_60.Q ),
    .y(_016_)
  );
  al_nand2ft _253_ (
    .a(_015_),
    .b(_016_),
    .y(_017_)
  );
  al_nand3fft _254_ (
    .a(_013_),
    .b(_014_),
    .c(_017_),
    .y(_018_)
  );
  al_inv _255_ (
    .a(\DFF_56.Q ),
    .y(_019_)
  );
  al_or3 _256_ (
    .a(\DFF_57.Q ),
    .b(\DFF_58.Q ),
    .c(\DFF_59.Q ),
    .y(_020_)
  );
  al_oa21ttf _257_ (
    .a(\DFF_60.Q ),
    .b(_020_),
    .c(_019_),
    .y(_021_)
  );
  al_or3 _258_ (
    .a(\DFF_56.Q ),
    .b(\DFF_60.Q ),
    .c(_020_),
    .y(_022_)
  );
  al_nor2ft _259_ (
    .a(_022_),
    .b(_021_),
    .y(_023_)
  );
  al_and3ftt _260_ (
    .a(_018_),
    .b(_012_),
    .c(_023_),
    .y(_024_)
  );
  al_and2ft _261_ (
    .a(\DFF_44.Q ),
    .b(G16),
    .y(_025_)
  );
  al_nand3 _262_ (
    .a(_006_),
    .b(_025_),
    .c(_024_),
    .y(_026_)
  );
  al_and2 _263_ (
    .a(\DFF_68.Q ),
    .b(_026_),
    .y(_027_)
  );
  al_inv _264_ (
    .a(\DFF_12.Q ),
    .y(_028_)
  );
  al_mux2h _265_ (
    .a(\DFF_13.Q ),
    .b(_028_),
    .s(\DFF_70.Q ),
    .y(_029_)
  );
  al_mux2l _266_ (
    .a(\DFF_16.Q ),
    .b(_029_),
    .s(_027_),
    .y(_030_)
  );
  al_oa21ttf _267_ (
    .a(\DFF_41.Q ),
    .b(_030_),
    .c(_005_),
    .y(\DFF_41.D )
  );
  al_inv _268_ (
    .a(\DFF_45.Q ),
    .y(_031_)
  );
  al_or3 _269_ (
    .a(\DFF_48.Q ),
    .b(\DFF_46.Q ),
    .c(\DFF_47.Q ),
    .y(_032_)
  );
  al_ao21ftf _270_ (
    .a(\DFF_49.Q ),
    .b(_032_),
    .c(_031_),
    .y(_033_)
  );
  al_oai21ftt _271_ (
    .a(\DFF_50.Q ),
    .b(\DFF_48.Q ),
    .c(\DFF_46.Q ),
    .y(_034_)
  );
  al_ao21ftf _272_ (
    .a(\DFF_46.Q ),
    .b(\DFF_50.Q ),
    .c(_034_),
    .y(_035_)
  );
  al_oa21ftt _273_ (
    .a(\DFF_49.Q ),
    .b(\DFF_48.Q ),
    .c(\DFF_45.Q ),
    .y(_036_)
  );
  al_nand3ftt _274_ (
    .a(\DFF_48.Q ),
    .b(\DFF_47.Q ),
    .c(\DFF_51.Q ),
    .y(_037_)
  );
  al_or2 _275_ (
    .a(\DFF_47.Q ),
    .b(\DFF_51.Q ),
    .y(_038_)
  );
  al_aoi21 _276_ (
    .a(_037_),
    .b(_038_),
    .c(_036_),
    .y(_039_)
  );
  al_nand3ftt _277_ (
    .a(_035_),
    .b(_033_),
    .c(_039_),
    .y(_040_)
  );
  al_mux2l _278_ (
    .a(\DFF_42.Q ),
    .b(\DFF_41.Q ),
    .s(_040_),
    .y(_041_)
  );
  al_and2 _279_ (
    .a(G14),
    .b(_041_),
    .y(\DFF_42.D )
  );
  al_aoi21ftf _280_ (
    .a(\DFF_43.Q ),
    .b(_040_),
    .c(G14),
    .y(\DFF_43.D )
  );
  al_mux2l _281_ (
    .a(\DFF_44.Q ),
    .b(\DFF_43.Q ),
    .s(_040_),
    .y(_042_)
  );
  al_and2 _282_ (
    .a(G14),
    .b(_042_),
    .y(\DFF_44.D )
  );
  al_inv _283_ (
    .a(\DFF_31.Q ),
    .y(_043_)
  );
  al_inv _284_ (
    .a(\DFF_37.Q ),
    .y(_044_)
  );
  al_inv _285_ (
    .a(\DFF_36.Q ),
    .y(_045_)
  );
  al_inv _286_ (
    .a(\DFF_11.Q ),
    .y(_046_)
  );
  al_inv _287_ (
    .a(\DFF_7.Q ),
    .y(_047_)
  );
  al_inv _288_ (
    .a(\DFF_70.Q ),
    .y(_048_)
  );
  al_inv _289_ (
    .a(\DFF_5.Q ),
    .y(_049_)
  );
  al_inv _290_ (
    .a(\DFF_2.Q ),
    .y(_050_)
  );
  al_or2 _291_ (
    .a(\DFF_68.Q ),
    .b(G4),
    .y(_051_)
  );
  al_inv _292_ (
    .a(\DFF_68.Q ),
    .y(_052_)
  );
  al_nand2ft _293_ (
    .a(\DFF_68.Q ),
    .b(G8),
    .y(_053_)
  );
  al_ao21ftf _294_ (
    .a(\DFF_42.Q ),
    .b(\DFF_68.Q ),
    .c(_053_),
    .y(_054_)
  );
  al_mux2l _295_ (
    .a(\DFF_62.Q ),
    .b(\DFF_63.Q ),
    .s(_054_),
    .y(_055_)
  );
  al_nand3fft _296_ (
    .a(_052_),
    .b(_019_),
    .c(_055_),
    .y(_056_)
  );
  al_and3 _297_ (
    .a(\DFF_24.Q ),
    .b(_051_),
    .c(_056_),
    .y(_057_)
  );
  al_or2 _298_ (
    .a(\DFF_68.Q ),
    .b(G3),
    .y(_058_)
  );
  al_nand2 _299_ (
    .a(\DFF_42.Q ),
    .b(\DFF_68.Q ),
    .y(_059_)
  );
  al_or2 _300_ (
    .a(\DFF_68.Q ),
    .b(G8),
    .y(_060_)
  );
  al_nand3ftt _301_ (
    .a(\DFF_62.Q ),
    .b(_060_),
    .c(_059_),
    .y(_061_)
  );
  al_nand2ft _302_ (
    .a(\DFF_42.Q ),
    .b(\DFF_68.Q ),
    .y(_062_)
  );
  al_nand3ftt _303_ (
    .a(\DFF_63.Q ),
    .b(_053_),
    .c(_062_),
    .y(_063_)
  );
  al_and2 _304_ (
    .a(\DFF_68.Q ),
    .b(\DFF_55.Q ),
    .y(_064_)
  );
  al_nand3 _305_ (
    .a(_064_),
    .b(_063_),
    .c(_061_),
    .y(_065_)
  );
  al_and3 _306_ (
    .a(\DFF_23.Q ),
    .b(_058_),
    .c(_065_),
    .y(_066_)
  );
  al_or2 _307_ (
    .a(\DFF_68.Q ),
    .b(G2),
    .y(_067_)
  );
  al_and2 _308_ (
    .a(\DFF_68.Q ),
    .b(\DFF_54.Q ),
    .y(_068_)
  );
  al_nand3 _309_ (
    .a(_068_),
    .b(_063_),
    .c(_061_),
    .y(_069_)
  );
  al_and2 _310_ (
    .a(_067_),
    .b(_069_),
    .y(_070_)
  );
  al_ao21 _311_ (
    .a(\DFF_22.Q ),
    .b(_070_),
    .c(_066_),
    .y(_071_)
  );
  al_and2 _312_ (
    .a(\DFF_68.Q ),
    .b(\DFF_52.Q ),
    .y(_072_)
  );
  al_nand3 _313_ (
    .a(_072_),
    .b(_063_),
    .c(_061_),
    .y(_073_)
  );
  al_or2 _314_ (
    .a(\DFF_68.Q ),
    .b(G0),
    .y(_074_)
  );
  al_and3 _315_ (
    .a(\DFF_20.Q ),
    .b(_074_),
    .c(_073_),
    .y(_075_)
  );
  al_and2 _316_ (
    .a(\DFF_68.Q ),
    .b(\DFF_53.Q ),
    .y(_076_)
  );
  al_nand3 _317_ (
    .a(_076_),
    .b(_063_),
    .c(_061_),
    .y(_077_)
  );
  al_or2 _318_ (
    .a(\DFF_68.Q ),
    .b(G1),
    .y(_078_)
  );
  al_ao21 _319_ (
    .a(_078_),
    .b(_077_),
    .c(\DFF_21.Q ),
    .y(_079_)
  );
  al_nand3 _320_ (
    .a(\DFF_21.Q ),
    .b(_078_),
    .c(_077_),
    .y(_080_)
  );
  al_nand3ftt _321_ (
    .a(_075_),
    .b(_079_),
    .c(_080_),
    .y(_081_)
  );
  al_nand2 _322_ (
    .a(_078_),
    .b(_077_),
    .y(_082_)
  );
  al_ao21 _323_ (
    .a(_067_),
    .b(_069_),
    .c(\DFF_22.Q ),
    .y(_083_)
  );
  al_aoi21ftf _324_ (
    .a(\DFF_21.Q ),
    .b(_082_),
    .c(_083_),
    .y(_084_)
  );
  al_ao21 _325_ (
    .a(_084_),
    .b(_081_),
    .c(_071_),
    .y(_085_)
  );
  al_inv _326_ (
    .a(\DFF_24.Q ),
    .y(_086_)
  );
  al_nand2 _327_ (
    .a(_051_),
    .b(_056_),
    .y(_087_)
  );
  al_aoi21 _328_ (
    .a(_058_),
    .b(_065_),
    .c(\DFF_23.Q ),
    .y(_088_)
  );
  al_aoi21 _329_ (
    .a(_086_),
    .b(_087_),
    .c(_088_),
    .y(_089_)
  );
  al_aoi21 _330_ (
    .a(_089_),
    .b(_085_),
    .c(_057_),
    .y(_090_)
  );
  al_and3 _331_ (
    .a(_050_),
    .b(\DFF_3.Q ),
    .c(_090_),
    .y(_091_)
  );
  al_and3 _332_ (
    .a(_049_),
    .b(\DFF_4.Q ),
    .c(_091_),
    .y(_092_)
  );
  al_ao21 _333_ (
    .a(\DFF_6.Q ),
    .b(_092_),
    .c(_048_),
    .y(_093_)
  );
  al_and3 _334_ (
    .a(_047_),
    .b(\DFF_8.Q ),
    .c(_093_),
    .y(_094_)
  );
  al_and3 _335_ (
    .a(\DFF_9.Q ),
    .b(\DFF_10.Q ),
    .c(_094_),
    .y(_095_)
  );
  al_nand3fft _336_ (
    .a(\DFF_12.Q ),
    .b(_046_),
    .c(_095_),
    .y(_096_)
  );
  al_nand2 _337_ (
    .a(\DFF_70.Q ),
    .b(_096_),
    .y(_097_)
  );
  al_inv _338_ (
    .a(\DFF_19.Q ),
    .y(_098_)
  );
  al_aoi21 _339_ (
    .a(\DFF_70.Q ),
    .b(_096_),
    .c(\DFF_17.Q ),
    .y(_099_)
  );
  al_nand3fft _340_ (
    .a(\DFF_18.Q ),
    .b(_098_),
    .c(_099_),
    .y(_100_)
  );
  al_aoi21 _341_ (
    .a(\DFF_69.Q ),
    .b(_100_),
    .c(\DFF_14.Q ),
    .y(_101_)
  );
  al_and3 _342_ (
    .a(\DFF_16.Q ),
    .b(\DFF_15.Q ),
    .c(_101_),
    .y(_102_)
  );
  al_mux2h _343_ (
    .a(_097_),
    .b(_102_),
    .s(_027_),
    .y(_103_)
  );
  al_nand3fft _344_ (
    .a(_044_),
    .b(_045_),
    .c(_103_),
    .y(_104_)
  );
  al_aoi21 _345_ (
    .a(\DFF_69.Q ),
    .b(_104_),
    .c(_043_),
    .y(_105_)
  );
  al_and2 _346_ (
    .a(\DFF_69.Q ),
    .b(\DFF_40.Q ),
    .y(_106_)
  );
  al_nand3 _347_ (
    .a(\DFF_39.Q ),
    .b(_106_),
    .c(_105_),
    .y(_107_)
  );
  al_inv _348_ (
    .a(\DFF_69.Q ),
    .y(_108_)
  );
  al_oa21ftf _349_ (
    .a(_108_),
    .b(_104_),
    .c(_052_),
    .y(_109_)
  );
  al_nand3 _350_ (
    .a(_031_),
    .b(_109_),
    .c(_107_),
    .y(_110_)
  );
  al_aoi21 _351_ (
    .a(_109_),
    .b(_107_),
    .c(_031_),
    .y(_111_)
  );
  al_and2 _352_ (
    .a(G14),
    .b(_040_),
    .y(_112_)
  );
  al_inv _353_ (
    .a(_112_),
    .y(_113_)
  );
  al_and3fft _354_ (
    .a(_113_),
    .b(_111_),
    .c(_110_),
    .y(\DFF_45.D )
  );
  al_nand2 _355_ (
    .a(_109_),
    .b(_107_),
    .y(_114_)
  );
  al_and3 _356_ (
    .a(\DFF_45.Q ),
    .b(\DFF_46.Q ),
    .c(_114_),
    .y(_115_)
  );
  al_aoi21 _357_ (
    .a(\DFF_45.Q ),
    .b(_114_),
    .c(\DFF_46.Q ),
    .y(_116_)
  );
  al_nor3ftt _358_ (
    .a(_112_),
    .b(_115_),
    .c(_116_),
    .y(\DFF_46.D )
  );
  al_inv _359_ (
    .a(\DFF_46.Q ),
    .y(_117_)
  );
  al_inv _360_ (
    .a(\DFF_47.Q ),
    .y(_118_)
  );
  al_nand3fft _361_ (
    .a(_117_),
    .b(_118_),
    .c(_111_),
    .y(_119_)
  );
  al_ao21 _362_ (
    .a(\DFF_46.Q ),
    .b(_111_),
    .c(\DFF_47.Q ),
    .y(_120_)
  );
  al_and3 _363_ (
    .a(_112_),
    .b(_119_),
    .c(_120_),
    .y(\DFF_47.D )
  );
  al_nand2 _364_ (
    .a(\DFF_48.Q ),
    .b(_119_),
    .y(_121_)
  );
  al_nand3fft _365_ (
    .a(\DFF_48.Q ),
    .b(_118_),
    .c(_115_),
    .y(_122_)
  );
  al_aoi21 _366_ (
    .a(_122_),
    .b(_121_),
    .c(_113_),
    .y(\DFF_48.D )
  );
  al_oa21ftf _367_ (
    .a(\DFF_68.Q ),
    .b(_040_),
    .c(_005_),
    .y(_123_)
  );
  al_mux2l _368_ (
    .a(G3),
    .b(G0),
    .s(\DFF_41.Q ),
    .y(_124_)
  );
  al_mux2l _369_ (
    .a(\DFF_49.Q ),
    .b(_124_),
    .s(_123_),
    .y(\DFF_49.D )
  );
  al_mux2l _370_ (
    .a(G4),
    .b(G1),
    .s(\DFF_41.Q ),
    .y(_125_)
  );
  al_mux2l _371_ (
    .a(\DFF_50.Q ),
    .b(_125_),
    .s(_123_),
    .y(\DFF_50.D )
  );
  al_mux2l _372_ (
    .a(G5),
    .b(G2),
    .s(\DFF_41.Q ),
    .y(_126_)
  );
  al_mux2l _373_ (
    .a(\DFF_51.Q ),
    .b(_126_),
    .s(_123_),
    .y(\DFF_51.D )
  );
  al_and2 _374_ (
    .a(\DFF_15.Q ),
    .b(_101_),
    .y(_127_)
  );
  al_nand3ftt _375_ (
    .a(\DFF_16.Q ),
    .b(_027_),
    .c(_127_),
    .y(_128_)
  );
  al_nand3fft _376_ (
    .a(_028_),
    .b(_046_),
    .c(_095_),
    .y(_129_)
  );
  al_ao21 _377_ (
    .a(\DFF_70.Q ),
    .b(_129_),
    .c(_027_),
    .y(_130_)
  );
  al_aoi21 _378_ (
    .a(_130_),
    .b(_128_),
    .c(_024_),
    .y(_131_)
  );
  al_nand3fft _379_ (
    .a(_052_),
    .b(_005_),
    .c(_040_),
    .y(_132_)
  );
  al_ao21ftf _380_ (
    .a(G9),
    .b(_052_),
    .c(_132_),
    .y(_133_)
  );
  al_aoi21ttf _381_ (
    .a(\DFF_52.Q ),
    .b(_131_),
    .c(_133_),
    .y(_134_)
  );
  al_oa21 _382_ (
    .a(\DFF_52.Q ),
    .b(_131_),
    .c(_134_),
    .y(\DFF_52.D )
  );
  al_and3 _383_ (
    .a(\DFF_52.Q ),
    .b(\DFF_53.Q ),
    .c(_131_),
    .y(_135_)
  );
  al_aoi21 _384_ (
    .a(\DFF_52.Q ),
    .b(_131_),
    .c(\DFF_53.Q ),
    .y(_136_)
  );
  al_nor3ftt _385_ (
    .a(_133_),
    .b(_135_),
    .c(_136_),
    .y(\DFF_53.D )
  );
  al_and2 _386_ (
    .a(\DFF_54.Q ),
    .b(_135_),
    .y(_137_)
  );
  al_or2 _387_ (
    .a(\DFF_54.Q ),
    .b(_135_),
    .y(_138_)
  );
  al_nor3fft _388_ (
    .a(_133_),
    .b(_138_),
    .c(_137_),
    .y(\DFF_54.D )
  );
  al_nand3 _389_ (
    .a(\DFF_54.Q ),
    .b(\DFF_55.Q ),
    .c(_135_),
    .y(_139_)
  );
  al_ao21 _390_ (
    .a(\DFF_54.Q ),
    .b(_135_),
    .c(\DFF_55.Q ),
    .y(_140_)
  );
  al_and3 _391_ (
    .a(_133_),
    .b(_139_),
    .c(_140_),
    .y(\DFF_55.D )
  );
  al_nand2 _392_ (
    .a(\DFF_56.Q ),
    .b(_139_),
    .y(_141_)
  );
  al_nand3 _393_ (
    .a(_019_),
    .b(\DFF_55.Q ),
    .c(_137_),
    .y(_142_)
  );
  al_aoi21ttf _394_ (
    .a(_141_),
    .b(_142_),
    .c(_133_),
    .y(\DFF_56.D )
  );
  al_oa21ftf _395_ (
    .a(\DFF_69.Q ),
    .b(_040_),
    .c(_005_),
    .y(_143_)
  );
  al_mux2l _396_ (
    .a(\DFF_57.Q ),
    .b(G6),
    .s(_143_),
    .y(\DFF_57.D )
  );
  al_mux2l _397_ (
    .a(\DFF_58.Q ),
    .b(G7),
    .s(_143_),
    .y(\DFF_58.D )
  );
  al_mux2l _398_ (
    .a(\DFF_59.Q ),
    .b(G8),
    .s(_143_),
    .y(\DFF_59.D )
  );
  al_mux2l _399_ (
    .a(\DFF_60.Q ),
    .b(G9),
    .s(_143_),
    .y(\DFF_60.D )
  );
  al_oai21ftt _400_ (
    .a(_024_),
    .b(_030_),
    .c(_133_),
    .y(_144_)
  );
  al_oa21ftf _401_ (
    .a(_006_),
    .b(_131_),
    .c(_144_),
    .y(\DFF_61.D )
  );
  al_mux2l _402_ (
    .a(\DFF_62.Q ),
    .b(G10),
    .s(_143_),
    .y(\DFF_62.D )
  );
  al_mux2l _403_ (
    .a(\DFF_63.Q ),
    .b(G11),
    .s(_143_),
    .y(\DFF_63.D )
  );
  al_and2 _404_ (
    .a(G13),
    .b(G14),
    .y(\DFF_64.D )
  );
  al_oa21 _405_ (
    .a(G11),
    .b(\DFF_65.Q ),
    .c(G14),
    .y(_145_)
  );
  al_aoi21ttf _406_ (
    .a(\DFF_72.Q ),
    .b(G11),
    .c(_145_),
    .y(\DFF_65.D )
  );
  al_mux2l _407_ (
    .a(\DFF_65.Q ),
    .b(\DFF_66.Q ),
    .s(G11),
    .y(_146_)
  );
  al_and2 _408_ (
    .a(G14),
    .b(_146_),
    .y(\DFF_66.D )
  );
  al_mux2l _409_ (
    .a(\DFF_66.Q ),
    .b(\DFF_67.Q ),
    .s(G11),
    .y(_147_)
  );
  al_and2 _410_ (
    .a(G14),
    .b(_147_),
    .y(\DFF_67.D )
  );
  al_nand3 _411_ (
    .a(\DFF_40.Q ),
    .b(\DFF_39.Q ),
    .c(_105_),
    .y(_148_)
  );
  al_and3ftt _412_ (
    .a(\DFF_72.Q ),
    .b(\DFF_6.Q ),
    .c(_092_),
    .y(_149_)
  );
  al_oa21ftf _413_ (
    .a(\DFF_65.Q ),
    .b(_096_),
    .c(_149_),
    .y(_150_)
  );
  al_oa21ftf _414_ (
    .a(\DFF_66.Q ),
    .b(_100_),
    .c(\DFF_68.Q ),
    .y(_151_)
  );
  al_nand2 _415_ (
    .a(_150_),
    .b(_151_),
    .y(_152_)
  );
  al_oa21ftf _416_ (
    .a(\DFF_67.Q ),
    .b(_148_),
    .c(_152_),
    .y(G702)
  );
  al_aoi21ftt _417_ (
    .a(G6),
    .b(_052_),
    .c(_027_),
    .y(_153_)
  );
  al_nand3fft _418_ (
    .a(_052_),
    .b(\DFF_61.Q ),
    .c(_024_),
    .y(_154_)
  );
  al_aoi21ftf _419_ (
    .a(G5),
    .b(_052_),
    .c(_154_),
    .y(_155_)
  );
  al_aoi21 _420_ (
    .a(_074_),
    .b(_073_),
    .c(\DFF_20.Q ),
    .y(_156_)
  );
  al_and3fft _421_ (
    .a(_156_),
    .b(_057_),
    .c(_083_),
    .y(_157_)
  );
  al_nand3fft _422_ (
    .a(_071_),
    .b(_081_),
    .c(_089_),
    .y(_158_)
  );
  al_oai21ftf _423_ (
    .a(_157_),
    .b(_158_),
    .c(_155_),
    .y(_159_)
  );
  al_ao21ttf _424_ (
    .a(_030_),
    .b(_159_),
    .c(_090_),
    .y(_160_)
  );
  al_oai21ftt _425_ (
    .a(\DFF_37.Q ),
    .b(\DFF_69.Q ),
    .c(\DFF_68.Q ),
    .y(_161_)
  );
  al_nor2 _426_ (
    .a(\DFF_13.Q ),
    .b(\DFF_68.Q ),
    .y(_162_)
  );
  al_oai21ttf _427_ (
    .a(_161_),
    .b(_106_),
    .c(_162_),
    .y(_163_)
  );
  al_aoi21 _428_ (
    .a(_163_),
    .b(_153_),
    .c(_005_),
    .y(_164_)
  );
  al_aoi21ftf _429_ (
    .a(_153_),
    .b(_160_),
    .c(_164_),
    .y(\DFF_71.D )
  );
  al_oa21 _430_ (
    .a(\DFF_72.Q ),
    .b(G11),
    .c(G14),
    .y(_165_)
  );
  al_aoi21ttf _431_ (
    .a(G11),
    .b(\DFF_67.Q ),
    .c(_165_),
    .y(\DFF_72.D )
  );
  al_and3 _432_ (
    .a(G14),
    .b(\DFF_61.Q ),
    .c(_055_),
    .y(_166_)
  );
  al_and2 _433_ (
    .a(_166_),
    .b(_030_),
    .y(\DFF_73.D )
  );
  al_aoi21 _434_ (
    .a(G14),
    .b(_040_),
    .c(\DFF_68.Q ),
    .y(G727)
  );
  al_oai21 _435_ (
    .a(\DFF_68.Q ),
    .b(G10),
    .c(\DFF_64.Q ),
    .y(_167_)
  );
  al_nand3 _436_ (
    .a(G13),
    .b(G14),
    .c(_167_),
    .y(\DFF_68.D )
  );
  al_or2 _437_ (
    .a(\DFF_69.Q ),
    .b(G10),
    .y(_168_)
  );
  al_nand2ft _438_ (
    .a(\DFF_64.Q ),
    .b(G13),
    .y(_169_)
  );
  al_aoi21ftf _439_ (
    .a(\DFF_68.Q ),
    .b(G10),
    .c(_169_),
    .y(_170_)
  );
  al_ao21ttf _440_ (
    .a(_168_),
    .b(_170_),
    .c(\DFF_64.D ),
    .y(\DFF_69.D )
  );
  al_mux2l _441_ (
    .a(\DFF_69.Q ),
    .b(\DFF_70.Q ),
    .s(G10),
    .y(_171_)
  );
  al_ao21ttf _442_ (
    .a(_169_),
    .b(_171_),
    .c(\DFF_64.D ),
    .y(\DFF_70.D )
  );
  al_nand2 _443_ (
    .a(_050_),
    .b(_090_),
    .y(_172_)
  );
  al_or2 _444_ (
    .a(_050_),
    .b(_090_),
    .y(_173_)
  );
  al_aoi21 _445_ (
    .a(_172_),
    .b(_173_),
    .c(_005_),
    .y(\DFF_2.D )
  );
  al_aoi21 _446_ (
    .a(_050_),
    .b(_090_),
    .c(\DFF_3.Q ),
    .y(_174_)
  );
  al_nor3ftt _447_ (
    .a(G14),
    .b(_091_),
    .c(_174_),
    .y(\DFF_3.D )
  );
  al_and2 _448_ (
    .a(\DFF_4.Q ),
    .b(_091_),
    .y(_175_)
  );
  al_or2 _449_ (
    .a(\DFF_4.Q ),
    .b(_091_),
    .y(_176_)
  );
  al_nor3fft _450_ (
    .a(G14),
    .b(_176_),
    .c(_175_),
    .y(\DFF_4.D )
  );
  al_ao21 _451_ (
    .a(\DFF_4.Q ),
    .b(_091_),
    .c(_049_),
    .y(_177_)
  );
  al_aoi21ftt _452_ (
    .a(_092_),
    .b(_177_),
    .c(_005_),
    .y(\DFF_5.D )
  );
  al_nand3 _453_ (
    .a(_049_),
    .b(\DFF_6.Q ),
    .c(_175_),
    .y(_178_)
  );
  al_or2 _454_ (
    .a(\DFF_6.Q ),
    .b(_092_),
    .y(_179_)
  );
  al_and3 _455_ (
    .a(G14),
    .b(_178_),
    .c(_179_),
    .y(\DFF_6.D )
  );
  al_aoi21 _456_ (
    .a(\DFF_70.Q ),
    .b(_178_),
    .c(\DFF_7.Q ),
    .y(_180_)
  );
  al_nand3fft _457_ (
    .a(_047_),
    .b(_048_),
    .c(_178_),
    .y(_181_)
  );
  al_oa21ftf _458_ (
    .a(_181_),
    .b(_180_),
    .c(_005_),
    .y(\DFF_7.D )
  );
  al_aoi21 _459_ (
    .a(_047_),
    .b(_093_),
    .c(\DFF_8.Q ),
    .y(_182_)
  );
  al_nor3ftt _460_ (
    .a(G14),
    .b(_094_),
    .c(_182_),
    .y(\DFF_8.D )
  );
  al_and3 _461_ (
    .a(\DFF_8.Q ),
    .b(\DFF_9.Q ),
    .c(_180_),
    .y(_183_)
  );
  al_or2 _462_ (
    .a(\DFF_9.Q ),
    .b(_094_),
    .y(_184_)
  );
  al_nor3fft _463_ (
    .a(G14),
    .b(_184_),
    .c(_183_),
    .y(\DFF_9.D )
  );
  al_aoi21 _464_ (
    .a(\DFF_9.Q ),
    .b(_094_),
    .c(\DFF_10.Q ),
    .y(_185_)
  );
  al_nor3ftt _465_ (
    .a(G14),
    .b(_095_),
    .c(_185_),
    .y(\DFF_10.D )
  );
  al_aoi21 _466_ (
    .a(\DFF_11.Q ),
    .b(_095_),
    .c(_005_),
    .y(_186_)
  );
  al_aoi21ftf _467_ (
    .a(_095_),
    .b(_046_),
    .c(_186_),
    .y(\DFF_11.D )
  );
  al_ao21 _468_ (
    .a(\DFF_11.Q ),
    .b(_095_),
    .c(\DFF_12.Q ),
    .y(_187_)
  );
  al_and3 _469_ (
    .a(G14),
    .b(_129_),
    .c(_187_),
    .y(\DFF_12.D )
  );
  al_and2ft _470_ (
    .a(\DFF_13.Q ),
    .b(G14),
    .y(\DFF_13.D )
  );
  al_nand3 _471_ (
    .a(\DFF_14.Q ),
    .b(\DFF_69.Q ),
    .c(_100_),
    .y(_188_)
  );
  al_oa21ftf _472_ (
    .a(_188_),
    .b(_101_),
    .c(_005_),
    .y(\DFF_14.D )
  );
  al_or2 _473_ (
    .a(\DFF_15.Q ),
    .b(_101_),
    .y(_189_)
  );
  al_nor3fft _474_ (
    .a(G14),
    .b(_189_),
    .c(_127_),
    .y(\DFF_15.D )
  );
  al_aoi21 _475_ (
    .a(\DFF_15.Q ),
    .b(_101_),
    .c(\DFF_16.Q ),
    .y(_190_)
  );
  al_nor3ftt _476_ (
    .a(G14),
    .b(_102_),
    .c(_190_),
    .y(\DFF_16.D )
  );
  al_inv _477_ (
    .a(\DFF_17.Q ),
    .y(_191_)
  );
  al_nand3fft _478_ (
    .a(_048_),
    .b(_191_),
    .c(_096_),
    .y(_192_)
  );
  al_oa21ftf _479_ (
    .a(_192_),
    .b(_099_),
    .c(_005_),
    .y(\DFF_17.D )
  );
  al_nand3fft _480_ (
    .a(\DFF_17.Q ),
    .b(\DFF_18.Q ),
    .c(_097_),
    .y(_193_)
  );
  al_inv _481_ (
    .a(\DFF_18.Q ),
    .y(_194_)
  );
  al_ao21 _482_ (
    .a(_191_),
    .b(_097_),
    .c(_194_),
    .y(_195_)
  );
  al_aoi21 _483_ (
    .a(_193_),
    .b(_195_),
    .c(_005_),
    .y(\DFF_18.D )
  );
  al_ao21 _484_ (
    .a(_194_),
    .b(_099_),
    .c(\DFF_19.Q ),
    .y(_196_)
  );
  al_and3 _485_ (
    .a(G14),
    .b(_100_),
    .c(_196_),
    .y(\DFF_19.D )
  );
  al_ao21ftf _486_ (
    .a(G7),
    .b(_052_),
    .c(_132_),
    .y(_197_)
  );
  al_and3ftt _487_ (
    .a(\DFF_1.D ),
    .b(\DFF_20.Q ),
    .c(_001_),
    .y(_198_)
  );
  al_ao21ftt _488_ (
    .a(\DFF_1.D ),
    .b(_001_),
    .c(\DFF_20.Q ),
    .y(_199_)
  );
  al_and3ftt _489_ (
    .a(_198_),
    .b(_199_),
    .c(_197_),
    .y(\DFF_20.D )
  );
  al_and2 _490_ (
    .a(\DFF_21.Q ),
    .b(_198_),
    .y(_200_)
  );
  al_or2 _491_ (
    .a(\DFF_21.Q ),
    .b(_198_),
    .y(_201_)
  );
  al_and3ftt _492_ (
    .a(_200_),
    .b(_201_),
    .c(_197_),
    .y(\DFF_21.D )
  );
  al_nand3 _493_ (
    .a(\DFF_21.Q ),
    .b(\DFF_22.Q ),
    .c(_198_),
    .y(_202_)
  );
  al_ao21 _494_ (
    .a(\DFF_21.Q ),
    .b(_198_),
    .c(\DFF_22.Q ),
    .y(_203_)
  );
  al_and3 _495_ (
    .a(_202_),
    .b(_203_),
    .c(_197_),
    .y(\DFF_22.D )
  );
  al_nand3 _496_ (
    .a(\DFF_22.Q ),
    .b(\DFF_23.Q ),
    .c(_200_),
    .y(_204_)
  );
  al_and2ft _497_ (
    .a(\DFF_23.Q ),
    .b(_202_),
    .y(_205_)
  );
  al_and3ftt _498_ (
    .a(_205_),
    .b(_197_),
    .c(_204_),
    .y(\DFF_23.D )
  );
  al_aoi21ttf _499_ (
    .a(_086_),
    .b(_204_),
    .c(_197_),
    .y(_206_)
  );
  al_aoi21ftf _500_ (
    .a(_204_),
    .b(\DFF_24.Q ),
    .c(_206_),
    .y(\DFF_24.D )
  );
  al_aoi21ttf _501_ (
    .a(\DFF_70.Q ),
    .b(_096_),
    .c(\DFF_32.Q ),
    .y(_207_)
  );
  al_ao21 _502_ (
    .a(\DFF_34.Q ),
    .b(_207_),
    .c(_108_),
    .y(_208_)
  );
  al_mux2l _503_ (
    .a(G12),
    .b(\DFF_25.Q ),
    .s(_208_),
    .y(_209_)
  );
  al_and2 _504_ (
    .a(G14),
    .b(_209_),
    .y(\DFF_25.D )
  );
  al_mux2l _505_ (
    .a(\DFF_25.Q ),
    .b(\DFF_26.Q ),
    .s(_208_),
    .y(_210_)
  );
  al_and2 _506_ (
    .a(G14),
    .b(_210_),
    .y(\DFF_26.D )
  );
  al_mux2l _507_ (
    .a(\DFF_26.Q ),
    .b(\DFF_27.Q ),
    .s(_208_),
    .y(_211_)
  );
  al_and2 _508_ (
    .a(G14),
    .b(_211_),
    .y(\DFF_27.D )
  );
  al_mux2l _509_ (
    .a(\DFF_27.Q ),
    .b(\DFF_28.Q ),
    .s(_208_),
    .y(_212_)
  );
  al_and2 _510_ (
    .a(G14),
    .b(_212_),
    .y(\DFF_28.D )
  );
  al_nand2 _511_ (
    .a(\DFF_69.Q ),
    .b(_104_),
    .y(_213_)
  );
  al_aoi21 _512_ (
    .a(\DFF_31.Q ),
    .b(_213_),
    .c(_005_),
    .y(_214_)
  );
  al_nand3fft _513_ (
    .a(_108_),
    .b(\DFF_29.Q ),
    .c(_104_),
    .y(_215_)
  );
  al_inv _514_ (
    .a(\DFF_29.Q ),
    .y(_216_)
  );
  al_ao21 _515_ (
    .a(\DFF_69.Q ),
    .b(_104_),
    .c(_216_),
    .y(_217_)
  );
  al_and3 _516_ (
    .a(_215_),
    .b(_217_),
    .c(_214_),
    .y(\DFF_29.D )
  );
  al_inv _517_ (
    .a(\DFF_30.Q ),
    .y(_218_)
  );
  al_nand3fft _518_ (
    .a(_216_),
    .b(_218_),
    .c(_213_),
    .y(_219_)
  );
  al_nand2 _519_ (
    .a(_218_),
    .b(_217_),
    .y(_220_)
  );
  al_and3 _520_ (
    .a(_219_),
    .b(_220_),
    .c(_214_),
    .y(\DFF_30.D )
  );
  al_aoi21ftf _521_ (
    .a(\DFF_31.Q ),
    .b(_219_),
    .c(_214_),
    .y(\DFF_31.D )
  );
  al_nand3fft _522_ (
    .a(_048_),
    .b(\DFF_32.Q ),
    .c(_096_),
    .y(_221_)
  );
  al_and3fft _523_ (
    .a(_005_),
    .b(_207_),
    .c(_221_),
    .y(\DFF_32.D )
  );
  al_aoi21 _524_ (
    .a(\DFF_34.Q ),
    .b(_207_),
    .c(_005_),
    .y(_222_)
  );
  al_nand3 _525_ (
    .a(\DFF_32.Q ),
    .b(\DFF_33.Q ),
    .c(_097_),
    .y(_223_)
  );
  al_ao21 _526_ (
    .a(\DFF_32.Q ),
    .b(_097_),
    .c(\DFF_33.Q ),
    .y(_224_)
  );
  al_and3 _527_ (
    .a(_223_),
    .b(_224_),
    .c(_222_),
    .y(\DFF_33.D )
  );
  al_aoi21ftf _528_ (
    .a(\DFF_34.Q ),
    .b(_223_),
    .c(_222_),
    .y(\DFF_34.D )
  );
  al_aoi21 _529_ (
    .a(\DFF_36.Q ),
    .b(_103_),
    .c(_005_),
    .y(_225_)
  );
  al_nand2 _530_ (
    .a(\DFF_35.Q ),
    .b(_103_),
    .y(_226_)
  );
  al_or2 _531_ (
    .a(\DFF_35.Q ),
    .b(_103_),
    .y(_227_)
  );
  al_and3 _532_ (
    .a(_226_),
    .b(_227_),
    .c(_225_),
    .y(\DFF_35.D )
  );
  al_aoi21ftf _533_ (
    .a(\DFF_36.Q ),
    .b(_226_),
    .c(_225_),
    .y(\DFF_36.D )
  );
  al_ao21 _534_ (
    .a(\DFF_36.Q ),
    .b(_103_),
    .c(\DFF_37.Q ),
    .y(_228_)
  );
  al_and3 _535_ (
    .a(G14),
    .b(_104_),
    .c(_228_),
    .y(\DFF_37.D )
  );
  al_aoi21 _536_ (
    .a(\DFF_39.Q ),
    .b(_105_),
    .c(_005_),
    .y(_229_)
  );
  al_nand3 _537_ (
    .a(\DFF_38.Q ),
    .b(\DFF_31.Q ),
    .c(_213_),
    .y(_230_)
  );
  al_ao21 _538_ (
    .a(\DFF_31.Q ),
    .b(_213_),
    .c(\DFF_38.Q ),
    .y(_231_)
  );
  al_and3 _539_ (
    .a(_230_),
    .b(_231_),
    .c(_229_),
    .y(\DFF_38.D )
  );
  al_aoi21ftf _540_ (
    .a(\DFF_39.Q ),
    .b(_230_),
    .c(_229_),
    .y(\DFF_39.D )
  );
  al_ao21 _541_ (
    .a(\DFF_39.Q ),
    .b(_105_),
    .c(\DFF_40.Q ),
    .y(_232_)
  );
  al_and3 _542_ (
    .a(G14),
    .b(_148_),
    .c(_232_),
    .y(\DFF_40.D )
  );
  al_dffl _543_ (
    .clk(CK),
    .d(\DFF_0.D ),
    .q(\DFF_0.Q )
  );
  al_dffl _544_ (
    .clk(CK),
    .d(\DFF_1.D ),
    .q(\DFF_1.Q )
  );
  al_dffl _545_ (
    .clk(CK),
    .d(\DFF_2.D ),
    .q(\DFF_2.Q )
  );
  al_dffl _546_ (
    .clk(CK),
    .d(\DFF_3.D ),
    .q(\DFF_3.Q )
  );
  al_dffl _547_ (
    .clk(CK),
    .d(\DFF_4.D ),
    .q(\DFF_4.Q )
  );
  al_dffl _548_ (
    .clk(CK),
    .d(\DFF_5.D ),
    .q(\DFF_5.Q )
  );
  al_dffl _549_ (
    .clk(CK),
    .d(\DFF_6.D ),
    .q(\DFF_6.Q )
  );
  al_dffl _550_ (
    .clk(CK),
    .d(\DFF_7.D ),
    .q(\DFF_7.Q )
  );
  al_dffl _551_ (
    .clk(CK),
    .d(\DFF_8.D ),
    .q(\DFF_8.Q )
  );
  al_dffl _552_ (
    .clk(CK),
    .d(\DFF_9.D ),
    .q(\DFF_9.Q )
  );
  al_dffl _553_ (
    .clk(CK),
    .d(\DFF_10.D ),
    .q(\DFF_10.Q )
  );
  al_dffl _554_ (
    .clk(CK),
    .d(\DFF_11.D ),
    .q(\DFF_11.Q )
  );
  al_dffl _555_ (
    .clk(CK),
    .d(\DFF_12.D ),
    .q(\DFF_12.Q )
  );
  al_dffl _556_ (
    .clk(CK),
    .d(\DFF_13.D ),
    .q(\DFF_13.Q )
  );
  al_dffl _557_ (
    .clk(CK),
    .d(\DFF_14.D ),
    .q(\DFF_14.Q )
  );
  al_dffl _558_ (
    .clk(CK),
    .d(\DFF_15.D ),
    .q(\DFF_15.Q )
  );
  al_dffl _559_ (
    .clk(CK),
    .d(\DFF_16.D ),
    .q(\DFF_16.Q )
  );
  al_dffl _560_ (
    .clk(CK),
    .d(\DFF_17.D ),
    .q(\DFF_17.Q )
  );
  al_dffl _561_ (
    .clk(CK),
    .d(\DFF_18.D ),
    .q(\DFF_18.Q )
  );
  al_dffl _562_ (
    .clk(CK),
    .d(\DFF_19.D ),
    .q(\DFF_19.Q )
  );
  al_dffl _563_ (
    .clk(CK),
    .d(\DFF_20.D ),
    .q(\DFF_20.Q )
  );
  al_dffl _564_ (
    .clk(CK),
    .d(\DFF_21.D ),
    .q(\DFF_21.Q )
  );
  al_dffl _565_ (
    .clk(CK),
    .d(\DFF_22.D ),
    .q(\DFF_22.Q )
  );
  al_dffl _566_ (
    .clk(CK),
    .d(\DFF_23.D ),
    .q(\DFF_23.Q )
  );
  al_dffl _567_ (
    .clk(CK),
    .d(\DFF_24.D ),
    .q(\DFF_24.Q )
  );
  al_dffl _568_ (
    .clk(CK),
    .d(\DFF_25.D ),
    .q(\DFF_25.Q )
  );
  al_dffl _569_ (
    .clk(CK),
    .d(\DFF_26.D ),
    .q(\DFF_26.Q )
  );
  al_dffl _570_ (
    .clk(CK),
    .d(\DFF_27.D ),
    .q(\DFF_27.Q )
  );
  al_dffl _571_ (
    .clk(CK),
    .d(\DFF_28.D ),
    .q(\DFF_28.Q )
  );
  al_dffl _572_ (
    .clk(CK),
    .d(\DFF_29.D ),
    .q(\DFF_29.Q )
  );
  al_dffl _573_ (
    .clk(CK),
    .d(\DFF_30.D ),
    .q(\DFF_30.Q )
  );
  al_dffl _574_ (
    .clk(CK),
    .d(\DFF_31.D ),
    .q(\DFF_31.Q )
  );
  al_dffl _575_ (
    .clk(CK),
    .d(\DFF_32.D ),
    .q(\DFF_32.Q )
  );
  al_dffl _576_ (
    .clk(CK),
    .d(\DFF_33.D ),
    .q(\DFF_33.Q )
  );
  al_dffl _577_ (
    .clk(CK),
    .d(\DFF_34.D ),
    .q(\DFF_34.Q )
  );
  al_dffl _578_ (
    .clk(CK),
    .d(\DFF_35.D ),
    .q(\DFF_35.Q )
  );
  al_dffl _579_ (
    .clk(CK),
    .d(\DFF_36.D ),
    .q(\DFF_36.Q )
  );
  al_dffl _580_ (
    .clk(CK),
    .d(\DFF_37.D ),
    .q(\DFF_37.Q )
  );
  al_dffl _581_ (
    .clk(CK),
    .d(\DFF_38.D ),
    .q(\DFF_38.Q )
  );
  al_dffl _582_ (
    .clk(CK),
    .d(\DFF_39.D ),
    .q(\DFF_39.Q )
  );
  al_dffl _583_ (
    .clk(CK),
    .d(\DFF_40.D ),
    .q(\DFF_40.Q )
  );
  al_dffl _584_ (
    .clk(CK),
    .d(\DFF_41.D ),
    .q(\DFF_41.Q )
  );
  al_dffl _585_ (
    .clk(CK),
    .d(\DFF_42.D ),
    .q(\DFF_42.Q )
  );
  al_dffl _586_ (
    .clk(CK),
    .d(\DFF_43.D ),
    .q(\DFF_43.Q )
  );
  al_dffl _587_ (
    .clk(CK),
    .d(\DFF_44.D ),
    .q(\DFF_44.Q )
  );
  al_dffl _588_ (
    .clk(CK),
    .d(\DFF_45.D ),
    .q(\DFF_45.Q )
  );
  al_dffl _589_ (
    .clk(CK),
    .d(\DFF_46.D ),
    .q(\DFF_46.Q )
  );
  al_dffl _590_ (
    .clk(CK),
    .d(\DFF_47.D ),
    .q(\DFF_47.Q )
  );
  al_dffl _591_ (
    .clk(CK),
    .d(\DFF_48.D ),
    .q(\DFF_48.Q )
  );
  al_dffl _592_ (
    .clk(CK),
    .d(\DFF_49.D ),
    .q(\DFF_49.Q )
  );
  al_dffl _593_ (
    .clk(CK),
    .d(\DFF_50.D ),
    .q(\DFF_50.Q )
  );
  al_dffl _594_ (
    .clk(CK),
    .d(\DFF_51.D ),
    .q(\DFF_51.Q )
  );
  al_dffl _595_ (
    .clk(CK),
    .d(\DFF_52.D ),
    .q(\DFF_52.Q )
  );
  al_dffl _596_ (
    .clk(CK),
    .d(\DFF_53.D ),
    .q(\DFF_53.Q )
  );
  al_dffl _597_ (
    .clk(CK),
    .d(\DFF_54.D ),
    .q(\DFF_54.Q )
  );
  al_dffl _598_ (
    .clk(CK),
    .d(\DFF_55.D ),
    .q(\DFF_55.Q )
  );
  al_dffl _599_ (
    .clk(CK),
    .d(\DFF_56.D ),
    .q(\DFF_56.Q )
  );
  al_dffl _600_ (
    .clk(CK),
    .d(\DFF_57.D ),
    .q(\DFF_57.Q )
  );
  al_dffl _601_ (
    .clk(CK),
    .d(\DFF_58.D ),
    .q(\DFF_58.Q )
  );
  al_dffl _602_ (
    .clk(CK),
    .d(\DFF_59.D ),
    .q(\DFF_59.Q )
  );
  al_dffl _603_ (
    .clk(CK),
    .d(\DFF_60.D ),
    .q(\DFF_60.Q )
  );
  al_dffl _604_ (
    .clk(CK),
    .d(\DFF_61.D ),
    .q(\DFF_61.Q )
  );
  al_dffl _605_ (
    .clk(CK),
    .d(\DFF_62.D ),
    .q(\DFF_62.Q )
  );
  al_dffl _606_ (
    .clk(CK),
    .d(\DFF_63.D ),
    .q(\DFF_63.Q )
  );
  al_dffl _607_ (
    .clk(CK),
    .d(\DFF_64.D ),
    .q(\DFF_64.Q )
  );
  al_dffl _608_ (
    .clk(CK),
    .d(\DFF_65.D ),
    .q(\DFF_65.Q )
  );
  al_dffl _609_ (
    .clk(CK),
    .d(\DFF_66.D ),
    .q(\DFF_66.Q )
  );
  al_dffl _610_ (
    .clk(CK),
    .d(\DFF_67.D ),
    .q(\DFF_67.Q )
  );
  al_dffl _611_ (
    .clk(CK),
    .d(\DFF_68.D ),
    .q(\DFF_68.Q )
  );
  al_dffl _612_ (
    .clk(CK),
    .d(\DFF_69.D ),
    .q(\DFF_69.Q )
  );
  al_dffl _613_ (
    .clk(CK),
    .d(\DFF_70.D ),
    .q(\DFF_70.Q )
  );
  al_dffl _614_ (
    .clk(CK),
    .d(\DFF_71.D ),
    .q(\DFF_71.Q )
  );
  al_dffl _615_ (
    .clk(CK),
    .d(\DFF_72.D ),
    .q(\DFF_72.Q )
  );
  al_dffl _616_ (
    .clk(CK),
    .d(\DFF_73.D ),
    .q(\DFF_73.Q )
  );
  assign \DFF_0.CK  = CK;
  assign \DFF_1.CK  = CK;
  assign \DFF_10.CK  = CK;
  assign \DFF_11.CK  = CK;
  assign \DFF_12.CK  = CK;
  assign \DFF_13.CK  = CK;
  assign \DFF_14.CK  = CK;
  assign \DFF_15.CK  = CK;
  assign \DFF_16.CK  = CK;
  assign \DFF_17.CK  = CK;
  assign \DFF_18.CK  = CK;
  assign \DFF_19.CK  = CK;
  assign \DFF_2.CK  = CK;
  assign \DFF_20.CK  = CK;
  assign \DFF_21.CK  = CK;
  assign \DFF_22.CK  = CK;
  assign \DFF_23.CK  = CK;
  assign \DFF_24.CK  = CK;
  assign \DFF_25.CK  = CK;
  assign \DFF_26.CK  = CK;
  assign \DFF_27.CK  = CK;
  assign \DFF_28.CK  = CK;
  assign \DFF_29.CK  = CK;
  assign \DFF_3.CK  = CK;
  assign \DFF_30.CK  = CK;
  assign \DFF_31.CK  = CK;
  assign \DFF_32.CK  = CK;
  assign \DFF_33.CK  = CK;
  assign \DFF_34.CK  = CK;
  assign \DFF_35.CK  = CK;
  assign \DFF_36.CK  = CK;
  assign \DFF_37.CK  = CK;
  assign \DFF_38.CK  = CK;
  assign \DFF_39.CK  = CK;
  assign \DFF_4.CK  = CK;
  assign \DFF_40.CK  = CK;
  assign \DFF_41.CK  = CK;
  assign \DFF_42.CK  = CK;
  assign \DFF_43.CK  = CK;
  assign \DFF_44.CK  = CK;
  assign \DFF_45.CK  = CK;
  assign \DFF_46.CK  = CK;
  assign \DFF_47.CK  = CK;
  assign \DFF_48.CK  = CK;
  assign \DFF_49.CK  = CK;
  assign \DFF_5.CK  = CK;
  assign \DFF_50.CK  = CK;
  assign \DFF_51.CK  = CK;
  assign \DFF_52.CK  = CK;
  assign \DFF_53.CK  = CK;
  assign \DFF_54.CK  = CK;
  assign \DFF_55.CK  = CK;
  assign \DFF_56.CK  = CK;
  assign \DFF_57.CK  = CK;
  assign \DFF_58.CK  = CK;
  assign \DFF_59.CK  = CK;
  assign \DFF_6.CK  = CK;
  assign \DFF_60.CK  = CK;
  assign \DFF_61.CK  = CK;
  assign \DFF_62.CK  = CK;
  assign \DFF_63.CK  = CK;
  assign \DFF_64.CK  = CK;
  assign \DFF_65.CK  = CK;
  assign \DFF_66.CK  = CK;
  assign \DFF_67.CK  = CK;
  assign \DFF_68.CK  = CK;
  assign \DFF_69.CK  = CK;
  assign \DFF_7.CK  = CK;
  assign \DFF_70.CK  = CK;
  assign \DFF_71.CK  = CK;
  assign \DFF_72.CK  = CK;
  assign \DFF_73.CK  = CK;
  assign \DFF_8.CK  = CK;
  assign \DFF_9.CK  = CK;
  assign G108 = G14;
  assign G109 = \DFF_2.D ;
  assign G112 = G14;
  assign G113 = \DFF_3.D ;
  assign G117 = G14;
  assign G118 = \DFF_4.D ;
  assign G124 = G14;
  assign G125 = \DFF_5.D ;
  assign G128 = G14;
  assign G129 = \DFF_6.D ;
  assign G139 = G14;
  assign G140 = \DFF_7.D ;
  assign G143 = G14;
  assign G144 = \DFF_8.D ;
  assign G148 = G14;
  assign G149 = \DFF_9.D ;
  assign G153 = G14;
  assign G154 = \DFF_10.D ;
  assign G158 = G14;
  assign G159 = \DFF_11.D ;
  assign G165 = G14;
  assign G166 = \DFF_12.D ;
  assign G174 = G14;
  assign G175 = \DFF_13.D ;
  assign G179 = \DFF_70.Q ;
  assign G188 = G14;
  assign G189 = \DFF_14.D ;
  assign G192 = G14;
  assign G193 = \DFF_15.D ;
  assign G197 = G14;
  assign G198 = \DFF_16.D ;
  assign G207 = G14;
  assign G208 = \DFF_17.D ;
  assign G213 = G14;
  assign G214 = \DFF_18.D ;
  assign G217 = G14;
  assign G218 = \DFF_19.D ;
  assign G22 = \DFF_0.Q ;
  assign G23 = \DFF_1.Q ;
  assign G237 = \DFF_20.D ;
  assign G24 = \DFF_2.Q ;
  assign G242 = \DFF_21.D ;
  assign G247 = \DFF_22.D ;
  assign G25 = \DFF_3.Q ;
  assign G252 = \DFF_23.D ;
  assign G26 = \DFF_4.Q ;
  assign G260 = \DFF_24.D ;
  assign G27 = \DFF_5.Q ;
  assign G28 = \DFF_6.Q ;
  assign G29 = \DFF_7.Q ;
  assign G30 = \DFF_8.Q ;
  assign G302 = G14;
  assign G303 = \DFF_25.D ;
  assign G308 = G14;
  assign G309 = \DFF_26.D ;
  assign G31 = \DFF_9.Q ;
  assign G314 = G14;
  assign G315 = \DFF_27.D ;
  assign G32 = \DFF_10.Q ;
  assign G320 = G14;
  assign G321 = \DFF_28.D ;
  assign G328 = \DFF_1.D ;
  assign G328BF = \DFF_1.D ;
  assign G33 = \DFF_11.Q ;
  assign G332 = \DFF_0.D ;
  assign G332BF = \DFF_0.D ;
  assign G34 = \DFF_12.Q ;
  assign G343 = \DFF_69.Q ;
  assign G347 = \DFF_69.Q ;
  assign G35 = \DFF_13.Q ;
  assign G351 = \DFF_68.Q ;
  assign G36 = \DFF_14.Q ;
  assign G360 = \DFF_29.D ;
  assign G365 = \DFF_30.D ;
  assign G37 = \DFF_15.Q ;
  assign G373 = \DFF_31.D ;
  assign G379 = \DFF_32.D ;
  assign G38 = \DFF_16.Q ;
  assign G384 = \DFF_33.D ;
  assign G39 = \DFF_17.Q ;
  assign G392 = \DFF_34.D ;
  assign G397 = \DFF_35.D ;
  assign G40 = \DFF_18.Q ;
  assign G405 = \DFF_36.D ;
  assign G407 = G14;
  assign G408 = \DFF_37.D ;
  assign G41 = \DFF_19.Q ;
  assign G416 = \DFF_38.D ;
  assign G42 = \DFF_20.Q ;
  assign G424 = \DFF_39.D ;
  assign G426 = G14;
  assign G427 = \DFF_40.D ;
  assign G43 = \DFF_21.Q ;
  assign G437 = G14;
  assign G438 = \DFF_41.D ;
  assign G44 = \DFF_22.Q ;
  assign G440 = G14;
  assign G441 = \DFF_42.D ;
  assign G446 = G14;
  assign G447 = \DFF_43.D ;
  assign G45 = \DFF_23.Q ;
  assign G450 = G14;
  assign G451 = \DFF_44.D ;
  assign G459 = \DFF_45.D ;
  assign G46 = \DFF_24.Q ;
  assign G464 = \DFF_46.D ;
  assign G469 = \DFF_47.D ;
  assign G47 = \DFF_25.Q ;
  assign G477 = \DFF_48.D ;
  assign G48 = \DFF_26.Q ;
  assign G486 = G14;
  assign G49 = \DFF_27.Q ;
  assign G494 = \DFF_49.D ;
  assign G498 = \DFF_50.D ;
  assign G50 = \DFF_28.Q ;
  assign G503 = \DFF_51.D ;
  assign G504 = \DFF_41.Q ;
  assign G507 = \DFF_41.Q ;
  assign G51 = \DFF_29.Q ;
  assign G510 = \DFF_41.Q ;
  assign G52 = \DFF_30.Q ;
  assign G526 = \DFF_52.D ;
  assign G53 = \DFF_31.Q ;
  assign G531 = \DFF_53.D ;
  assign G536 = \DFF_54.D ;
  assign G54 = \DFF_32.Q ;
  assign G541 = \DFF_55.D ;
  assign G548 = \DFF_56.D ;
  assign G55 = \DFF_33.Q ;
  assign G56 = \DFF_34.Q ;
  assign G565 = \DFF_57.D ;
  assign G569 = \DFF_58.D ;
  assign G57 = \DFF_35.Q ;
  assign G573 = \DFF_59.D ;
  assign G577 = \DFF_60.D ;
  assign G58 = \DFF_36.Q ;
  assign G59 = \DFF_37.Q ;
  assign G590 = \DFF_61.D ;
  assign G60 = \DFF_38.Q ;
  assign G608 = \DFF_62.D ;
  assign G61 = \DFF_39.Q ;
  assign G613 = \DFF_63.D ;
  assign G617 = \DFF_68.Q ;
  assign G62 = \DFF_40.Q ;
  assign G620 = \DFF_68.Q ;
  assign G623 = \DFF_68.Q ;
  assign G626 = \DFF_68.Q ;
  assign G629 = \DFF_68.Q ;
  assign G63 = \DFF_41.Q ;
  assign G632 = \DFF_68.Q ;
  assign G635 = \DFF_68.Q ;
  assign G638 = \DFF_68.Q ;
  assign G64 = \DFF_42.Q ;
  assign G641 = \DFF_68.Q ;
  assign G644 = \DFF_68.Q ;
  assign G65 = \DFF_43.Q ;
  assign G656 = G14;
  assign G657 = \DFF_64.D ;
  assign G659 = G13;
  assign G66 = \DFF_44.Q ;
  assign G662 = G14;
  assign G663 = \DFF_65.D ;
  assign G668 = G14;
  assign G669 = \DFF_66.D ;
  assign G67 = \DFF_45.Q ;
  assign G674 = G14;
  assign G675 = \DFF_67.D ;
  assign G678 = G11;
  assign G68 = \DFF_46.Q ;
  assign G682 = \DFF_68.D ;
  assign G687 = \DFF_69.D ;
  assign G69 = \DFF_47.Q ;
  assign G693 = \DFF_70.D ;
  assign G696 = G10;
  assign G70 = \DFF_48.Q ;
  assign G701 = G701BF;
  assign G704 = G14;
  assign G705 = \DFF_71.D ;
  assign G706 = G14;
  assign G707 = \DFF_72.D ;
  assign G71 = \DFF_49.Q ;
  assign G711 = G14;
  assign G713 = \DFF_73.D ;
  assign G714 = G15;
  assign G715 = G6;
  assign G716 = G7;
  assign G717 = G8;
  assign G718 = G9;
  assign G719 = G12;
  assign G72 = \DFF_50.Q ;
  assign G720 = G0;
  assign G721 = G1;
  assign G722 = G2;
  assign G723 = G3;
  assign G724 = G4;
  assign G725 = G5;
  assign G726 = \DFF_71.Q ;
  assign G728 = G16;
  assign G729 = \DFF_73.Q ;
  assign G73 = \DFF_51.Q ;
  assign G74 = \DFF_52.Q ;
  assign G75 = \DFF_53.Q ;
  assign G76 = \DFF_54.Q ;
  assign G77 = \DFF_55.Q ;
  assign G78 = \DFF_56.Q ;
  assign G79 = \DFF_57.Q ;
  assign G80 = \DFF_58.Q ;
  assign G81 = \DFF_59.Q ;
  assign G82 = \DFF_60.Q ;
  assign G83 = \DFF_61.Q ;
  assign G84 = \DFF_62.Q ;
  assign G85 = \DFF_63.Q ;
  assign G86 = \DFF_64.Q ;
  assign G87 = \DFF_65.Q ;
  assign G88 = \DFF_66.Q ;
  assign G89 = \DFF_67.Q ;
  assign G90 = \DFF_68.Q ;
  assign G91 = \DFF_69.Q ;
  assign G92 = \DFF_70.Q ;
  assign G93 = \DFF_71.Q ;
  assign G94 = \DFF_72.Q ;
  assign G95 = \DFF_73.Q ;
  assign II1211 = G15;
endmodule
